
module AES_HPC2_BDDcudd_ClockGating_d1 ( plaintext_s0, key_s0, clk, start, 
        plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1, Synch
 );
  input [127:0] plaintext_s0;
  input [127:0] key_s0;
  input [127:0] plaintext_s1;
  input [127:0] key_s1;
  input [413:0] Fresh;
  output [127:0] ciphertext_s0;
  output [127:0] ciphertext_s1;
  input clk, start;
  output done, Synch;
  wire   signal_2390, signal_1413, signal_2389, signal_1493, signal_2393,
         signal_1412, signal_2392, signal_1492, signal_2396, signal_1411,
         signal_2395, signal_1491, signal_2399, signal_1410, signal_2398,
         signal_1490, signal_2402, signal_1409, signal_2401, signal_1489,
         signal_2405, signal_1408, signal_2404, signal_1488, signal_2408,
         signal_1407, signal_2407, signal_1487, signal_2411, signal_1406,
         signal_2410, signal_1486, signal_399, signal_400, signal_421,
         signal_420, signal_419, signal_418, signal_429, signal_431,
         signal_433, signal_435, signal_437, signal_439, signal_441,
         signal_3786, signal_465, signal_2562, signal_1677, signal_3787,
         signal_467, signal_2565, signal_1676, signal_3788, signal_469,
         signal_2568, signal_1675, signal_3789, signal_471, signal_2571,
         signal_1674, signal_3790, signal_473, signal_2574, signal_1673,
         signal_3791, signal_475, signal_2577, signal_1672, signal_3792,
         signal_477, signal_2580, signal_1671, signal_3793, signal_479,
         signal_2583, signal_1670, signal_3794, signal_481, signal_2586,
         signal_1669, signal_3795, signal_483, signal_2589, signal_1668,
         signal_3796, signal_485, signal_2592, signal_1667, signal_3797,
         signal_487, signal_2595, signal_1666, signal_3798, signal_489,
         signal_2598, signal_1665, signal_3799, signal_491, signal_2601,
         signal_1664, signal_3800, signal_493, signal_2604, signal_1663,
         signal_3801, signal_495, signal_2607, signal_1662, signal_3802,
         signal_497, signal_2610, signal_1661, signal_3803, signal_499,
         signal_2613, signal_1660, signal_3804, signal_501, signal_2616,
         signal_1659, signal_3805, signal_503, signal_2619, signal_1658,
         signal_3806, signal_505, signal_2622, signal_1657, signal_3807,
         signal_507, signal_2625, signal_1656, signal_3808, signal_509,
         signal_2628, signal_1655, signal_3809, signal_511, signal_2631,
         signal_1654, signal_3810, signal_513, signal_3592, signal_1653,
         signal_3811, signal_515, signal_3594, signal_1652, signal_3812,
         signal_517, signal_3596, signal_1651, signal_3813, signal_519,
         signal_3598, signal_1650, signal_3814, signal_521, signal_3600,
         signal_1649, signal_3815, signal_523, signal_3602, signal_1648,
         signal_3816, signal_525, signal_3604, signal_1647, signal_3817,
         signal_527, signal_3606, signal_1646, signal_3818, signal_529,
         signal_2634, signal_1645, signal_3819, signal_531, signal_2637,
         signal_1644, signal_3820, signal_533, signal_2640, signal_1643,
         signal_3821, signal_535, signal_2643, signal_1642, signal_3822,
         signal_537, signal_2646, signal_1641, signal_3823, signal_539,
         signal_2649, signal_1640, signal_3824, signal_541, signal_2652,
         signal_1639, signal_3825, signal_543, signal_2655, signal_1638,
         signal_3826, signal_545, signal_2658, signal_1637, signal_3827,
         signal_547, signal_2661, signal_1636, signal_3828, signal_549,
         signal_2664, signal_1635, signal_3829, signal_551, signal_2667,
         signal_1634, signal_3830, signal_553, signal_2670, signal_1633,
         signal_3831, signal_555, signal_2673, signal_1632, signal_3832,
         signal_557, signal_2676, signal_1631, signal_3833, signal_559,
         signal_2679, signal_1630, signal_3834, signal_561, signal_2682,
         signal_1629, signal_3835, signal_563, signal_2685, signal_1628,
         signal_3836, signal_565, signal_2688, signal_1627, signal_3837,
         signal_567, signal_2691, signal_1626, signal_3838, signal_569,
         signal_2694, signal_1625, signal_3839, signal_571, signal_2697,
         signal_1624, signal_3840, signal_573, signal_2700, signal_1623,
         signal_3841, signal_575, signal_2703, signal_1622, signal_3842,
         signal_577, signal_3608, signal_1621, signal_3843, signal_579,
         signal_3610, signal_1620, signal_3844, signal_581, signal_3612,
         signal_1619, signal_3845, signal_583, signal_3614, signal_1618,
         signal_3846, signal_585, signal_3616, signal_1617, signal_3847,
         signal_587, signal_3618, signal_1616, signal_3848, signal_589,
         signal_3620, signal_1615, signal_3849, signal_591, signal_3622,
         signal_1614, signal_3850, signal_593, signal_2706, signal_1613,
         signal_3851, signal_595, signal_2709, signal_1612, signal_3852,
         signal_597, signal_2712, signal_1611, signal_3853, signal_599,
         signal_2715, signal_1610, signal_3854, signal_601, signal_2718,
         signal_1609, signal_3855, signal_603, signal_2721, signal_1608,
         signal_3856, signal_605, signal_2724, signal_1607, signal_3857,
         signal_607, signal_2727, signal_1606, signal_3858, signal_609,
         signal_2730, signal_1605, signal_3859, signal_611, signal_2733,
         signal_1604, signal_3860, signal_613, signal_2736, signal_1603,
         signal_3861, signal_615, signal_2739, signal_1602, signal_3862,
         signal_617, signal_2742, signal_1601, signal_3863, signal_619,
         signal_2745, signal_1600, signal_3864, signal_621, signal_2748,
         signal_1599, signal_3865, signal_623, signal_2751, signal_1598,
         signal_3866, signal_625, signal_2754, signal_1597, signal_3867,
         signal_627, signal_2757, signal_1596, signal_3868, signal_629,
         signal_2760, signal_1595, signal_3869, signal_631, signal_2763,
         signal_1594, signal_3870, signal_633, signal_2766, signal_1593,
         signal_3871, signal_635, signal_2769, signal_1592, signal_3872,
         signal_637, signal_2772, signal_1591, signal_3873, signal_639,
         signal_2775, signal_1590, signal_3874, signal_641, signal_3624,
         signal_1589, signal_3875, signal_643, signal_3626, signal_1588,
         signal_3876, signal_645, signal_3628, signal_1587, signal_3877,
         signal_647, signal_3630, signal_1586, signal_3878, signal_649,
         signal_3632, signal_1585, signal_3879, signal_651, signal_3634,
         signal_1584, signal_3880, signal_653, signal_3636, signal_1583,
         signal_3881, signal_655, signal_3638, signal_1582, signal_3882,
         signal_657, signal_2778, signal_1581, signal_3883, signal_659,
         signal_2781, signal_1580, signal_3884, signal_661, signal_2784,
         signal_1579, signal_3885, signal_663, signal_2787, signal_1578,
         signal_3886, signal_665, signal_2790, signal_1577, signal_3887,
         signal_667, signal_2793, signal_1576, signal_3888, signal_669,
         signal_2796, signal_1575, signal_3889, signal_671, signal_2799,
         signal_1574, signal_3890, signal_673, signal_2802, signal_1573,
         signal_3891, signal_675, signal_2805, signal_1572, signal_3892,
         signal_677, signal_2808, signal_1571, signal_3893, signal_679,
         signal_2811, signal_1570, signal_3894, signal_681, signal_2814,
         signal_1569, signal_3895, signal_683, signal_2817, signal_1568,
         signal_3896, signal_685, signal_2820, signal_1567, signal_3897,
         signal_687, signal_2823, signal_1566, signal_3898, signal_689,
         signal_2826, signal_1565, signal_3899, signal_691, signal_2829,
         signal_1564, signal_3900, signal_693, signal_2832, signal_1563,
         signal_3901, signal_695, signal_2835, signal_1562, signal_3902,
         signal_697, signal_2838, signal_1561, signal_3903, signal_699,
         signal_2841, signal_1560, signal_3904, signal_701, signal_2844,
         signal_1559, signal_3905, signal_703, signal_2847, signal_1558,
         signal_3434, signal_1549, signal_3282, signal_1429, signal_3435,
         signal_1548, signal_3283, signal_1428, signal_3436, signal_1547,
         signal_3284, signal_1427, signal_3437, signal_1546, signal_3285,
         signal_1426, signal_3438, signal_1545, signal_3286, signal_1425,
         signal_3439, signal_1544, signal_3287, signal_1424, signal_3440,
         signal_1543, signal_3288, signal_1423, signal_3441, signal_1542,
         signal_3289, signal_1422, signal_3442, signal_1541, signal_3274,
         signal_1437, signal_3443, signal_1540, signal_3275, signal_1436,
         signal_3444, signal_1539, signal_3276, signal_1435, signal_3445,
         signal_1538, signal_3277, signal_1434, signal_3446, signal_1537,
         signal_3278, signal_1433, signal_3447, signal_1536, signal_3279,
         signal_1432, signal_3448, signal_1535, signal_3280, signal_1431,
         signal_3449, signal_1534, signal_3281, signal_1430, signal_3450,
         signal_1533, signal_3266, signal_1445, signal_3451, signal_1532,
         signal_3267, signal_1444, signal_3452, signal_1531, signal_3268,
         signal_1443, signal_3453, signal_1530, signal_3269, signal_1442,
         signal_3454, signal_1529, signal_3270, signal_1441, signal_3455,
         signal_1528, signal_3271, signal_1440, signal_3456, signal_1527,
         signal_3272, signal_1439, signal_3457, signal_1526, signal_3273,
         signal_1438, signal_3262, signal_1453, signal_3231, signal_1485,
         signal_3263, signal_1452, signal_3255, signal_1484, signal_3240,
         signal_1451, signal_3229, signal_1483, signal_3264, signal_1450,
         signal_3254, signal_1482, signal_3265, signal_1449, signal_3253,
         signal_1481, signal_3241, signal_1448, signal_3226, signal_1480,
         signal_3242, signal_1447, signal_3225, signal_1479, signal_3243,
         signal_1446, signal_3224, signal_1478, signal_3223, signal_1477,
         signal_3252, signal_1476, signal_3221, signal_1475, signal_3251,
         signal_1474, signal_3250, signal_1473, signal_3218, signal_1472,
         signal_3217, signal_1471, signal_3216, signal_1470, signal_3215,
         signal_1469, signal_3249, signal_1468, signal_3213, signal_1467,
         signal_3248, signal_1466, signal_3247, signal_1465, signal_3210,
         signal_1464, signal_3209, signal_1463, signal_3208, signal_1462,
         signal_3207, signal_1461, signal_3246, signal_1460, signal_3205,
         signal_1459, signal_3245, signal_1458, signal_3244, signal_1457,
         signal_3202, signal_1456, signal_3201, signal_1455, signal_3200,
         signal_1454, signal_2413, signal_1686, signal_2412, signal_765,
         signal_2415, signal_1687, signal_2414, signal_764, signal_2417,
         signal_1688, signal_2416, signal_763, signal_2419, signal_1689,
         signal_2418, signal_762, signal_2421, signal_1690, signal_2420,
         signal_761, signal_2423, signal_1691, signal_2422, signal_760,
         signal_2425, signal_1692, signal_2424, signal_759, signal_2427,
         signal_1693, signal_2426, signal_758, signal_4122, signal_766,
         signal_3986, signal_767, signal_2897, signal_1877, signal_3907,
         signal_1933, signal_4123, signal_769, signal_3987, signal_770,
         signal_2900, signal_1876, signal_3909, signal_1932, signal_4124,
         signal_772, signal_3988, signal_773, signal_2903, signal_1875,
         signal_3911, signal_1931, signal_4125, signal_775, signal_3989,
         signal_776, signal_2906, signal_1874, signal_3913, signal_1930,
         signal_4126, signal_778, signal_3990, signal_779, signal_2909,
         signal_1873, signal_3915, signal_1929, signal_4127, signal_781,
         signal_3991, signal_782, signal_2912, signal_1872, signal_3917,
         signal_1928, signal_4128, signal_784, signal_3992, signal_785,
         signal_2915, signal_1871, signal_3919, signal_1927, signal_4129,
         signal_787, signal_3993, signal_788, signal_2918, signal_1870,
         signal_3921, signal_1926, signal_3994, signal_790, signal_3290,
         signal_791, signal_2921, signal_1861, signal_2850, signal_1925,
         signal_3995, signal_793, signal_3291, signal_794, signal_2924,
         signal_1860, signal_2853, signal_1924, signal_3996, signal_796,
         signal_3292, signal_797, signal_2927, signal_1859, signal_2856,
         signal_1923, signal_3997, signal_799, signal_3293, signal_800,
         signal_2930, signal_1858, signal_2859, signal_1922, signal_3998,
         signal_802, signal_3294, signal_803, signal_2933, signal_1857,
         signal_2862, signal_1921, signal_3999, signal_805, signal_3295,
         signal_806, signal_2936, signal_1856, signal_2865, signal_1920,
         signal_4000, signal_808, signal_3296, signal_809, signal_2939,
         signal_1855, signal_2868, signal_1919, signal_4001, signal_811,
         signal_3297, signal_812, signal_2942, signal_1854, signal_2871,
         signal_1918, signal_4002, signal_814, signal_3298, signal_815,
         signal_2849, signal_1909, signal_2945, signal_1845, signal_2874,
         signal_1917, signal_4003, signal_817, signal_3299, signal_818,
         signal_2852, signal_1908, signal_2948, signal_1844, signal_2877,
         signal_1916, signal_4004, signal_820, signal_3300, signal_821,
         signal_2855, signal_1907, signal_2951, signal_1843, signal_2880,
         signal_1915, signal_4005, signal_823, signal_3301, signal_824,
         signal_2858, signal_1906, signal_2954, signal_1842, signal_2883,
         signal_1914, signal_4006, signal_826, signal_3302, signal_827,
         signal_2861, signal_1905, signal_2957, signal_1841, signal_2886,
         signal_1913, signal_4007, signal_829, signal_3303, signal_830,
         signal_2864, signal_1904, signal_2960, signal_1840, signal_2889,
         signal_1912, signal_4008, signal_832, signal_3304, signal_833,
         signal_2867, signal_1903, signal_2963, signal_1839, signal_2892,
         signal_1911, signal_4009, signal_835, signal_3305, signal_836,
         signal_2870, signal_1902, signal_2966, signal_1838, signal_2895,
         signal_1910, signal_4010, signal_838, signal_3306, signal_839,
         signal_2873, signal_1893, signal_2969, signal_1509, signal_2898,
         signal_1901, signal_4011, signal_841, signal_3307, signal_842,
         signal_2876, signal_1892, signal_2972, signal_1508, signal_2901,
         signal_1900, signal_4012, signal_844, signal_3308, signal_845,
         signal_2879, signal_1891, signal_2975, signal_1507, signal_2904,
         signal_1899, signal_4013, signal_847, signal_3309, signal_848,
         signal_2882, signal_1890, signal_2978, signal_1506, signal_2907,
         signal_1898, signal_4014, signal_850, signal_3310, signal_851,
         signal_2885, signal_1889, signal_2981, signal_1505, signal_2910,
         signal_1897, signal_4015, signal_853, signal_3311, signal_854,
         signal_2888, signal_1888, signal_2984, signal_1504, signal_2913,
         signal_1896, signal_4016, signal_856, signal_3312, signal_857,
         signal_2891, signal_1887, signal_2987, signal_1503, signal_2916,
         signal_1895, signal_4017, signal_859, signal_3313, signal_860,
         signal_2894, signal_1886, signal_2990, signal_1502, signal_2919,
         signal_1894, signal_4018, signal_862, signal_3314, signal_863,
         signal_2993, signal_1821, signal_2922, signal_1885, signal_4019,
         signal_865, signal_3315, signal_866, signal_2996, signal_1820,
         signal_2925, signal_1884, signal_4020, signal_868, signal_3316,
         signal_869, signal_2999, signal_1819, signal_2928, signal_1883,
         signal_4021, signal_871, signal_3317, signal_872, signal_3002,
         signal_1818, signal_2931, signal_1882, signal_4022, signal_874,
         signal_3318, signal_875, signal_3005, signal_1817, signal_2934,
         signal_1881, signal_4023, signal_877, signal_3319, signal_878,
         signal_3008, signal_1816, signal_2937, signal_1880, signal_4024,
         signal_880, signal_3320, signal_881, signal_3011, signal_1815,
         signal_2940, signal_1879, signal_4025, signal_883, signal_3321,
         signal_884, signal_3014, signal_1814, signal_2943, signal_1878,
         signal_4026, signal_886, signal_3322, signal_887, signal_3017,
         signal_1805, signal_2946, signal_1869, signal_4027, signal_889,
         signal_3323, signal_890, signal_3020, signal_1804, signal_2949,
         signal_1868, signal_4028, signal_892, signal_3324, signal_893,
         signal_3023, signal_1803, signal_2952, signal_1867, signal_4029,
         signal_895, signal_3325, signal_896, signal_3026, signal_1802,
         signal_2955, signal_1866, signal_4030, signal_898, signal_3326,
         signal_899, signal_3029, signal_1801, signal_2958, signal_1865,
         signal_4031, signal_901, signal_3327, signal_902, signal_3032,
         signal_1800, signal_2961, signal_1864, signal_4032, signal_904,
         signal_3328, signal_905, signal_3035, signal_1799, signal_2964,
         signal_1863, signal_4033, signal_907, signal_3329, signal_908,
         signal_3038, signal_1798, signal_2967, signal_1862, signal_3639,
         signal_910, signal_3330, signal_911, signal_3041, signal_1789,
         signal_2970, signal_1853, signal_3640, signal_913, signal_3331,
         signal_914, signal_3044, signal_1788, signal_2973, signal_1852,
         signal_3641, signal_916, signal_3332, signal_917, signal_3047,
         signal_1787, signal_2976, signal_1851, signal_3642, signal_919,
         signal_3333, signal_920, signal_3050, signal_1786, signal_2979,
         signal_1850, signal_3643, signal_922, signal_3334, signal_923,
         signal_3053, signal_1785, signal_2982, signal_1849, signal_3644,
         signal_925, signal_3335, signal_926, signal_3056, signal_1784,
         signal_2985, signal_1848, signal_3645, signal_928, signal_3336,
         signal_929, signal_3059, signal_1783, signal_2988, signal_1847,
         signal_3646, signal_931, signal_3337, signal_932, signal_3062,
         signal_1782, signal_2991, signal_1846, signal_3647, signal_934,
         signal_3338, signal_935, signal_3065, signal_1773, signal_2994,
         signal_1837, signal_3648, signal_937, signal_3339, signal_938,
         signal_3068, signal_1772, signal_2997, signal_1836, signal_3649,
         signal_940, signal_3340, signal_941, signal_3071, signal_1771,
         signal_3000, signal_1835, signal_3650, signal_943, signal_3341,
         signal_944, signal_3074, signal_1770, signal_3003, signal_1834,
         signal_3651, signal_946, signal_3342, signal_947, signal_3077,
         signal_1769, signal_3006, signal_1833, signal_3652, signal_949,
         signal_3343, signal_950, signal_3080, signal_1768, signal_3009,
         signal_1832, signal_3653, signal_952, signal_3344, signal_953,
         signal_3083, signal_1767, signal_3012, signal_1831, signal_3654,
         signal_955, signal_3345, signal_956, signal_3086, signal_1766,
         signal_3015, signal_1830, signal_4034, signal_958, signal_3346,
         signal_959, signal_3089, signal_1749, signal_3018, signal_1829,
         signal_4035, signal_961, signal_3347, signal_962, signal_3092,
         signal_1748, signal_3021, signal_1828, signal_4036, signal_964,
         signal_3348, signal_965, signal_3095, signal_1747, signal_3024,
         signal_1827, signal_4037, signal_967, signal_3349, signal_968,
         signal_3098, signal_1746, signal_3027, signal_1826, signal_4038,
         signal_970, signal_3350, signal_971, signal_3101, signal_1745,
         signal_3030, signal_1825, signal_4039, signal_973, signal_3351,
         signal_974, signal_3104, signal_1744, signal_3033, signal_1824,
         signal_4040, signal_976, signal_3352, signal_977, signal_3107,
         signal_1743, signal_3036, signal_1823, signal_4041, signal_979,
         signal_3353, signal_980, signal_3110, signal_1742, signal_3039,
         signal_1822, signal_4042, signal_982, signal_3354, signal_983,
         signal_3113, signal_1733, signal_3042, signal_1813, signal_4043,
         signal_985, signal_3355, signal_986, signal_3116, signal_1732,
         signal_3045, signal_1812, signal_4044, signal_988, signal_3356,
         signal_989, signal_3119, signal_1731, signal_3048, signal_1811,
         signal_4045, signal_991, signal_3357, signal_992, signal_3122,
         signal_1730, signal_3051, signal_1810, signal_4046, signal_994,
         signal_3358, signal_995, signal_3125, signal_1729, signal_3054,
         signal_1809, signal_4047, signal_997, signal_3359, signal_998,
         signal_3128, signal_1728, signal_3057, signal_1808, signal_4048,
         signal_1000, signal_3360, signal_1001, signal_3131, signal_1727,
         signal_3060, signal_1807, signal_4049, signal_1003, signal_3361,
         signal_1004, signal_3134, signal_1726, signal_3063, signal_1806,
         signal_4050, signal_1006, signal_3362, signal_1007, signal_3137,
         signal_1717, signal_3066, signal_1797, signal_4051, signal_1009,
         signal_3363, signal_1010, signal_3140, signal_1716, signal_3069,
         signal_1796, signal_4052, signal_1012, signal_3364, signal_1013,
         signal_3143, signal_1715, signal_3072, signal_1795, signal_4053,
         signal_1015, signal_3365, signal_1016, signal_3146, signal_1714,
         signal_3075, signal_1794, signal_4054, signal_1018, signal_3366,
         signal_1019, signal_3149, signal_1713, signal_3078, signal_1793,
         signal_4055, signal_1021, signal_3367, signal_1022, signal_3152,
         signal_1712, signal_3081, signal_1792, signal_4056, signal_1024,
         signal_3368, signal_1025, signal_3155, signal_1711, signal_3084,
         signal_1791, signal_4057, signal_1027, signal_3369, signal_1028,
         signal_3158, signal_1710, signal_3087, signal_1790, signal_4058,
         signal_1030, signal_3370, signal_1031, signal_3161, signal_1701,
         signal_3090, signal_1781, signal_4059, signal_1033, signal_3371,
         signal_1034, signal_3164, signal_1700, signal_3093, signal_1780,
         signal_4060, signal_1036, signal_3372, signal_1037, signal_3167,
         signal_1699, signal_3096, signal_1779, signal_4061, signal_1039,
         signal_3373, signal_1040, signal_3170, signal_1698, signal_3099,
         signal_1778, signal_4062, signal_1042, signal_3374, signal_1043,
         signal_3173, signal_1697, signal_3102, signal_1777, signal_4063,
         signal_1045, signal_3375, signal_1046, signal_3176, signal_1696,
         signal_3105, signal_1776, signal_4064, signal_1048, signal_3376,
         signal_1049, signal_3179, signal_1695, signal_3108, signal_1775,
         signal_4065, signal_1051, signal_3377, signal_1052, signal_3182,
         signal_1694, signal_3111, signal_1774, signal_4066, signal_1078,
         signal_3378, signal_1079, signal_3138, signal_1741, signal_4067,
         signal_1081, signal_3379, signal_1082, signal_3141, signal_1740,
         signal_4068, signal_1084, signal_3380, signal_1085, signal_3144,
         signal_1739, signal_4069, signal_1087, signal_3381, signal_1088,
         signal_3147, signal_1738, signal_4070, signal_1090, signal_3382,
         signal_1091, signal_3150, signal_1737, signal_4071, signal_1093,
         signal_3383, signal_1094, signal_3153, signal_1736, signal_4072,
         signal_1096, signal_3384, signal_1097, signal_3156, signal_1735,
         signal_4073, signal_1099, signal_3385, signal_1100, signal_3159,
         signal_1734, signal_4074, signal_1102, signal_3386, signal_1103,
         signal_3162, signal_1725, signal_4075, signal_1105, signal_3387,
         signal_1106, signal_3165, signal_1724, signal_4076, signal_1108,
         signal_3388, signal_1109, signal_3168, signal_1723, signal_4077,
         signal_1111, signal_3389, signal_1112, signal_3171, signal_1722,
         signal_4078, signal_1114, signal_3390, signal_1115, signal_3174,
         signal_1721, signal_4079, signal_1117, signal_3391, signal_1118,
         signal_3177, signal_1720, signal_4080, signal_1120, signal_3392,
         signal_1121, signal_3180, signal_1719, signal_4081, signal_1123,
         signal_3393, signal_1124, signal_3183, signal_1718, signal_4082,
         signal_1126, signal_3394, signal_1127, signal_3185, signal_1709,
         signal_4083, signal_1129, signal_3395, signal_1130, signal_3187,
         signal_1708, signal_4084, signal_1132, signal_3396, signal_1133,
         signal_3189, signal_1707, signal_4085, signal_1135, signal_3397,
         signal_1136, signal_3191, signal_1706, signal_4086, signal_1138,
         signal_3398, signal_1139, signal_3193, signal_1705, signal_4087,
         signal_1141, signal_3399, signal_1142, signal_3195, signal_1704,
         signal_4088, signal_1144, signal_3400, signal_1145, signal_3197,
         signal_1703, signal_4089, signal_1147, signal_3401, signal_1148,
         signal_3199, signal_1702, signal_3655, signal_1685, signal_3656,
         signal_1684, signal_3657, signal_1683, signal_3658, signal_1682,
         signal_3659, signal_1681, signal_3660, signal_1680, signal_3661,
         signal_1679, signal_3662, signal_1678, signal_3114, signal_1765,
         signal_3117, signal_1764, signal_3120, signal_1763, signal_3123,
         signal_1762, signal_3126, signal_1761, signal_3129, signal_1760,
         signal_3132, signal_1759, signal_3135, signal_1758, signal_2430,
         signal_1151, signal_2528, signal_1150, signal_2457, signal_1934,
         signal_2433, signal_1153, signal_2529, signal_1152, signal_2459,
         signal_1935, signal_2436, signal_1155, signal_2530, signal_1154,
         signal_2461, signal_1936, signal_2439, signal_1157, signal_3203,
         signal_1156, signal_2533, signal_1937, signal_2452, signal_1942,
         signal_2442, signal_1159, signal_3204, signal_1158, signal_2534,
         signal_1938, signal_2453, signal_1943, signal_2445, signal_1161,
         signal_2531, signal_1160, signal_2464, signal_1939, signal_2448,
         signal_1163, signal_3206, signal_1162, signal_2535, signal_1940,
         signal_2454, signal_1945, signal_2451, signal_1165, signal_2532,
         signal_1164, signal_2466, signal_1941, signal_2468, signal_1946,
         signal_2469, signal_1947, signal_2470, signal_1949, signal_2471,
         signal_1167, signal_2536, signal_1166, signal_2482, signal_1950,
         signal_2472, signal_1169, signal_2537, signal_1168, signal_2483,
         signal_1951, signal_2473, signal_1171, signal_2538, signal_1170,
         signal_2484, signal_1952, signal_2474, signal_1173, signal_3211,
         signal_1172, signal_2541, signal_1953, signal_2479, signal_1184,
         signal_2475, signal_1175, signal_3212, signal_1174, signal_2542,
         signal_1954, signal_2480, signal_1183, signal_2476, signal_1177,
         signal_2539, signal_1176, signal_2485, signal_1955, signal_2477,
         signal_1179, signal_3214, signal_1178, signal_2543, signal_1956,
         signal_2481, signal_1182, signal_2478, signal_1181, signal_2540,
         signal_1180, signal_2486, signal_1957, signal_2487, signal_1958,
         signal_2488, signal_1959, signal_2489, signal_1961, signal_2490,
         signal_1186, signal_2544, signal_1185, signal_2501, signal_1962,
         signal_2491, signal_1188, signal_2545, signal_1187, signal_2502,
         signal_1963, signal_2492, signal_1190, signal_2546, signal_1189,
         signal_2503, signal_1964, signal_2493, signal_1192, signal_3219,
         signal_1191, signal_2549, signal_1965, signal_2498, signal_1203,
         signal_2494, signal_1194, signal_3220, signal_1193, signal_2550,
         signal_1966, signal_2499, signal_1202, signal_2495, signal_1196,
         signal_2547, signal_1195, signal_2504, signal_1967, signal_2496,
         signal_1198, signal_3222, signal_1197, signal_2551, signal_1968,
         signal_2500, signal_1201, signal_2497, signal_1200, signal_2548,
         signal_1199, signal_2505, signal_1969, signal_2506, signal_1970,
         signal_2507, signal_1971, signal_2508, signal_1973, signal_2509,
         signal_1205, signal_2552, signal_1204, signal_2520, signal_1974,
         signal_2510, signal_1207, signal_2553, signal_1206, signal_2521,
         signal_1975, signal_2511, signal_1209, signal_2554, signal_1208,
         signal_2522, signal_1976, signal_2512, signal_1211, signal_3227,
         signal_1210, signal_2557, signal_1977, signal_2517, signal_1222,
         signal_2513, signal_1213, signal_3228, signal_1212, signal_2558,
         signal_1978, signal_2518, signal_1221, signal_2514, signal_1215,
         signal_2555, signal_1214, signal_2523, signal_1979, signal_2515,
         signal_1217, signal_3230, signal_1216, signal_2559, signal_1980,
         signal_2519, signal_1220, signal_2516, signal_1219, signal_2556,
         signal_1218, signal_2524, signal_1981, signal_2525, signal_1225,
         signal_2526, signal_1224, signal_2527, signal_1223, signal_1494,
         signal_1495, signal_1273, signal_1496, signal_1272, signal_1497,
         signal_1498, signal_1499, signal_1500, signal_1501, signal_1269,
         signal_1274, signal_1270, signal_1254, signal_1275, signal_1266,
         signal_1268, signal_1264, signal_1262, signal_1260, signal_1259,
         signal_1258, signal_1256, signal_1271, signal_3232, signal_1517,
         signal_3233, signal_1516, signal_3234, signal_1515, signal_3235,
         signal_1514, signal_3236, signal_1513, signal_3237, signal_1512,
         signal_3238, signal_1511, signal_3239, signal_1510, signal_4640,
         signal_3256, signal_1982, signal_3257, signal_1983, signal_3258,
         signal_1984, signal_3259, signal_1985, signal_3260, signal_1986,
         signal_3261, signal_1987, signal_3402, signal_1988, signal_3403,
         signal_1989, signal_3404, signal_1990, signal_3405, signal_1991,
         signal_3406, signal_1992, signal_3407, signal_1993, signal_3408,
         signal_1994, signal_3409, signal_1995, signal_3410, signal_1996,
         signal_3411, signal_1997, signal_3412, signal_1998, signal_3413,
         signal_1999, signal_3414, signal_2000, signal_3415, signal_2001,
         signal_3416, signal_2002, signal_3417, signal_2003, signal_3418,
         signal_2004, signal_3419, signal_2005, signal_3420, signal_2006,
         signal_3421, signal_2007, signal_3422, signal_2008, signal_3423,
         signal_2009, signal_3424, signal_2010, signal_3425, signal_2011,
         signal_3426, signal_2012, signal_3427, signal_2013, signal_3428,
         signal_2014, signal_3429, signal_2015, signal_3430, signal_2016,
         signal_3431, signal_2017, signal_3432, signal_2018, signal_3433,
         signal_2019, signal_3458, signal_2020, signal_3459, signal_2021,
         signal_3460, signal_2022, signal_3461, signal_2023, signal_3462,
         signal_2024, signal_3463, signal_2025, signal_3464, signal_2026,
         signal_3465, signal_2027, signal_3466, signal_2028, signal_3467,
         signal_2029, signal_3468, signal_2030, signal_3469, signal_2031,
         signal_3470, signal_2032, signal_3471, signal_2033, signal_3472,
         signal_2034, signal_3473, signal_2035, signal_3474, signal_2036,
         signal_3475, signal_2037, signal_3476, signal_2038, signal_3477,
         signal_2039, signal_3478, signal_2040, signal_3479, signal_2041,
         signal_3480, signal_2042, signal_3481, signal_2043, signal_3482,
         signal_2044, signal_3483, signal_2045, signal_3484, signal_2046,
         signal_3485, signal_2047, signal_3486, signal_2048, signal_3487,
         signal_2049, signal_3488, signal_2050, signal_3489, signal_2051,
         signal_3490, signal_2052, signal_3491, signal_2053, signal_3492,
         signal_2054, signal_3493, signal_2055, signal_3494, signal_2056,
         signal_3495, signal_2057, signal_3496, signal_2058, signal_3497,
         signal_2059, signal_3498, signal_2060, signal_3499, signal_2061,
         signal_3500, signal_2062, signal_3501, signal_2063, signal_3502,
         signal_2064, signal_3503, signal_2065, signal_3504, signal_2066,
         signal_3505, signal_2067, signal_3506, signal_2068, signal_3507,
         signal_2069, signal_3508, signal_2070, signal_3509, signal_2071,
         signal_3510, signal_2072, signal_3511, signal_2073, signal_3512,
         signal_2074, signal_3513, signal_2075, signal_3514, signal_2076,
         signal_3515, signal_2077, signal_3516, signal_2078, signal_3517,
         signal_2079, signal_3518, signal_2080, signal_3519, signal_2081,
         signal_3520, signal_2082, signal_3521, signal_2083, signal_3522,
         signal_2084, signal_3523, signal_2085, signal_3524, signal_2086,
         signal_3525, signal_2087, signal_3526, signal_2088, signal_3527,
         signal_2089, signal_3528, signal_2090, signal_3529, signal_2091,
         signal_3530, signal_2092, signal_3531, signal_2093, signal_3532,
         signal_2094, signal_3533, signal_2095, signal_3534, signal_2096,
         signal_3535, signal_2097, signal_3536, signal_2098, signal_3537,
         signal_2099, signal_3538, signal_2100, signal_3539, signal_2101,
         signal_3540, signal_2102, signal_3541, signal_2103, signal_3542,
         signal_2104, signal_3543, signal_2105, signal_3544, signal_2106,
         signal_3545, signal_2107, signal_3546, signal_2108, signal_3547,
         signal_2109, signal_3548, signal_2110, signal_3549, signal_2111,
         signal_3550, signal_2112, signal_3551, signal_2113, signal_3552,
         signal_2114, signal_3553, signal_2115, signal_3554, signal_2116,
         signal_3555, signal_2117, signal_3556, signal_2118, signal_3557,
         signal_2119, signal_3558, signal_2120, signal_3559, signal_2121,
         signal_3560, signal_2122, signal_3561, signal_2123, signal_3562,
         signal_2124, signal_3563, signal_2125, signal_3564, signal_2126,
         signal_3565, signal_2127, signal_3566, signal_2128, signal_3567,
         signal_2129, signal_3568, signal_2130, signal_3569, signal_2131,
         signal_3570, signal_2132, signal_3571, signal_2133, signal_3572,
         signal_2134, signal_3573, signal_2135, signal_3574, signal_2136,
         signal_3575, signal_2137, signal_3576, signal_2138, signal_3577,
         signal_2139, signal_3578, signal_2140, signal_3579, signal_2141,
         signal_3580, signal_2142, signal_3581, signal_2143, signal_3582,
         signal_2144, signal_3583, signal_2145, signal_3584, signal_2146,
         signal_3585, signal_2147, signal_3586, signal_2148, signal_3587,
         signal_2149, signal_3588, signal_2150, signal_3589, signal_2151,
         signal_3590, signal_2152, signal_3663, signal_2153, signal_3664,
         signal_2154, signal_3665, signal_2155, signal_3666, signal_2156,
         signal_3667, signal_2157, signal_3668, signal_2158, signal_3669,
         signal_2159, signal_3670, signal_2160, signal_3671, signal_2161,
         signal_3672, signal_2162, signal_3673, signal_2163, signal_3674,
         signal_2164, signal_3675, signal_2165, signal_3676, signal_2166,
         signal_3677, signal_2167, signal_3678, signal_2168, signal_3679,
         signal_2169, signal_3680, signal_2170, signal_3681, signal_2171,
         signal_3682, signal_2172, signal_3683, signal_2173, signal_3684,
         signal_2174, signal_3685, signal_2175, signal_3686, signal_2176,
         signal_3687, signal_2177, signal_3688, signal_2178, signal_3689,
         signal_2179, signal_3690, signal_2180, signal_3691, signal_2181,
         signal_3692, signal_2182, signal_3693, signal_2183, signal_3694,
         signal_2184, signal_3695, signal_2185, signal_3696, signal_2186,
         signal_3697, signal_2187, signal_3698, signal_2188, signal_3699,
         signal_2189, signal_3700, signal_2190, signal_3701, signal_2191,
         signal_3702, signal_2192, signal_3703, signal_2193, signal_3704,
         signal_2194, signal_3705, signal_2195, signal_3706, signal_2196,
         signal_3707, signal_2197, signal_3708, signal_2198, signal_3709,
         signal_2199, signal_3710, signal_2200, signal_3711, signal_2201,
         signal_3712, signal_2202, signal_3713, signal_2203, signal_3714,
         signal_2204, signal_3715, signal_2205, signal_3716, signal_2206,
         signal_3717, signal_2207, signal_3718, signal_2208, signal_3719,
         signal_2209, signal_3720, signal_2210, signal_3721, signal_2211,
         signal_3722, signal_2212, signal_3723, signal_2213, signal_3724,
         signal_2214, signal_3725, signal_2215, signal_3726, signal_2216,
         signal_3727, signal_2217, signal_3728, signal_2218, signal_3729,
         signal_2219, signal_3730, signal_2220, signal_3731, signal_2221,
         signal_3732, signal_2222, signal_3733, signal_2223, signal_3734,
         signal_2224, signal_3735, signal_2225, signal_3736, signal_2226,
         signal_3737, signal_2227, signal_3738, signal_2228, signal_3739,
         signal_2229, signal_3740, signal_2230, signal_3741, signal_2231,
         signal_3742, signal_2232, signal_3743, signal_2233, signal_3744,
         signal_2234, signal_3745, signal_2235, signal_3746, signal_2236,
         signal_3747, signal_2237, signal_3748, signal_2238, signal_3749,
         signal_2239, signal_3750, signal_2240, signal_3751, signal_2241,
         signal_3752, signal_2242, signal_3753, signal_2243, signal_3754,
         signal_2244, signal_3755, signal_2245, signal_3756, signal_2246,
         signal_3757, signal_2247, signal_3758, signal_2248, signal_3759,
         signal_2249, signal_3760, signal_2250, signal_3761, signal_2251,
         signal_3762, signal_2252, signal_3763, signal_2253, signal_3764,
         signal_2254, signal_3765, signal_2255, signal_3766, signal_2256,
         signal_3767, signal_2257, signal_3768, signal_2258, signal_3769,
         signal_2259, signal_3770, signal_2260, signal_3771, signal_2261,
         signal_3772, signal_2262, signal_3773, signal_2263, signal_3774,
         signal_2264, signal_3775, signal_2265, signal_3776, signal_2266,
         signal_3777, signal_2267, signal_3778, signal_2268, signal_3779,
         signal_2269, signal_3780, signal_2270, signal_3781, signal_2271,
         signal_3782, signal_2272, signal_3783, signal_2273, signal_3784,
         signal_2274, signal_3785, signal_2275, signal_3922, signal_2276,
         signal_3923, signal_2277, signal_3924, signal_2278, signal_3925,
         signal_2279, signal_3926, signal_2280, signal_3927, signal_2281,
         signal_3928, signal_2282, signal_3929, signal_2283, signal_3930,
         signal_2284, signal_3931, signal_2285, signal_3932, signal_2286,
         signal_3933, signal_2287, signal_3934, signal_2288, signal_3935,
         signal_2289, signal_3936, signal_2290, signal_3937, signal_2291,
         signal_3938, signal_2292, signal_3939, signal_2293, signal_3940,
         signal_2294, signal_3941, signal_2295, signal_3942, signal_2296,
         signal_3943, signal_2297, signal_3944, signal_2298, signal_3945,
         signal_2299, signal_3946, signal_2300, signal_3947, signal_2301,
         signal_3948, signal_2302, signal_3949, signal_2303, signal_3950,
         signal_2304, signal_3951, signal_2305, signal_3952, signal_2306,
         signal_3953, signal_2307, signal_3954, signal_2308, signal_3955,
         signal_2309, signal_3956, signal_2310, signal_3957, signal_2311,
         signal_3958, signal_2312, signal_3959, signal_2313, signal_3960,
         signal_2314, signal_3961, signal_2315, signal_3962, signal_2316,
         signal_3963, signal_2317, signal_3964, signal_2318, signal_3965,
         signal_2319, signal_3966, signal_2320, signal_3967, signal_2321,
         signal_3968, signal_2322, signal_3969, signal_2323, signal_3970,
         signal_2324, signal_3971, signal_2325, signal_3972, signal_2326,
         signal_3973, signal_2327, signal_3974, signal_2328, signal_3975,
         signal_2329, signal_3976, signal_2330, signal_3977, signal_2331,
         signal_3978, signal_2332, signal_3979, signal_2333, signal_3980,
         signal_2334, signal_3981, signal_2335, signal_3982, signal_2336,
         signal_3983, signal_2337, signal_3984, signal_2338, signal_3985,
         signal_2339, signal_4090, signal_2340, signal_4091, signal_2341,
         signal_4092, signal_2342, signal_4093, signal_2343, signal_4094,
         signal_2344, signal_4095, signal_2345, signal_4096, signal_2346,
         signal_4097, signal_2347, signal_4098, signal_2348, signal_4099,
         signal_2349, signal_4100, signal_2350, signal_4101, signal_2351,
         signal_4102, signal_2352, signal_4103, signal_2353, signal_4104,
         signal_2354, signal_4105, signal_2355, signal_4106, signal_2356,
         signal_4107, signal_2357, signal_4108, signal_2358, signal_4109,
         signal_2359, signal_4110, signal_2360, signal_4111, signal_2361,
         signal_4112, signal_2362, signal_4113, signal_2363, signal_4114,
         signal_2364, signal_4115, signal_2365, signal_4116, signal_2366,
         signal_4117, signal_2367, signal_4118, signal_2368, signal_4119,
         signal_2369, signal_4120, signal_2370, signal_4121, signal_2371,
         signal_4130, signal_2372, signal_4131, signal_2373, signal_4132,
         signal_2374, signal_4133, signal_2375, signal_4134, signal_2376,
         signal_4135, signal_2377, signal_4136, signal_2378, signal_4137,
         signal_2379, signal_4138, signal_2380, signal_4139, signal_2381,
         signal_4140, signal_2382, signal_4141, signal_2383, signal_4142,
         signal_2384, signal_4143, signal_2385, signal_4144, signal_2386,
         signal_4145, signal_2387, signal_4154, signal_1421, signal_4146,
         signal_1405, signal_4155, signal_1420, signal_4151, signal_1404,
         signal_4156, signal_1419, signal_4148, signal_1403, signal_4157,
         signal_1418, signal_4150, signal_1402, signal_4158, signal_1417,
         signal_4152, signal_1401, signal_4159, signal_1416, signal_4153,
         signal_1400, signal_4160, signal_1415, signal_4147, signal_1399,
         signal_4161, signal_1414, signal_4149, signal_1398, signal_4210,
         signal_705, signal_4187, signal_1557, signal_4211, signal_707,
         signal_4189, signal_1556, signal_4212, signal_709, signal_4191,
         signal_1555, signal_4213, signal_711, signal_4193, signal_1554,
         signal_4214, signal_713, signal_4195, signal_1553, signal_4215,
         signal_715, signal_4197, signal_1552, signal_4216, signal_717,
         signal_4199, signal_1551, signal_4217, signal_719, signal_4201,
         signal_1550, signal_4170, signal_1525, signal_4171, signal_1524,
         signal_4172, signal_1523, signal_4173, signal_1522, signal_4174,
         signal_1521, signal_4175, signal_1520, signal_4176, signal_1519,
         signal_4177, signal_1518, signal_4178, signal_1750, signal_4162,
         signal_724, signal_4179, signal_1751, signal_4163, signal_725,
         signal_4180, signal_1752, signal_4164, signal_726, signal_4181,
         signal_1753, signal_4165, signal_727, signal_4182, signal_1754,
         signal_4166, signal_728, signal_4183, signal_1755, signal_4167,
         signal_729, signal_4184, signal_1756, signal_4168, signal_730,
         signal_4185, signal_1757, signal_4169, signal_731, signal_4218,
         signal_1054, signal_4202, signal_1055, signal_4219, signal_1057,
         signal_4203, signal_1058, signal_4220, signal_1060, signal_4204,
         signal_1061, signal_4221, signal_1063, signal_4205, signal_1064,
         signal_4222, signal_1066, signal_4206, signal_1067, signal_4223,
         signal_1069, signal_4207, signal_1070, signal_4224, signal_1072,
         signal_4208, signal_1073, signal_4225, signal_1075, signal_4209,
         signal_1076, n29, n35, n42, n242, n253, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, cell_2128_n17,
         cell_2128_n34, cell_2128_n33, cell_2128_n32, cell_2128_n31,
         cell_2128_n30, cell_2128_n29, cell_2128_n28, cell_2128_n27,
         cell_2128_n26, cell_2128_n25, cell_2128_n24, cell_2128_n23,
         cell_2128_n22, cell_2128_n21, cell_2128_n20, cell_2128_n19,
         cell_2128_n18, cell_2128_n16, cell_2128_n15, cell_2128_n14,
         cell_2128_n13, cell_2128_n12, cell_2128_n11, cell_2128_n10,
         cell_2128_n9, cell_2128_n8, cell_2128_n7, cell_2128_n6, cell_2128_n5,
         cell_2128_n4, cell_2128_n3, cell_2128_n2, cell_2128_n1,
         cell_2128_LatchedEnable, cell_2128_N19, cell_2128_ShiftRegister_17_,
         cell_1714_a_HPC2_and_n9, cell_1714_a_HPC2_and_n8,
         cell_1714_a_HPC2_and_n7, cell_1714_a_HPC2_and_p_0_out_0__1_,
         cell_1714_a_HPC2_and_p_0_out_1__0_,
         cell_1714_a_HPC2_and_p_1_out_0__1_,
         cell_1714_a_HPC2_and_p_1_out_1__0_,
         cell_1714_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1714_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1714_a_HPC2_and_p_1_in_0__1_, cell_1714_a_HPC2_and_p_1_in_1__0_,
         cell_1714_a_HPC2_and_s_out_0__1_, cell_1714_a_HPC2_and_s_out_1__0_,
         cell_1714_a_HPC2_and_p_0_in_0__1_, cell_1714_a_HPC2_and_p_0_in_1__0_,
         cell_1714_a_HPC2_and_s_in_0__1_, cell_1714_a_HPC2_and_s_in_1__0_,
         cell_1714_a_HPC2_and_z_0__0_, cell_1714_a_HPC2_and_z_1__1_,
         cell_1715_a_HPC2_and_n9, cell_1715_a_HPC2_and_n8,
         cell_1715_a_HPC2_and_n7, cell_1715_a_HPC2_and_p_0_out_0__1_,
         cell_1715_a_HPC2_and_p_0_out_1__0_,
         cell_1715_a_HPC2_and_p_1_out_0__1_,
         cell_1715_a_HPC2_and_p_1_out_1__0_,
         cell_1715_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1715_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1715_a_HPC2_and_p_1_in_0__1_, cell_1715_a_HPC2_and_p_1_in_1__0_,
         cell_1715_a_HPC2_and_s_out_0__1_, cell_1715_a_HPC2_and_s_out_1__0_,
         cell_1715_a_HPC2_and_p_0_in_0__1_, cell_1715_a_HPC2_and_p_0_in_1__0_,
         cell_1715_a_HPC2_and_s_in_0__1_, cell_1715_a_HPC2_and_s_in_1__0_,
         cell_1715_a_HPC2_and_z_0__0_, cell_1715_a_HPC2_and_z_1__1_,
         cell_1716_a_HPC2_and_n9, cell_1716_a_HPC2_and_n8,
         cell_1716_a_HPC2_and_n7, cell_1716_a_HPC2_and_p_0_out_0__1_,
         cell_1716_a_HPC2_and_p_0_out_1__0_,
         cell_1716_a_HPC2_and_p_1_out_0__1_,
         cell_1716_a_HPC2_and_p_1_out_1__0_,
         cell_1716_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1716_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1716_a_HPC2_and_p_1_in_0__1_, cell_1716_a_HPC2_and_p_1_in_1__0_,
         cell_1716_a_HPC2_and_s_out_0__1_, cell_1716_a_HPC2_and_s_out_1__0_,
         cell_1716_a_HPC2_and_p_0_in_0__1_, cell_1716_a_HPC2_and_p_0_in_1__0_,
         cell_1716_a_HPC2_and_s_in_0__1_, cell_1716_a_HPC2_and_s_in_1__0_,
         cell_1716_a_HPC2_and_z_0__0_, cell_1716_a_HPC2_and_z_1__1_,
         cell_1717_a_HPC2_and_n9, cell_1717_a_HPC2_and_n8,
         cell_1717_a_HPC2_and_n7, cell_1717_a_HPC2_and_p_0_out_0__1_,
         cell_1717_a_HPC2_and_p_0_out_1__0_,
         cell_1717_a_HPC2_and_p_1_out_0__1_,
         cell_1717_a_HPC2_and_p_1_out_1__0_,
         cell_1717_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1717_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1717_a_HPC2_and_p_1_in_0__1_, cell_1717_a_HPC2_and_p_1_in_1__0_,
         cell_1717_a_HPC2_and_s_out_0__1_, cell_1717_a_HPC2_and_s_out_1__0_,
         cell_1717_a_HPC2_and_p_0_in_0__1_, cell_1717_a_HPC2_and_p_0_in_1__0_,
         cell_1717_a_HPC2_and_s_in_0__1_, cell_1717_a_HPC2_and_s_in_1__0_,
         cell_1717_a_HPC2_and_z_0__0_, cell_1717_a_HPC2_and_z_1__1_,
         cell_1718_a_HPC2_and_n9, cell_1718_a_HPC2_and_n8,
         cell_1718_a_HPC2_and_n7, cell_1718_a_HPC2_and_p_0_out_0__1_,
         cell_1718_a_HPC2_and_p_0_out_1__0_,
         cell_1718_a_HPC2_and_p_1_out_0__1_,
         cell_1718_a_HPC2_and_p_1_out_1__0_,
         cell_1718_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1718_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1718_a_HPC2_and_p_1_in_0__1_, cell_1718_a_HPC2_and_p_1_in_1__0_,
         cell_1718_a_HPC2_and_s_out_0__1_, cell_1718_a_HPC2_and_s_out_1__0_,
         cell_1718_a_HPC2_and_p_0_in_0__1_, cell_1718_a_HPC2_and_p_0_in_1__0_,
         cell_1718_a_HPC2_and_s_in_0__1_, cell_1718_a_HPC2_and_s_in_1__0_,
         cell_1718_a_HPC2_and_z_0__0_, cell_1718_a_HPC2_and_z_1__1_,
         cell_1719_a_HPC2_and_n9, cell_1719_a_HPC2_and_n8,
         cell_1719_a_HPC2_and_n7, cell_1719_a_HPC2_and_p_0_out_0__1_,
         cell_1719_a_HPC2_and_p_0_out_1__0_,
         cell_1719_a_HPC2_and_p_1_out_0__1_,
         cell_1719_a_HPC2_and_p_1_out_1__0_,
         cell_1719_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1719_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1719_a_HPC2_and_p_1_in_0__1_, cell_1719_a_HPC2_and_p_1_in_1__0_,
         cell_1719_a_HPC2_and_s_out_0__1_, cell_1719_a_HPC2_and_s_out_1__0_,
         cell_1719_a_HPC2_and_p_0_in_0__1_, cell_1719_a_HPC2_and_p_0_in_1__0_,
         cell_1719_a_HPC2_and_s_in_0__1_, cell_1719_a_HPC2_and_s_in_1__0_,
         cell_1719_a_HPC2_and_z_0__0_, cell_1719_a_HPC2_and_z_1__1_,
         cell_1720_a_HPC2_and_n9, cell_1720_a_HPC2_and_n8,
         cell_1720_a_HPC2_and_n7, cell_1720_a_HPC2_and_p_0_out_0__1_,
         cell_1720_a_HPC2_and_p_0_out_1__0_,
         cell_1720_a_HPC2_and_p_1_out_0__1_,
         cell_1720_a_HPC2_and_p_1_out_1__0_,
         cell_1720_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1720_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1720_a_HPC2_and_p_1_in_0__1_, cell_1720_a_HPC2_and_p_1_in_1__0_,
         cell_1720_a_HPC2_and_s_out_0__1_, cell_1720_a_HPC2_and_s_out_1__0_,
         cell_1720_a_HPC2_and_p_0_in_0__1_, cell_1720_a_HPC2_and_p_0_in_1__0_,
         cell_1720_a_HPC2_and_s_in_0__1_, cell_1720_a_HPC2_and_s_in_1__0_,
         cell_1720_a_HPC2_and_z_0__0_, cell_1720_a_HPC2_and_z_1__1_,
         cell_1721_a_HPC2_and_n9, cell_1721_a_HPC2_and_n8,
         cell_1721_a_HPC2_and_n7, cell_1721_a_HPC2_and_p_0_out_0__1_,
         cell_1721_a_HPC2_and_p_0_out_1__0_,
         cell_1721_a_HPC2_and_p_1_out_0__1_,
         cell_1721_a_HPC2_and_p_1_out_1__0_,
         cell_1721_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1721_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1721_a_HPC2_and_p_1_in_0__1_, cell_1721_a_HPC2_and_p_1_in_1__0_,
         cell_1721_a_HPC2_and_s_out_0__1_, cell_1721_a_HPC2_and_s_out_1__0_,
         cell_1721_a_HPC2_and_p_0_in_0__1_, cell_1721_a_HPC2_and_p_0_in_1__0_,
         cell_1721_a_HPC2_and_s_in_0__1_, cell_1721_a_HPC2_and_s_in_1__0_,
         cell_1721_a_HPC2_and_z_0__0_, cell_1721_a_HPC2_and_z_1__1_,
         cell_1722_a_HPC2_and_n9, cell_1722_a_HPC2_and_n8,
         cell_1722_a_HPC2_and_n7, cell_1722_a_HPC2_and_p_0_out_0__1_,
         cell_1722_a_HPC2_and_p_0_out_1__0_,
         cell_1722_a_HPC2_and_p_1_out_0__1_,
         cell_1722_a_HPC2_and_p_1_out_1__0_,
         cell_1722_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1722_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1722_a_HPC2_and_p_1_in_0__1_, cell_1722_a_HPC2_and_p_1_in_1__0_,
         cell_1722_a_HPC2_and_s_out_0__1_, cell_1722_a_HPC2_and_s_out_1__0_,
         cell_1722_a_HPC2_and_p_0_in_0__1_, cell_1722_a_HPC2_and_p_0_in_1__0_,
         cell_1722_a_HPC2_and_s_in_0__1_, cell_1722_a_HPC2_and_s_in_1__0_,
         cell_1722_a_HPC2_and_z_0__0_, cell_1722_a_HPC2_and_z_1__1_,
         cell_1723_a_HPC2_and_n9, cell_1723_a_HPC2_and_n8,
         cell_1723_a_HPC2_and_n7, cell_1723_a_HPC2_and_p_0_out_0__1_,
         cell_1723_a_HPC2_and_p_0_out_1__0_,
         cell_1723_a_HPC2_and_p_1_out_0__1_,
         cell_1723_a_HPC2_and_p_1_out_1__0_,
         cell_1723_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1723_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1723_a_HPC2_and_p_1_in_0__1_, cell_1723_a_HPC2_and_p_1_in_1__0_,
         cell_1723_a_HPC2_and_s_out_0__1_, cell_1723_a_HPC2_and_s_out_1__0_,
         cell_1723_a_HPC2_and_p_0_in_0__1_, cell_1723_a_HPC2_and_p_0_in_1__0_,
         cell_1723_a_HPC2_and_s_in_0__1_, cell_1723_a_HPC2_and_s_in_1__0_,
         cell_1723_a_HPC2_and_z_0__0_, cell_1723_a_HPC2_and_z_1__1_,
         cell_1724_n6, cell_1724_n5, cell_1724_a_HPC2_and_n9,
         cell_1724_a_HPC2_and_n8, cell_1724_a_HPC2_and_n7,
         cell_1724_a_HPC2_and_p_0_out_0__1_,
         cell_1724_a_HPC2_and_p_0_out_1__0_,
         cell_1724_a_HPC2_and_p_1_out_0__1_,
         cell_1724_a_HPC2_and_p_1_out_1__0_,
         cell_1724_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1724_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1724_a_HPC2_and_p_1_in_0__1_, cell_1724_a_HPC2_and_p_1_in_1__0_,
         cell_1724_a_HPC2_and_s_out_0__1_, cell_1724_a_HPC2_and_s_out_1__0_,
         cell_1724_a_HPC2_and_p_0_in_0__1_, cell_1724_a_HPC2_and_p_0_in_1__0_,
         cell_1724_a_HPC2_and_s_in_0__1_, cell_1724_a_HPC2_and_s_in_1__0_,
         cell_1724_a_HPC2_and_z_0__0_, cell_1724_a_HPC2_and_z_1__1_,
         cell_1725_a_HPC2_and_n9, cell_1725_a_HPC2_and_n8,
         cell_1725_a_HPC2_and_n7, cell_1725_a_HPC2_and_p_0_out_0__1_,
         cell_1725_a_HPC2_and_p_0_out_1__0_,
         cell_1725_a_HPC2_and_p_1_out_0__1_,
         cell_1725_a_HPC2_and_p_1_out_1__0_,
         cell_1725_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1725_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1725_a_HPC2_and_p_1_in_0__1_, cell_1725_a_HPC2_and_p_1_in_1__0_,
         cell_1725_a_HPC2_and_s_out_0__1_, cell_1725_a_HPC2_and_s_out_1__0_,
         cell_1725_a_HPC2_and_p_0_in_0__1_, cell_1725_a_HPC2_and_p_0_in_1__0_,
         cell_1725_a_HPC2_and_s_in_0__1_, cell_1725_a_HPC2_and_s_in_1__0_,
         cell_1725_a_HPC2_and_z_0__0_, cell_1725_a_HPC2_and_z_1__1_,
         cell_1726_a_HPC2_and_n9, cell_1726_a_HPC2_and_n8,
         cell_1726_a_HPC2_and_n7, cell_1726_a_HPC2_and_p_0_out_0__1_,
         cell_1726_a_HPC2_and_p_0_out_1__0_,
         cell_1726_a_HPC2_and_p_1_out_0__1_,
         cell_1726_a_HPC2_and_p_1_out_1__0_,
         cell_1726_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1726_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1726_a_HPC2_and_p_1_in_0__1_, cell_1726_a_HPC2_and_p_1_in_1__0_,
         cell_1726_a_HPC2_and_s_out_0__1_, cell_1726_a_HPC2_and_s_out_1__0_,
         cell_1726_a_HPC2_and_p_0_in_0__1_, cell_1726_a_HPC2_and_p_0_in_1__0_,
         cell_1726_a_HPC2_and_s_in_0__1_, cell_1726_a_HPC2_and_s_in_1__0_,
         cell_1726_a_HPC2_and_z_0__0_, cell_1726_a_HPC2_and_z_1__1_,
         cell_1727_a_HPC2_and_n9, cell_1727_a_HPC2_and_n8,
         cell_1727_a_HPC2_and_n7, cell_1727_a_HPC2_and_p_0_out_0__1_,
         cell_1727_a_HPC2_and_p_0_out_1__0_,
         cell_1727_a_HPC2_and_p_1_out_0__1_,
         cell_1727_a_HPC2_and_p_1_out_1__0_,
         cell_1727_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1727_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1727_a_HPC2_and_p_1_in_0__1_, cell_1727_a_HPC2_and_p_1_in_1__0_,
         cell_1727_a_HPC2_and_s_out_0__1_, cell_1727_a_HPC2_and_s_out_1__0_,
         cell_1727_a_HPC2_and_p_0_in_0__1_, cell_1727_a_HPC2_and_p_0_in_1__0_,
         cell_1727_a_HPC2_and_s_in_0__1_, cell_1727_a_HPC2_and_s_in_1__0_,
         cell_1727_a_HPC2_and_z_0__0_, cell_1727_a_HPC2_and_z_1__1_,
         cell_1728_a_HPC2_and_n9, cell_1728_a_HPC2_and_n8,
         cell_1728_a_HPC2_and_n7, cell_1728_a_HPC2_and_p_0_out_0__1_,
         cell_1728_a_HPC2_and_p_0_out_1__0_,
         cell_1728_a_HPC2_and_p_1_out_0__1_,
         cell_1728_a_HPC2_and_p_1_out_1__0_,
         cell_1728_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1728_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1728_a_HPC2_and_p_1_in_0__1_, cell_1728_a_HPC2_and_p_1_in_1__0_,
         cell_1728_a_HPC2_and_s_out_0__1_, cell_1728_a_HPC2_and_s_out_1__0_,
         cell_1728_a_HPC2_and_p_0_in_0__1_, cell_1728_a_HPC2_and_p_0_in_1__0_,
         cell_1728_a_HPC2_and_s_in_0__1_, cell_1728_a_HPC2_and_s_in_1__0_,
         cell_1728_a_HPC2_and_z_0__0_, cell_1728_a_HPC2_and_z_1__1_,
         cell_1729_a_HPC2_and_n9, cell_1729_a_HPC2_and_n8,
         cell_1729_a_HPC2_and_n7, cell_1729_a_HPC2_and_p_0_out_0__1_,
         cell_1729_a_HPC2_and_p_0_out_1__0_,
         cell_1729_a_HPC2_and_p_1_out_0__1_,
         cell_1729_a_HPC2_and_p_1_out_1__0_,
         cell_1729_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1729_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1729_a_HPC2_and_p_1_in_0__1_, cell_1729_a_HPC2_and_p_1_in_1__0_,
         cell_1729_a_HPC2_and_s_out_0__1_, cell_1729_a_HPC2_and_s_out_1__0_,
         cell_1729_a_HPC2_and_p_0_in_0__1_, cell_1729_a_HPC2_and_p_0_in_1__0_,
         cell_1729_a_HPC2_and_s_in_0__1_, cell_1729_a_HPC2_and_s_in_1__0_,
         cell_1729_a_HPC2_and_z_0__0_, cell_1729_a_HPC2_and_z_1__1_,
         cell_1730_a_HPC2_and_n9, cell_1730_a_HPC2_and_n8,
         cell_1730_a_HPC2_and_n7, cell_1730_a_HPC2_and_p_0_out_0__1_,
         cell_1730_a_HPC2_and_p_0_out_1__0_,
         cell_1730_a_HPC2_and_p_1_out_0__1_,
         cell_1730_a_HPC2_and_p_1_out_1__0_,
         cell_1730_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1730_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1730_a_HPC2_and_p_1_in_0__1_, cell_1730_a_HPC2_and_p_1_in_1__0_,
         cell_1730_a_HPC2_and_s_out_0__1_, cell_1730_a_HPC2_and_s_out_1__0_,
         cell_1730_a_HPC2_and_p_0_in_0__1_, cell_1730_a_HPC2_and_p_0_in_1__0_,
         cell_1730_a_HPC2_and_s_in_0__1_, cell_1730_a_HPC2_and_s_in_1__0_,
         cell_1730_a_HPC2_and_z_0__0_, cell_1730_a_HPC2_and_z_1__1_,
         cell_1731_a_HPC2_and_n9, cell_1731_a_HPC2_and_n8,
         cell_1731_a_HPC2_and_n7, cell_1731_a_HPC2_and_p_0_out_0__1_,
         cell_1731_a_HPC2_and_p_0_out_1__0_,
         cell_1731_a_HPC2_and_p_1_out_0__1_,
         cell_1731_a_HPC2_and_p_1_out_1__0_,
         cell_1731_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1731_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1731_a_HPC2_and_p_1_in_0__1_, cell_1731_a_HPC2_and_p_1_in_1__0_,
         cell_1731_a_HPC2_and_s_out_0__1_, cell_1731_a_HPC2_and_s_out_1__0_,
         cell_1731_a_HPC2_and_p_0_in_0__1_, cell_1731_a_HPC2_and_p_0_in_1__0_,
         cell_1731_a_HPC2_and_s_in_0__1_, cell_1731_a_HPC2_and_s_in_1__0_,
         cell_1731_a_HPC2_and_z_0__0_, cell_1731_a_HPC2_and_z_1__1_,
         cell_1732_a_HPC2_and_n9, cell_1732_a_HPC2_and_n8,
         cell_1732_a_HPC2_and_n7, cell_1732_a_HPC2_and_p_0_out_0__1_,
         cell_1732_a_HPC2_and_p_0_out_1__0_,
         cell_1732_a_HPC2_and_p_1_out_0__1_,
         cell_1732_a_HPC2_and_p_1_out_1__0_,
         cell_1732_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1732_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1732_a_HPC2_and_p_1_in_0__1_, cell_1732_a_HPC2_and_p_1_in_1__0_,
         cell_1732_a_HPC2_and_s_out_0__1_, cell_1732_a_HPC2_and_s_out_1__0_,
         cell_1732_a_HPC2_and_p_0_in_0__1_, cell_1732_a_HPC2_and_p_0_in_1__0_,
         cell_1732_a_HPC2_and_s_in_0__1_, cell_1732_a_HPC2_and_s_in_1__0_,
         cell_1732_a_HPC2_and_z_0__0_, cell_1732_a_HPC2_and_z_1__1_,
         cell_1733_a_HPC2_and_n9, cell_1733_a_HPC2_and_n8,
         cell_1733_a_HPC2_and_n7, cell_1733_a_HPC2_and_p_0_out_0__1_,
         cell_1733_a_HPC2_and_p_0_out_1__0_,
         cell_1733_a_HPC2_and_p_1_out_0__1_,
         cell_1733_a_HPC2_and_p_1_out_1__0_,
         cell_1733_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1733_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1733_a_HPC2_and_p_1_in_0__1_, cell_1733_a_HPC2_and_p_1_in_1__0_,
         cell_1733_a_HPC2_and_s_out_0__1_, cell_1733_a_HPC2_and_s_out_1__0_,
         cell_1733_a_HPC2_and_p_0_in_0__1_, cell_1733_a_HPC2_and_p_0_in_1__0_,
         cell_1733_a_HPC2_and_s_in_0__1_, cell_1733_a_HPC2_and_s_in_1__0_,
         cell_1733_a_HPC2_and_z_0__0_, cell_1733_a_HPC2_and_z_1__1_,
         cell_1734_a_HPC2_and_n9, cell_1734_a_HPC2_and_n8,
         cell_1734_a_HPC2_and_n7, cell_1734_a_HPC2_and_p_0_out_0__1_,
         cell_1734_a_HPC2_and_p_0_out_1__0_,
         cell_1734_a_HPC2_and_p_1_out_0__1_,
         cell_1734_a_HPC2_and_p_1_out_1__0_,
         cell_1734_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1734_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1734_a_HPC2_and_p_1_in_0__1_, cell_1734_a_HPC2_and_p_1_in_1__0_,
         cell_1734_a_HPC2_and_s_out_0__1_, cell_1734_a_HPC2_and_s_out_1__0_,
         cell_1734_a_HPC2_and_p_0_in_0__1_, cell_1734_a_HPC2_and_p_0_in_1__0_,
         cell_1734_a_HPC2_and_s_in_0__1_, cell_1734_a_HPC2_and_s_in_1__0_,
         cell_1734_a_HPC2_and_z_0__0_, cell_1734_a_HPC2_and_z_1__1_,
         cell_1735_a_HPC2_and_n9, cell_1735_a_HPC2_and_n8,
         cell_1735_a_HPC2_and_n7, cell_1735_a_HPC2_and_p_0_out_0__1_,
         cell_1735_a_HPC2_and_p_0_out_1__0_,
         cell_1735_a_HPC2_and_p_1_out_0__1_,
         cell_1735_a_HPC2_and_p_1_out_1__0_,
         cell_1735_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1735_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1735_a_HPC2_and_p_1_in_0__1_, cell_1735_a_HPC2_and_p_1_in_1__0_,
         cell_1735_a_HPC2_and_s_out_0__1_, cell_1735_a_HPC2_and_s_out_1__0_,
         cell_1735_a_HPC2_and_p_0_in_0__1_, cell_1735_a_HPC2_and_p_0_in_1__0_,
         cell_1735_a_HPC2_and_s_in_0__1_, cell_1735_a_HPC2_and_s_in_1__0_,
         cell_1735_a_HPC2_and_z_0__0_, cell_1735_a_HPC2_and_z_1__1_,
         cell_1736_a_HPC2_and_n9, cell_1736_a_HPC2_and_n8,
         cell_1736_a_HPC2_and_n7, cell_1736_a_HPC2_and_p_0_out_0__1_,
         cell_1736_a_HPC2_and_p_0_out_1__0_,
         cell_1736_a_HPC2_and_p_1_out_0__1_,
         cell_1736_a_HPC2_and_p_1_out_1__0_,
         cell_1736_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1736_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1736_a_HPC2_and_p_1_in_0__1_, cell_1736_a_HPC2_and_p_1_in_1__0_,
         cell_1736_a_HPC2_and_s_out_0__1_, cell_1736_a_HPC2_and_s_out_1__0_,
         cell_1736_a_HPC2_and_p_0_in_0__1_, cell_1736_a_HPC2_and_p_0_in_1__0_,
         cell_1736_a_HPC2_and_s_in_0__1_, cell_1736_a_HPC2_and_s_in_1__0_,
         cell_1736_a_HPC2_and_z_0__0_, cell_1736_a_HPC2_and_z_1__1_,
         cell_1737_a_HPC2_and_n9, cell_1737_a_HPC2_and_n8,
         cell_1737_a_HPC2_and_n7, cell_1737_a_HPC2_and_p_0_out_0__1_,
         cell_1737_a_HPC2_and_p_0_out_1__0_,
         cell_1737_a_HPC2_and_p_1_out_0__1_,
         cell_1737_a_HPC2_and_p_1_out_1__0_,
         cell_1737_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1737_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1737_a_HPC2_and_p_1_in_0__1_, cell_1737_a_HPC2_and_p_1_in_1__0_,
         cell_1737_a_HPC2_and_s_out_0__1_, cell_1737_a_HPC2_and_s_out_1__0_,
         cell_1737_a_HPC2_and_p_0_in_0__1_, cell_1737_a_HPC2_and_p_0_in_1__0_,
         cell_1737_a_HPC2_and_s_in_0__1_, cell_1737_a_HPC2_and_s_in_1__0_,
         cell_1737_a_HPC2_and_z_0__0_, cell_1737_a_HPC2_and_z_1__1_,
         cell_1738_a_HPC2_and_n9, cell_1738_a_HPC2_and_n8,
         cell_1738_a_HPC2_and_n7, cell_1738_a_HPC2_and_p_0_out_0__1_,
         cell_1738_a_HPC2_and_p_0_out_1__0_,
         cell_1738_a_HPC2_and_p_1_out_0__1_,
         cell_1738_a_HPC2_and_p_1_out_1__0_,
         cell_1738_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1738_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1738_a_HPC2_and_p_1_in_0__1_, cell_1738_a_HPC2_and_p_1_in_1__0_,
         cell_1738_a_HPC2_and_s_out_0__1_, cell_1738_a_HPC2_and_s_out_1__0_,
         cell_1738_a_HPC2_and_p_0_in_0__1_, cell_1738_a_HPC2_and_p_0_in_1__0_,
         cell_1738_a_HPC2_and_s_in_0__1_, cell_1738_a_HPC2_and_s_in_1__0_,
         cell_1738_a_HPC2_and_z_0__0_, cell_1738_a_HPC2_and_z_1__1_,
         cell_1739_a_HPC2_and_n9, cell_1739_a_HPC2_and_n8,
         cell_1739_a_HPC2_and_n7, cell_1739_a_HPC2_and_p_0_out_0__1_,
         cell_1739_a_HPC2_and_p_0_out_1__0_,
         cell_1739_a_HPC2_and_p_1_out_0__1_,
         cell_1739_a_HPC2_and_p_1_out_1__0_,
         cell_1739_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1739_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1739_a_HPC2_and_p_1_in_0__1_, cell_1739_a_HPC2_and_p_1_in_1__0_,
         cell_1739_a_HPC2_and_s_out_0__1_, cell_1739_a_HPC2_and_s_out_1__0_,
         cell_1739_a_HPC2_and_p_0_in_0__1_, cell_1739_a_HPC2_and_p_0_in_1__0_,
         cell_1739_a_HPC2_and_s_in_0__1_, cell_1739_a_HPC2_and_s_in_1__0_,
         cell_1739_a_HPC2_and_z_0__0_, cell_1739_a_HPC2_and_z_1__1_,
         cell_1740_a_HPC2_and_n9, cell_1740_a_HPC2_and_n8,
         cell_1740_a_HPC2_and_n7, cell_1740_a_HPC2_and_p_0_out_0__1_,
         cell_1740_a_HPC2_and_p_0_out_1__0_,
         cell_1740_a_HPC2_and_p_1_out_0__1_,
         cell_1740_a_HPC2_and_p_1_out_1__0_,
         cell_1740_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1740_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1740_a_HPC2_and_p_1_in_0__1_, cell_1740_a_HPC2_and_p_1_in_1__0_,
         cell_1740_a_HPC2_and_s_out_0__1_, cell_1740_a_HPC2_and_s_out_1__0_,
         cell_1740_a_HPC2_and_p_0_in_0__1_, cell_1740_a_HPC2_and_p_0_in_1__0_,
         cell_1740_a_HPC2_and_s_in_0__1_, cell_1740_a_HPC2_and_s_in_1__0_,
         cell_1740_a_HPC2_and_z_0__0_, cell_1740_a_HPC2_and_z_1__1_,
         cell_1741_a_HPC2_and_n9, cell_1741_a_HPC2_and_n8,
         cell_1741_a_HPC2_and_n7, cell_1741_a_HPC2_and_p_0_out_0__1_,
         cell_1741_a_HPC2_and_p_0_out_1__0_,
         cell_1741_a_HPC2_and_p_1_out_0__1_,
         cell_1741_a_HPC2_and_p_1_out_1__0_,
         cell_1741_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1741_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1741_a_HPC2_and_p_1_in_0__1_, cell_1741_a_HPC2_and_p_1_in_1__0_,
         cell_1741_a_HPC2_and_s_out_0__1_, cell_1741_a_HPC2_and_s_out_1__0_,
         cell_1741_a_HPC2_and_p_0_in_0__1_, cell_1741_a_HPC2_and_p_0_in_1__0_,
         cell_1741_a_HPC2_and_s_in_0__1_, cell_1741_a_HPC2_and_s_in_1__0_,
         cell_1741_a_HPC2_and_z_0__0_, cell_1741_a_HPC2_and_z_1__1_,
         cell_1742_a_HPC2_and_n9, cell_1742_a_HPC2_and_n8,
         cell_1742_a_HPC2_and_n7, cell_1742_a_HPC2_and_p_0_out_0__1_,
         cell_1742_a_HPC2_and_p_0_out_1__0_,
         cell_1742_a_HPC2_and_p_1_out_0__1_,
         cell_1742_a_HPC2_and_p_1_out_1__0_,
         cell_1742_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1742_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1742_a_HPC2_and_p_1_in_0__1_, cell_1742_a_HPC2_and_p_1_in_1__0_,
         cell_1742_a_HPC2_and_s_out_0__1_, cell_1742_a_HPC2_and_s_out_1__0_,
         cell_1742_a_HPC2_and_p_0_in_0__1_, cell_1742_a_HPC2_and_p_0_in_1__0_,
         cell_1742_a_HPC2_and_s_in_0__1_, cell_1742_a_HPC2_and_s_in_1__0_,
         cell_1742_a_HPC2_and_z_0__0_, cell_1742_a_HPC2_and_z_1__1_,
         cell_1743_a_HPC2_and_n9, cell_1743_a_HPC2_and_n8,
         cell_1743_a_HPC2_and_n7, cell_1743_a_HPC2_and_p_0_out_0__1_,
         cell_1743_a_HPC2_and_p_0_out_1__0_,
         cell_1743_a_HPC2_and_p_1_out_0__1_,
         cell_1743_a_HPC2_and_p_1_out_1__0_,
         cell_1743_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1743_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1743_a_HPC2_and_p_1_in_0__1_, cell_1743_a_HPC2_and_p_1_in_1__0_,
         cell_1743_a_HPC2_and_s_out_0__1_, cell_1743_a_HPC2_and_s_out_1__0_,
         cell_1743_a_HPC2_and_p_0_in_0__1_, cell_1743_a_HPC2_and_p_0_in_1__0_,
         cell_1743_a_HPC2_and_s_in_0__1_, cell_1743_a_HPC2_and_s_in_1__0_,
         cell_1743_a_HPC2_and_z_0__0_, cell_1743_a_HPC2_and_z_1__1_,
         cell_1744_a_HPC2_and_n9, cell_1744_a_HPC2_and_n8,
         cell_1744_a_HPC2_and_n7, cell_1744_a_HPC2_and_p_0_out_0__1_,
         cell_1744_a_HPC2_and_p_0_out_1__0_,
         cell_1744_a_HPC2_and_p_1_out_0__1_,
         cell_1744_a_HPC2_and_p_1_out_1__0_,
         cell_1744_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1744_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1744_a_HPC2_and_p_1_in_0__1_, cell_1744_a_HPC2_and_p_1_in_1__0_,
         cell_1744_a_HPC2_and_s_out_0__1_, cell_1744_a_HPC2_and_s_out_1__0_,
         cell_1744_a_HPC2_and_p_0_in_0__1_, cell_1744_a_HPC2_and_p_0_in_1__0_,
         cell_1744_a_HPC2_and_s_in_0__1_, cell_1744_a_HPC2_and_s_in_1__0_,
         cell_1744_a_HPC2_and_z_0__0_, cell_1744_a_HPC2_and_z_1__1_,
         cell_1745_a_HPC2_and_n9, cell_1745_a_HPC2_and_n8,
         cell_1745_a_HPC2_and_n7, cell_1745_a_HPC2_and_p_0_out_0__1_,
         cell_1745_a_HPC2_and_p_0_out_1__0_,
         cell_1745_a_HPC2_and_p_1_out_0__1_,
         cell_1745_a_HPC2_and_p_1_out_1__0_,
         cell_1745_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1745_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1745_a_HPC2_and_p_1_in_0__1_, cell_1745_a_HPC2_and_p_1_in_1__0_,
         cell_1745_a_HPC2_and_s_out_0__1_, cell_1745_a_HPC2_and_s_out_1__0_,
         cell_1745_a_HPC2_and_p_0_in_0__1_, cell_1745_a_HPC2_and_p_0_in_1__0_,
         cell_1745_a_HPC2_and_s_in_0__1_, cell_1745_a_HPC2_and_s_in_1__0_,
         cell_1745_a_HPC2_and_z_0__0_, cell_1745_a_HPC2_and_z_1__1_,
         cell_1746_a_HPC2_and_n9, cell_1746_a_HPC2_and_n8,
         cell_1746_a_HPC2_and_n7, cell_1746_a_HPC2_and_p_0_out_0__1_,
         cell_1746_a_HPC2_and_p_0_out_1__0_,
         cell_1746_a_HPC2_and_p_1_out_0__1_,
         cell_1746_a_HPC2_and_p_1_out_1__0_,
         cell_1746_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1746_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1746_a_HPC2_and_p_1_in_0__1_, cell_1746_a_HPC2_and_p_1_in_1__0_,
         cell_1746_a_HPC2_and_s_out_0__1_, cell_1746_a_HPC2_and_s_out_1__0_,
         cell_1746_a_HPC2_and_p_0_in_0__1_, cell_1746_a_HPC2_and_p_0_in_1__0_,
         cell_1746_a_HPC2_and_s_in_0__1_, cell_1746_a_HPC2_and_s_in_1__0_,
         cell_1746_a_HPC2_and_z_0__0_, cell_1746_a_HPC2_and_z_1__1_,
         cell_1747_a_HPC2_and_n9, cell_1747_a_HPC2_and_n8,
         cell_1747_a_HPC2_and_n7, cell_1747_a_HPC2_and_p_0_out_0__1_,
         cell_1747_a_HPC2_and_p_0_out_1__0_,
         cell_1747_a_HPC2_and_p_1_out_0__1_,
         cell_1747_a_HPC2_and_p_1_out_1__0_,
         cell_1747_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1747_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1747_a_HPC2_and_p_1_in_0__1_, cell_1747_a_HPC2_and_p_1_in_1__0_,
         cell_1747_a_HPC2_and_s_out_0__1_, cell_1747_a_HPC2_and_s_out_1__0_,
         cell_1747_a_HPC2_and_p_0_in_0__1_, cell_1747_a_HPC2_and_p_0_in_1__0_,
         cell_1747_a_HPC2_and_s_in_0__1_, cell_1747_a_HPC2_and_s_in_1__0_,
         cell_1747_a_HPC2_and_z_0__0_, cell_1747_a_HPC2_and_z_1__1_,
         cell_1748_a_HPC2_and_n9, cell_1748_a_HPC2_and_n8,
         cell_1748_a_HPC2_and_n7, cell_1748_a_HPC2_and_p_0_out_0__1_,
         cell_1748_a_HPC2_and_p_0_out_1__0_,
         cell_1748_a_HPC2_and_p_1_out_0__1_,
         cell_1748_a_HPC2_and_p_1_out_1__0_,
         cell_1748_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1748_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1748_a_HPC2_and_p_1_in_0__1_, cell_1748_a_HPC2_and_p_1_in_1__0_,
         cell_1748_a_HPC2_and_s_out_0__1_, cell_1748_a_HPC2_and_s_out_1__0_,
         cell_1748_a_HPC2_and_p_0_in_0__1_, cell_1748_a_HPC2_and_p_0_in_1__0_,
         cell_1748_a_HPC2_and_s_in_0__1_, cell_1748_a_HPC2_and_s_in_1__0_,
         cell_1748_a_HPC2_and_z_0__0_, cell_1748_a_HPC2_and_z_1__1_,
         cell_1749_a_HPC2_and_n9, cell_1749_a_HPC2_and_n8,
         cell_1749_a_HPC2_and_n7, cell_1749_a_HPC2_and_p_0_out_0__1_,
         cell_1749_a_HPC2_and_p_0_out_1__0_,
         cell_1749_a_HPC2_and_p_1_out_0__1_,
         cell_1749_a_HPC2_and_p_1_out_1__0_,
         cell_1749_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1749_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1749_a_HPC2_and_p_1_in_0__1_, cell_1749_a_HPC2_and_p_1_in_1__0_,
         cell_1749_a_HPC2_and_s_out_0__1_, cell_1749_a_HPC2_and_s_out_1__0_,
         cell_1749_a_HPC2_and_p_0_in_0__1_, cell_1749_a_HPC2_and_p_0_in_1__0_,
         cell_1749_a_HPC2_and_s_in_0__1_, cell_1749_a_HPC2_and_s_in_1__0_,
         cell_1749_a_HPC2_and_z_0__0_, cell_1749_a_HPC2_and_z_1__1_,
         cell_1750_a_HPC2_and_n9, cell_1750_a_HPC2_and_n8,
         cell_1750_a_HPC2_and_n7, cell_1750_a_HPC2_and_p_0_out_0__1_,
         cell_1750_a_HPC2_and_p_0_out_1__0_,
         cell_1750_a_HPC2_and_p_1_out_0__1_,
         cell_1750_a_HPC2_and_p_1_out_1__0_,
         cell_1750_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1750_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1750_a_HPC2_and_p_1_in_0__1_, cell_1750_a_HPC2_and_p_1_in_1__0_,
         cell_1750_a_HPC2_and_s_out_0__1_, cell_1750_a_HPC2_and_s_out_1__0_,
         cell_1750_a_HPC2_and_p_0_in_0__1_, cell_1750_a_HPC2_and_p_0_in_1__0_,
         cell_1750_a_HPC2_and_s_in_0__1_, cell_1750_a_HPC2_and_s_in_1__0_,
         cell_1750_a_HPC2_and_z_0__0_, cell_1750_a_HPC2_and_z_1__1_,
         cell_1751_a_HPC2_and_n9, cell_1751_a_HPC2_and_n8,
         cell_1751_a_HPC2_and_n7, cell_1751_a_HPC2_and_p_0_out_0__1_,
         cell_1751_a_HPC2_and_p_0_out_1__0_,
         cell_1751_a_HPC2_and_p_1_out_0__1_,
         cell_1751_a_HPC2_and_p_1_out_1__0_,
         cell_1751_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1751_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1751_a_HPC2_and_p_1_in_0__1_, cell_1751_a_HPC2_and_p_1_in_1__0_,
         cell_1751_a_HPC2_and_s_out_0__1_, cell_1751_a_HPC2_and_s_out_1__0_,
         cell_1751_a_HPC2_and_p_0_in_0__1_, cell_1751_a_HPC2_and_p_0_in_1__0_,
         cell_1751_a_HPC2_and_s_in_0__1_, cell_1751_a_HPC2_and_s_in_1__0_,
         cell_1751_a_HPC2_and_z_0__0_, cell_1751_a_HPC2_and_z_1__1_,
         cell_1752_a_HPC2_and_n9, cell_1752_a_HPC2_and_n8,
         cell_1752_a_HPC2_and_n7, cell_1752_a_HPC2_and_p_0_out_0__1_,
         cell_1752_a_HPC2_and_p_0_out_1__0_,
         cell_1752_a_HPC2_and_p_1_out_0__1_,
         cell_1752_a_HPC2_and_p_1_out_1__0_,
         cell_1752_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1752_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1752_a_HPC2_and_p_1_in_0__1_, cell_1752_a_HPC2_and_p_1_in_1__0_,
         cell_1752_a_HPC2_and_s_out_0__1_, cell_1752_a_HPC2_and_s_out_1__0_,
         cell_1752_a_HPC2_and_p_0_in_0__1_, cell_1752_a_HPC2_and_p_0_in_1__0_,
         cell_1752_a_HPC2_and_s_in_0__1_, cell_1752_a_HPC2_and_s_in_1__0_,
         cell_1752_a_HPC2_and_z_0__0_, cell_1752_a_HPC2_and_z_1__1_,
         cell_1753_a_HPC2_and_n9, cell_1753_a_HPC2_and_n8,
         cell_1753_a_HPC2_and_n7, cell_1753_a_HPC2_and_p_0_out_0__1_,
         cell_1753_a_HPC2_and_p_0_out_1__0_,
         cell_1753_a_HPC2_and_p_1_out_0__1_,
         cell_1753_a_HPC2_and_p_1_out_1__0_,
         cell_1753_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1753_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1753_a_HPC2_and_p_1_in_0__1_, cell_1753_a_HPC2_and_p_1_in_1__0_,
         cell_1753_a_HPC2_and_s_out_0__1_, cell_1753_a_HPC2_and_s_out_1__0_,
         cell_1753_a_HPC2_and_p_0_in_0__1_, cell_1753_a_HPC2_and_p_0_in_1__0_,
         cell_1753_a_HPC2_and_s_in_0__1_, cell_1753_a_HPC2_and_s_in_1__0_,
         cell_1753_a_HPC2_and_z_0__0_, cell_1753_a_HPC2_and_z_1__1_,
         cell_1754_a_HPC2_and_n9, cell_1754_a_HPC2_and_n8,
         cell_1754_a_HPC2_and_n7, cell_1754_a_HPC2_and_p_0_out_0__1_,
         cell_1754_a_HPC2_and_p_0_out_1__0_,
         cell_1754_a_HPC2_and_p_1_out_0__1_,
         cell_1754_a_HPC2_and_p_1_out_1__0_,
         cell_1754_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1754_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1754_a_HPC2_and_p_1_in_0__1_, cell_1754_a_HPC2_and_p_1_in_1__0_,
         cell_1754_a_HPC2_and_s_out_0__1_, cell_1754_a_HPC2_and_s_out_1__0_,
         cell_1754_a_HPC2_and_p_0_in_0__1_, cell_1754_a_HPC2_and_p_0_in_1__0_,
         cell_1754_a_HPC2_and_s_in_0__1_, cell_1754_a_HPC2_and_s_in_1__0_,
         cell_1754_a_HPC2_and_z_0__0_, cell_1754_a_HPC2_and_z_1__1_,
         cell_1755_a_HPC2_and_n9, cell_1755_a_HPC2_and_n8,
         cell_1755_a_HPC2_and_n7, cell_1755_a_HPC2_and_p_0_out_0__1_,
         cell_1755_a_HPC2_and_p_0_out_1__0_,
         cell_1755_a_HPC2_and_p_1_out_0__1_,
         cell_1755_a_HPC2_and_p_1_out_1__0_,
         cell_1755_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1755_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1755_a_HPC2_and_p_1_in_0__1_, cell_1755_a_HPC2_and_p_1_in_1__0_,
         cell_1755_a_HPC2_and_s_out_0__1_, cell_1755_a_HPC2_and_s_out_1__0_,
         cell_1755_a_HPC2_and_p_0_in_0__1_, cell_1755_a_HPC2_and_p_0_in_1__0_,
         cell_1755_a_HPC2_and_s_in_0__1_, cell_1755_a_HPC2_and_s_in_1__0_,
         cell_1755_a_HPC2_and_z_0__0_, cell_1755_a_HPC2_and_z_1__1_,
         cell_1756_a_HPC2_and_n9, cell_1756_a_HPC2_and_n8,
         cell_1756_a_HPC2_and_n7, cell_1756_a_HPC2_and_p_0_out_0__1_,
         cell_1756_a_HPC2_and_p_0_out_1__0_,
         cell_1756_a_HPC2_and_p_1_out_0__1_,
         cell_1756_a_HPC2_and_p_1_out_1__0_,
         cell_1756_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1756_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1756_a_HPC2_and_p_1_in_0__1_, cell_1756_a_HPC2_and_p_1_in_1__0_,
         cell_1756_a_HPC2_and_s_out_0__1_, cell_1756_a_HPC2_and_s_out_1__0_,
         cell_1756_a_HPC2_and_p_0_in_0__1_, cell_1756_a_HPC2_and_p_0_in_1__0_,
         cell_1756_a_HPC2_and_s_in_0__1_, cell_1756_a_HPC2_and_s_in_1__0_,
         cell_1756_a_HPC2_and_z_0__0_, cell_1756_a_HPC2_and_z_1__1_,
         cell_1757_a_HPC2_and_n9, cell_1757_a_HPC2_and_n8,
         cell_1757_a_HPC2_and_n7, cell_1757_a_HPC2_and_p_0_out_0__1_,
         cell_1757_a_HPC2_and_p_0_out_1__0_,
         cell_1757_a_HPC2_and_p_1_out_0__1_,
         cell_1757_a_HPC2_and_p_1_out_1__0_,
         cell_1757_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1757_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1757_a_HPC2_and_p_1_in_0__1_, cell_1757_a_HPC2_and_p_1_in_1__0_,
         cell_1757_a_HPC2_and_s_out_0__1_, cell_1757_a_HPC2_and_s_out_1__0_,
         cell_1757_a_HPC2_and_p_0_in_0__1_, cell_1757_a_HPC2_and_p_0_in_1__0_,
         cell_1757_a_HPC2_and_s_in_0__1_, cell_1757_a_HPC2_and_s_in_1__0_,
         cell_1757_a_HPC2_and_z_0__0_, cell_1757_a_HPC2_and_z_1__1_,
         cell_1758_a_HPC2_and_n9, cell_1758_a_HPC2_and_n8,
         cell_1758_a_HPC2_and_n7, cell_1758_a_HPC2_and_p_0_out_0__1_,
         cell_1758_a_HPC2_and_p_0_out_1__0_,
         cell_1758_a_HPC2_and_p_1_out_0__1_,
         cell_1758_a_HPC2_and_p_1_out_1__0_,
         cell_1758_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1758_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1758_a_HPC2_and_p_1_in_0__1_, cell_1758_a_HPC2_and_p_1_in_1__0_,
         cell_1758_a_HPC2_and_s_out_0__1_, cell_1758_a_HPC2_and_s_out_1__0_,
         cell_1758_a_HPC2_and_p_0_in_0__1_, cell_1758_a_HPC2_and_p_0_in_1__0_,
         cell_1758_a_HPC2_and_s_in_0__1_, cell_1758_a_HPC2_and_s_in_1__0_,
         cell_1758_a_HPC2_and_z_0__0_, cell_1758_a_HPC2_and_z_1__1_,
         cell_1759_a_HPC2_and_n9, cell_1759_a_HPC2_and_n8,
         cell_1759_a_HPC2_and_n7, cell_1759_a_HPC2_and_p_0_out_0__1_,
         cell_1759_a_HPC2_and_p_0_out_1__0_,
         cell_1759_a_HPC2_and_p_1_out_0__1_,
         cell_1759_a_HPC2_and_p_1_out_1__0_,
         cell_1759_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1759_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1759_a_HPC2_and_p_1_in_0__1_, cell_1759_a_HPC2_and_p_1_in_1__0_,
         cell_1759_a_HPC2_and_s_out_0__1_, cell_1759_a_HPC2_and_s_out_1__0_,
         cell_1759_a_HPC2_and_p_0_in_0__1_, cell_1759_a_HPC2_and_p_0_in_1__0_,
         cell_1759_a_HPC2_and_s_in_0__1_, cell_1759_a_HPC2_and_s_in_1__0_,
         cell_1759_a_HPC2_and_z_0__0_, cell_1759_a_HPC2_and_z_1__1_,
         cell_1760_n4, cell_1760_n3, cell_1760_a_HPC2_and_n9,
         cell_1760_a_HPC2_and_n8, cell_1760_a_HPC2_and_n7,
         cell_1760_a_HPC2_and_p_0_out_0__1_,
         cell_1760_a_HPC2_and_p_0_out_1__0_,
         cell_1760_a_HPC2_and_p_1_out_0__1_,
         cell_1760_a_HPC2_and_p_1_out_1__0_,
         cell_1760_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1760_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1760_a_HPC2_and_p_1_in_0__1_, cell_1760_a_HPC2_and_p_1_in_1__0_,
         cell_1760_a_HPC2_and_s_out_0__1_, cell_1760_a_HPC2_and_s_out_1__0_,
         cell_1760_a_HPC2_and_p_0_in_0__1_, cell_1760_a_HPC2_and_p_0_in_1__0_,
         cell_1760_a_HPC2_and_s_in_0__1_, cell_1760_a_HPC2_and_s_in_1__0_,
         cell_1760_a_HPC2_and_z_0__0_, cell_1760_a_HPC2_and_z_1__1_,
         cell_1761_a_HPC2_and_n9, cell_1761_a_HPC2_and_n8,
         cell_1761_a_HPC2_and_n7, cell_1761_a_HPC2_and_p_0_out_0__1_,
         cell_1761_a_HPC2_and_p_0_out_1__0_,
         cell_1761_a_HPC2_and_p_1_out_0__1_,
         cell_1761_a_HPC2_and_p_1_out_1__0_,
         cell_1761_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1761_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1761_a_HPC2_and_p_1_in_0__1_, cell_1761_a_HPC2_and_p_1_in_1__0_,
         cell_1761_a_HPC2_and_s_out_0__1_, cell_1761_a_HPC2_and_s_out_1__0_,
         cell_1761_a_HPC2_and_p_0_in_0__1_, cell_1761_a_HPC2_and_p_0_in_1__0_,
         cell_1761_a_HPC2_and_s_in_0__1_, cell_1761_a_HPC2_and_s_in_1__0_,
         cell_1761_a_HPC2_and_z_0__0_, cell_1761_a_HPC2_and_z_1__1_,
         cell_1762_a_HPC2_and_n9, cell_1762_a_HPC2_and_n8,
         cell_1762_a_HPC2_and_n7, cell_1762_a_HPC2_and_p_0_out_0__1_,
         cell_1762_a_HPC2_and_p_0_out_1__0_,
         cell_1762_a_HPC2_and_p_1_out_0__1_,
         cell_1762_a_HPC2_and_p_1_out_1__0_,
         cell_1762_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1762_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1762_a_HPC2_and_p_1_in_0__1_, cell_1762_a_HPC2_and_p_1_in_1__0_,
         cell_1762_a_HPC2_and_s_out_0__1_, cell_1762_a_HPC2_and_s_out_1__0_,
         cell_1762_a_HPC2_and_p_0_in_0__1_, cell_1762_a_HPC2_and_p_0_in_1__0_,
         cell_1762_a_HPC2_and_s_in_0__1_, cell_1762_a_HPC2_and_s_in_1__0_,
         cell_1762_a_HPC2_and_z_0__0_, cell_1762_a_HPC2_and_z_1__1_,
         cell_1763_a_HPC2_and_n9, cell_1763_a_HPC2_and_n8,
         cell_1763_a_HPC2_and_n7, cell_1763_a_HPC2_and_p_0_out_0__1_,
         cell_1763_a_HPC2_and_p_0_out_1__0_,
         cell_1763_a_HPC2_and_p_1_out_0__1_,
         cell_1763_a_HPC2_and_p_1_out_1__0_,
         cell_1763_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1763_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1763_a_HPC2_and_p_1_in_0__1_, cell_1763_a_HPC2_and_p_1_in_1__0_,
         cell_1763_a_HPC2_and_s_out_0__1_, cell_1763_a_HPC2_and_s_out_1__0_,
         cell_1763_a_HPC2_and_p_0_in_0__1_, cell_1763_a_HPC2_and_p_0_in_1__0_,
         cell_1763_a_HPC2_and_s_in_0__1_, cell_1763_a_HPC2_and_s_in_1__0_,
         cell_1763_a_HPC2_and_z_0__0_, cell_1763_a_HPC2_and_z_1__1_,
         cell_1764_a_HPC2_and_n9, cell_1764_a_HPC2_and_n8,
         cell_1764_a_HPC2_and_n7, cell_1764_a_HPC2_and_p_0_out_0__1_,
         cell_1764_a_HPC2_and_p_0_out_1__0_,
         cell_1764_a_HPC2_and_p_1_out_0__1_,
         cell_1764_a_HPC2_and_p_1_out_1__0_,
         cell_1764_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1764_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1764_a_HPC2_and_p_1_in_0__1_, cell_1764_a_HPC2_and_p_1_in_1__0_,
         cell_1764_a_HPC2_and_s_out_0__1_, cell_1764_a_HPC2_and_s_out_1__0_,
         cell_1764_a_HPC2_and_p_0_in_0__1_, cell_1764_a_HPC2_and_p_0_in_1__0_,
         cell_1764_a_HPC2_and_s_in_0__1_, cell_1764_a_HPC2_and_s_in_1__0_,
         cell_1764_a_HPC2_and_z_0__0_, cell_1764_a_HPC2_and_z_1__1_,
         cell_1765_a_HPC2_and_n9, cell_1765_a_HPC2_and_n8,
         cell_1765_a_HPC2_and_n7, cell_1765_a_HPC2_and_p_0_out_0__1_,
         cell_1765_a_HPC2_and_p_0_out_1__0_,
         cell_1765_a_HPC2_and_p_1_out_0__1_,
         cell_1765_a_HPC2_and_p_1_out_1__0_,
         cell_1765_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1765_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1765_a_HPC2_and_p_1_in_0__1_, cell_1765_a_HPC2_and_p_1_in_1__0_,
         cell_1765_a_HPC2_and_s_out_0__1_, cell_1765_a_HPC2_and_s_out_1__0_,
         cell_1765_a_HPC2_and_p_0_in_0__1_, cell_1765_a_HPC2_and_p_0_in_1__0_,
         cell_1765_a_HPC2_and_s_in_0__1_, cell_1765_a_HPC2_and_s_in_1__0_,
         cell_1765_a_HPC2_and_z_0__0_, cell_1765_a_HPC2_and_z_1__1_,
         cell_1766_a_HPC2_and_n9, cell_1766_a_HPC2_and_n8,
         cell_1766_a_HPC2_and_n7, cell_1766_a_HPC2_and_p_0_out_0__1_,
         cell_1766_a_HPC2_and_p_0_out_1__0_,
         cell_1766_a_HPC2_and_p_1_out_0__1_,
         cell_1766_a_HPC2_and_p_1_out_1__0_,
         cell_1766_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1766_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1766_a_HPC2_and_p_1_in_0__1_, cell_1766_a_HPC2_and_p_1_in_1__0_,
         cell_1766_a_HPC2_and_s_out_0__1_, cell_1766_a_HPC2_and_s_out_1__0_,
         cell_1766_a_HPC2_and_p_0_in_0__1_, cell_1766_a_HPC2_and_p_0_in_1__0_,
         cell_1766_a_HPC2_and_s_in_0__1_, cell_1766_a_HPC2_and_s_in_1__0_,
         cell_1766_a_HPC2_and_z_0__0_, cell_1766_a_HPC2_and_z_1__1_,
         cell_1767_a_HPC2_and_n9, cell_1767_a_HPC2_and_n8,
         cell_1767_a_HPC2_and_n7, cell_1767_a_HPC2_and_p_0_out_0__1_,
         cell_1767_a_HPC2_and_p_0_out_1__0_,
         cell_1767_a_HPC2_and_p_1_out_0__1_,
         cell_1767_a_HPC2_and_p_1_out_1__0_,
         cell_1767_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1767_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1767_a_HPC2_and_p_1_in_0__1_, cell_1767_a_HPC2_and_p_1_in_1__0_,
         cell_1767_a_HPC2_and_s_out_0__1_, cell_1767_a_HPC2_and_s_out_1__0_,
         cell_1767_a_HPC2_and_p_0_in_0__1_, cell_1767_a_HPC2_and_p_0_in_1__0_,
         cell_1767_a_HPC2_and_s_in_0__1_, cell_1767_a_HPC2_and_s_in_1__0_,
         cell_1767_a_HPC2_and_z_0__0_, cell_1767_a_HPC2_and_z_1__1_,
         cell_1768_a_HPC2_and_n9, cell_1768_a_HPC2_and_n8,
         cell_1768_a_HPC2_and_n7, cell_1768_a_HPC2_and_p_0_out_0__1_,
         cell_1768_a_HPC2_and_p_0_out_1__0_,
         cell_1768_a_HPC2_and_p_1_out_0__1_,
         cell_1768_a_HPC2_and_p_1_out_1__0_,
         cell_1768_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1768_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1768_a_HPC2_and_p_1_in_0__1_, cell_1768_a_HPC2_and_p_1_in_1__0_,
         cell_1768_a_HPC2_and_s_out_0__1_, cell_1768_a_HPC2_and_s_out_1__0_,
         cell_1768_a_HPC2_and_p_0_in_0__1_, cell_1768_a_HPC2_and_p_0_in_1__0_,
         cell_1768_a_HPC2_and_s_in_0__1_, cell_1768_a_HPC2_and_s_in_1__0_,
         cell_1768_a_HPC2_and_z_0__0_, cell_1768_a_HPC2_and_z_1__1_,
         cell_1769_a_HPC2_and_n9, cell_1769_a_HPC2_and_n8,
         cell_1769_a_HPC2_and_n7, cell_1769_a_HPC2_and_p_0_out_0__1_,
         cell_1769_a_HPC2_and_p_0_out_1__0_,
         cell_1769_a_HPC2_and_p_1_out_0__1_,
         cell_1769_a_HPC2_and_p_1_out_1__0_,
         cell_1769_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1769_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1769_a_HPC2_and_p_1_in_0__1_, cell_1769_a_HPC2_and_p_1_in_1__0_,
         cell_1769_a_HPC2_and_s_out_0__1_, cell_1769_a_HPC2_and_s_out_1__0_,
         cell_1769_a_HPC2_and_p_0_in_0__1_, cell_1769_a_HPC2_and_p_0_in_1__0_,
         cell_1769_a_HPC2_and_s_in_0__1_, cell_1769_a_HPC2_and_s_in_1__0_,
         cell_1769_a_HPC2_and_z_0__0_, cell_1769_a_HPC2_and_z_1__1_,
         cell_1770_a_HPC2_and_n9, cell_1770_a_HPC2_and_n8,
         cell_1770_a_HPC2_and_n7, cell_1770_a_HPC2_and_p_0_out_0__1_,
         cell_1770_a_HPC2_and_p_0_out_1__0_,
         cell_1770_a_HPC2_and_p_1_out_0__1_,
         cell_1770_a_HPC2_and_p_1_out_1__0_,
         cell_1770_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1770_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1770_a_HPC2_and_p_1_in_0__1_, cell_1770_a_HPC2_and_p_1_in_1__0_,
         cell_1770_a_HPC2_and_s_out_0__1_, cell_1770_a_HPC2_and_s_out_1__0_,
         cell_1770_a_HPC2_and_p_0_in_0__1_, cell_1770_a_HPC2_and_p_0_in_1__0_,
         cell_1770_a_HPC2_and_s_in_0__1_, cell_1770_a_HPC2_and_s_in_1__0_,
         cell_1770_a_HPC2_and_z_0__0_, cell_1770_a_HPC2_and_z_1__1_,
         cell_1771_a_HPC2_and_n9, cell_1771_a_HPC2_and_n8,
         cell_1771_a_HPC2_and_n7, cell_1771_a_HPC2_and_p_0_out_0__1_,
         cell_1771_a_HPC2_and_p_0_out_1__0_,
         cell_1771_a_HPC2_and_p_1_out_0__1_,
         cell_1771_a_HPC2_and_p_1_out_1__0_,
         cell_1771_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1771_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1771_a_HPC2_and_p_1_in_0__1_, cell_1771_a_HPC2_and_p_1_in_1__0_,
         cell_1771_a_HPC2_and_s_out_0__1_, cell_1771_a_HPC2_and_s_out_1__0_,
         cell_1771_a_HPC2_and_p_0_in_0__1_, cell_1771_a_HPC2_and_p_0_in_1__0_,
         cell_1771_a_HPC2_and_s_in_0__1_, cell_1771_a_HPC2_and_s_in_1__0_,
         cell_1771_a_HPC2_and_z_0__0_, cell_1771_a_HPC2_and_z_1__1_,
         cell_1772_a_HPC2_and_n9, cell_1772_a_HPC2_and_n8,
         cell_1772_a_HPC2_and_n7, cell_1772_a_HPC2_and_p_0_out_0__1_,
         cell_1772_a_HPC2_and_p_0_out_1__0_,
         cell_1772_a_HPC2_and_p_1_out_0__1_,
         cell_1772_a_HPC2_and_p_1_out_1__0_,
         cell_1772_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1772_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1772_a_HPC2_and_p_1_in_0__1_, cell_1772_a_HPC2_and_p_1_in_1__0_,
         cell_1772_a_HPC2_and_s_out_0__1_, cell_1772_a_HPC2_and_s_out_1__0_,
         cell_1772_a_HPC2_and_p_0_in_0__1_, cell_1772_a_HPC2_and_p_0_in_1__0_,
         cell_1772_a_HPC2_and_s_in_0__1_, cell_1772_a_HPC2_and_s_in_1__0_,
         cell_1772_a_HPC2_and_z_0__0_, cell_1772_a_HPC2_and_z_1__1_,
         cell_1773_a_HPC2_and_n9, cell_1773_a_HPC2_and_n8,
         cell_1773_a_HPC2_and_n7, cell_1773_a_HPC2_and_p_0_out_0__1_,
         cell_1773_a_HPC2_and_p_0_out_1__0_,
         cell_1773_a_HPC2_and_p_1_out_0__1_,
         cell_1773_a_HPC2_and_p_1_out_1__0_,
         cell_1773_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1773_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1773_a_HPC2_and_p_1_in_0__1_, cell_1773_a_HPC2_and_p_1_in_1__0_,
         cell_1773_a_HPC2_and_s_out_0__1_, cell_1773_a_HPC2_and_s_out_1__0_,
         cell_1773_a_HPC2_and_p_0_in_0__1_, cell_1773_a_HPC2_and_p_0_in_1__0_,
         cell_1773_a_HPC2_and_s_in_0__1_, cell_1773_a_HPC2_and_s_in_1__0_,
         cell_1773_a_HPC2_and_z_0__0_, cell_1773_a_HPC2_and_z_1__1_,
         cell_1774_a_HPC2_and_n9, cell_1774_a_HPC2_and_n8,
         cell_1774_a_HPC2_and_n7, cell_1774_a_HPC2_and_p_0_out_0__1_,
         cell_1774_a_HPC2_and_p_0_out_1__0_,
         cell_1774_a_HPC2_and_p_1_out_0__1_,
         cell_1774_a_HPC2_and_p_1_out_1__0_,
         cell_1774_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1774_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1774_a_HPC2_and_p_1_in_0__1_, cell_1774_a_HPC2_and_p_1_in_1__0_,
         cell_1774_a_HPC2_and_s_out_0__1_, cell_1774_a_HPC2_and_s_out_1__0_,
         cell_1774_a_HPC2_and_p_0_in_0__1_, cell_1774_a_HPC2_and_p_0_in_1__0_,
         cell_1774_a_HPC2_and_s_in_0__1_, cell_1774_a_HPC2_and_s_in_1__0_,
         cell_1774_a_HPC2_and_z_0__0_, cell_1774_a_HPC2_and_z_1__1_,
         cell_1775_a_HPC2_and_n9, cell_1775_a_HPC2_and_n8,
         cell_1775_a_HPC2_and_n7, cell_1775_a_HPC2_and_p_0_out_0__1_,
         cell_1775_a_HPC2_and_p_0_out_1__0_,
         cell_1775_a_HPC2_and_p_1_out_0__1_,
         cell_1775_a_HPC2_and_p_1_out_1__0_,
         cell_1775_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1775_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1775_a_HPC2_and_p_1_in_0__1_, cell_1775_a_HPC2_and_p_1_in_1__0_,
         cell_1775_a_HPC2_and_s_out_0__1_, cell_1775_a_HPC2_and_s_out_1__0_,
         cell_1775_a_HPC2_and_p_0_in_0__1_, cell_1775_a_HPC2_and_p_0_in_1__0_,
         cell_1775_a_HPC2_and_s_in_0__1_, cell_1775_a_HPC2_and_s_in_1__0_,
         cell_1775_a_HPC2_and_z_0__0_, cell_1775_a_HPC2_and_z_1__1_,
         cell_1776_a_HPC2_and_n9, cell_1776_a_HPC2_and_n8,
         cell_1776_a_HPC2_and_n7, cell_1776_a_HPC2_and_p_0_out_0__1_,
         cell_1776_a_HPC2_and_p_0_out_1__0_,
         cell_1776_a_HPC2_and_p_1_out_0__1_,
         cell_1776_a_HPC2_and_p_1_out_1__0_,
         cell_1776_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1776_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1776_a_HPC2_and_p_1_in_0__1_, cell_1776_a_HPC2_and_p_1_in_1__0_,
         cell_1776_a_HPC2_and_s_out_0__1_, cell_1776_a_HPC2_and_s_out_1__0_,
         cell_1776_a_HPC2_and_p_0_in_0__1_, cell_1776_a_HPC2_and_p_0_in_1__0_,
         cell_1776_a_HPC2_and_s_in_0__1_, cell_1776_a_HPC2_and_s_in_1__0_,
         cell_1776_a_HPC2_and_z_0__0_, cell_1776_a_HPC2_and_z_1__1_,
         cell_1777_a_HPC2_and_n9, cell_1777_a_HPC2_and_n8,
         cell_1777_a_HPC2_and_n7, cell_1777_a_HPC2_and_p_0_out_0__1_,
         cell_1777_a_HPC2_and_p_0_out_1__0_,
         cell_1777_a_HPC2_and_p_1_out_0__1_,
         cell_1777_a_HPC2_and_p_1_out_1__0_,
         cell_1777_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1777_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1777_a_HPC2_and_p_1_in_0__1_, cell_1777_a_HPC2_and_p_1_in_1__0_,
         cell_1777_a_HPC2_and_s_out_0__1_, cell_1777_a_HPC2_and_s_out_1__0_,
         cell_1777_a_HPC2_and_p_0_in_0__1_, cell_1777_a_HPC2_and_p_0_in_1__0_,
         cell_1777_a_HPC2_and_s_in_0__1_, cell_1777_a_HPC2_and_s_in_1__0_,
         cell_1777_a_HPC2_and_z_0__0_, cell_1777_a_HPC2_and_z_1__1_,
         cell_1778_a_HPC2_and_n9, cell_1778_a_HPC2_and_n8,
         cell_1778_a_HPC2_and_n7, cell_1778_a_HPC2_and_p_0_out_0__1_,
         cell_1778_a_HPC2_and_p_0_out_1__0_,
         cell_1778_a_HPC2_and_p_1_out_0__1_,
         cell_1778_a_HPC2_and_p_1_out_1__0_,
         cell_1778_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1778_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1778_a_HPC2_and_p_1_in_0__1_, cell_1778_a_HPC2_and_p_1_in_1__0_,
         cell_1778_a_HPC2_and_s_out_0__1_, cell_1778_a_HPC2_and_s_out_1__0_,
         cell_1778_a_HPC2_and_p_0_in_0__1_, cell_1778_a_HPC2_and_p_0_in_1__0_,
         cell_1778_a_HPC2_and_s_in_0__1_, cell_1778_a_HPC2_and_s_in_1__0_,
         cell_1778_a_HPC2_and_z_0__0_, cell_1778_a_HPC2_and_z_1__1_,
         cell_1779_a_HPC2_and_n9, cell_1779_a_HPC2_and_n8,
         cell_1779_a_HPC2_and_n7, cell_1779_a_HPC2_and_p_0_out_0__1_,
         cell_1779_a_HPC2_and_p_0_out_1__0_,
         cell_1779_a_HPC2_and_p_1_out_0__1_,
         cell_1779_a_HPC2_and_p_1_out_1__0_,
         cell_1779_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1779_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1779_a_HPC2_and_p_1_in_0__1_, cell_1779_a_HPC2_and_p_1_in_1__0_,
         cell_1779_a_HPC2_and_s_out_0__1_, cell_1779_a_HPC2_and_s_out_1__0_,
         cell_1779_a_HPC2_and_p_0_in_0__1_, cell_1779_a_HPC2_and_p_0_in_1__0_,
         cell_1779_a_HPC2_and_s_in_0__1_, cell_1779_a_HPC2_and_s_in_1__0_,
         cell_1779_a_HPC2_and_z_0__0_, cell_1779_a_HPC2_and_z_1__1_,
         cell_1780_a_HPC2_and_n9, cell_1780_a_HPC2_and_n8,
         cell_1780_a_HPC2_and_n7, cell_1780_a_HPC2_and_p_0_out_0__1_,
         cell_1780_a_HPC2_and_p_0_out_1__0_,
         cell_1780_a_HPC2_and_p_1_out_0__1_,
         cell_1780_a_HPC2_and_p_1_out_1__0_,
         cell_1780_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1780_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1780_a_HPC2_and_p_1_in_0__1_, cell_1780_a_HPC2_and_p_1_in_1__0_,
         cell_1780_a_HPC2_and_s_out_0__1_, cell_1780_a_HPC2_and_s_out_1__0_,
         cell_1780_a_HPC2_and_p_0_in_0__1_, cell_1780_a_HPC2_and_p_0_in_1__0_,
         cell_1780_a_HPC2_and_s_in_0__1_, cell_1780_a_HPC2_and_s_in_1__0_,
         cell_1780_a_HPC2_and_z_0__0_, cell_1780_a_HPC2_and_z_1__1_,
         cell_1781_a_HPC2_and_n9, cell_1781_a_HPC2_and_n8,
         cell_1781_a_HPC2_and_n7, cell_1781_a_HPC2_and_p_0_out_0__1_,
         cell_1781_a_HPC2_and_p_0_out_1__0_,
         cell_1781_a_HPC2_and_p_1_out_0__1_,
         cell_1781_a_HPC2_and_p_1_out_1__0_,
         cell_1781_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1781_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1781_a_HPC2_and_p_1_in_0__1_, cell_1781_a_HPC2_and_p_1_in_1__0_,
         cell_1781_a_HPC2_and_s_out_0__1_, cell_1781_a_HPC2_and_s_out_1__0_,
         cell_1781_a_HPC2_and_p_0_in_0__1_, cell_1781_a_HPC2_and_p_0_in_1__0_,
         cell_1781_a_HPC2_and_s_in_0__1_, cell_1781_a_HPC2_and_s_in_1__0_,
         cell_1781_a_HPC2_and_z_0__0_, cell_1781_a_HPC2_and_z_1__1_,
         cell_1782_a_HPC2_and_n9, cell_1782_a_HPC2_and_n8,
         cell_1782_a_HPC2_and_n7, cell_1782_a_HPC2_and_p_0_out_0__1_,
         cell_1782_a_HPC2_and_p_0_out_1__0_,
         cell_1782_a_HPC2_and_p_1_out_0__1_,
         cell_1782_a_HPC2_and_p_1_out_1__0_,
         cell_1782_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1782_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1782_a_HPC2_and_p_1_in_0__1_, cell_1782_a_HPC2_and_p_1_in_1__0_,
         cell_1782_a_HPC2_and_s_out_0__1_, cell_1782_a_HPC2_and_s_out_1__0_,
         cell_1782_a_HPC2_and_p_0_in_0__1_, cell_1782_a_HPC2_and_p_0_in_1__0_,
         cell_1782_a_HPC2_and_s_in_0__1_, cell_1782_a_HPC2_and_s_in_1__0_,
         cell_1782_a_HPC2_and_z_0__0_, cell_1782_a_HPC2_and_z_1__1_,
         cell_1783_a_HPC2_and_n9, cell_1783_a_HPC2_and_n8,
         cell_1783_a_HPC2_and_n7, cell_1783_a_HPC2_and_p_0_out_0__1_,
         cell_1783_a_HPC2_and_p_0_out_1__0_,
         cell_1783_a_HPC2_and_p_1_out_0__1_,
         cell_1783_a_HPC2_and_p_1_out_1__0_,
         cell_1783_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1783_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1783_a_HPC2_and_p_1_in_0__1_, cell_1783_a_HPC2_and_p_1_in_1__0_,
         cell_1783_a_HPC2_and_s_out_0__1_, cell_1783_a_HPC2_and_s_out_1__0_,
         cell_1783_a_HPC2_and_p_0_in_0__1_, cell_1783_a_HPC2_and_p_0_in_1__0_,
         cell_1783_a_HPC2_and_s_in_0__1_, cell_1783_a_HPC2_and_s_in_1__0_,
         cell_1783_a_HPC2_and_z_0__0_, cell_1783_a_HPC2_and_z_1__1_,
         cell_1784_a_HPC2_and_n9, cell_1784_a_HPC2_and_n8,
         cell_1784_a_HPC2_and_n7, cell_1784_a_HPC2_and_p_0_out_0__1_,
         cell_1784_a_HPC2_and_p_0_out_1__0_,
         cell_1784_a_HPC2_and_p_1_out_0__1_,
         cell_1784_a_HPC2_and_p_1_out_1__0_,
         cell_1784_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1784_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1784_a_HPC2_and_p_1_in_0__1_, cell_1784_a_HPC2_and_p_1_in_1__0_,
         cell_1784_a_HPC2_and_s_out_0__1_, cell_1784_a_HPC2_and_s_out_1__0_,
         cell_1784_a_HPC2_and_p_0_in_0__1_, cell_1784_a_HPC2_and_p_0_in_1__0_,
         cell_1784_a_HPC2_and_s_in_0__1_, cell_1784_a_HPC2_and_s_in_1__0_,
         cell_1784_a_HPC2_and_z_0__0_, cell_1784_a_HPC2_and_z_1__1_,
         cell_1785_a_HPC2_and_n9, cell_1785_a_HPC2_and_n8,
         cell_1785_a_HPC2_and_n7, cell_1785_a_HPC2_and_p_0_out_0__1_,
         cell_1785_a_HPC2_and_p_0_out_1__0_,
         cell_1785_a_HPC2_and_p_1_out_0__1_,
         cell_1785_a_HPC2_and_p_1_out_1__0_,
         cell_1785_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1785_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1785_a_HPC2_and_p_1_in_0__1_, cell_1785_a_HPC2_and_p_1_in_1__0_,
         cell_1785_a_HPC2_and_s_out_0__1_, cell_1785_a_HPC2_and_s_out_1__0_,
         cell_1785_a_HPC2_and_p_0_in_0__1_, cell_1785_a_HPC2_and_p_0_in_1__0_,
         cell_1785_a_HPC2_and_s_in_0__1_, cell_1785_a_HPC2_and_s_in_1__0_,
         cell_1785_a_HPC2_and_z_0__0_, cell_1785_a_HPC2_and_z_1__1_,
         cell_1786_a_HPC2_and_n9, cell_1786_a_HPC2_and_n8,
         cell_1786_a_HPC2_and_n7, cell_1786_a_HPC2_and_p_0_out_0__1_,
         cell_1786_a_HPC2_and_p_0_out_1__0_,
         cell_1786_a_HPC2_and_p_1_out_0__1_,
         cell_1786_a_HPC2_and_p_1_out_1__0_,
         cell_1786_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1786_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1786_a_HPC2_and_p_1_in_0__1_, cell_1786_a_HPC2_and_p_1_in_1__0_,
         cell_1786_a_HPC2_and_s_out_0__1_, cell_1786_a_HPC2_and_s_out_1__0_,
         cell_1786_a_HPC2_and_p_0_in_0__1_, cell_1786_a_HPC2_and_p_0_in_1__0_,
         cell_1786_a_HPC2_and_s_in_0__1_, cell_1786_a_HPC2_and_s_in_1__0_,
         cell_1786_a_HPC2_and_z_0__0_, cell_1786_a_HPC2_and_z_1__1_,
         cell_1787_a_HPC2_and_n9, cell_1787_a_HPC2_and_n8,
         cell_1787_a_HPC2_and_n7, cell_1787_a_HPC2_and_p_0_out_0__1_,
         cell_1787_a_HPC2_and_p_0_out_1__0_,
         cell_1787_a_HPC2_and_p_1_out_0__1_,
         cell_1787_a_HPC2_and_p_1_out_1__0_,
         cell_1787_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1787_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1787_a_HPC2_and_p_1_in_0__1_, cell_1787_a_HPC2_and_p_1_in_1__0_,
         cell_1787_a_HPC2_and_s_out_0__1_, cell_1787_a_HPC2_and_s_out_1__0_,
         cell_1787_a_HPC2_and_p_0_in_0__1_, cell_1787_a_HPC2_and_p_0_in_1__0_,
         cell_1787_a_HPC2_and_s_in_0__1_, cell_1787_a_HPC2_and_s_in_1__0_,
         cell_1787_a_HPC2_and_z_0__0_, cell_1787_a_HPC2_and_z_1__1_,
         cell_1788_a_HPC2_and_n9, cell_1788_a_HPC2_and_n8,
         cell_1788_a_HPC2_and_n7, cell_1788_a_HPC2_and_p_0_out_0__1_,
         cell_1788_a_HPC2_and_p_0_out_1__0_,
         cell_1788_a_HPC2_and_p_1_out_0__1_,
         cell_1788_a_HPC2_and_p_1_out_1__0_,
         cell_1788_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1788_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1788_a_HPC2_and_p_1_in_0__1_, cell_1788_a_HPC2_and_p_1_in_1__0_,
         cell_1788_a_HPC2_and_s_out_0__1_, cell_1788_a_HPC2_and_s_out_1__0_,
         cell_1788_a_HPC2_and_p_0_in_0__1_, cell_1788_a_HPC2_and_p_0_in_1__0_,
         cell_1788_a_HPC2_and_s_in_0__1_, cell_1788_a_HPC2_and_s_in_1__0_,
         cell_1788_a_HPC2_and_z_0__0_, cell_1788_a_HPC2_and_z_1__1_,
         cell_1789_a_HPC2_and_n9, cell_1789_a_HPC2_and_n8,
         cell_1789_a_HPC2_and_n7, cell_1789_a_HPC2_and_p_0_out_0__1_,
         cell_1789_a_HPC2_and_p_0_out_1__0_,
         cell_1789_a_HPC2_and_p_1_out_0__1_,
         cell_1789_a_HPC2_and_p_1_out_1__0_,
         cell_1789_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1789_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1789_a_HPC2_and_p_1_in_0__1_, cell_1789_a_HPC2_and_p_1_in_1__0_,
         cell_1789_a_HPC2_and_s_out_0__1_, cell_1789_a_HPC2_and_s_out_1__0_,
         cell_1789_a_HPC2_and_p_0_in_0__1_, cell_1789_a_HPC2_and_p_0_in_1__0_,
         cell_1789_a_HPC2_and_s_in_0__1_, cell_1789_a_HPC2_and_s_in_1__0_,
         cell_1789_a_HPC2_and_z_0__0_, cell_1789_a_HPC2_and_z_1__1_,
         cell_1790_a_HPC2_and_n9, cell_1790_a_HPC2_and_n8,
         cell_1790_a_HPC2_and_n7, cell_1790_a_HPC2_and_p_0_out_0__1_,
         cell_1790_a_HPC2_and_p_0_out_1__0_,
         cell_1790_a_HPC2_and_p_1_out_0__1_,
         cell_1790_a_HPC2_and_p_1_out_1__0_,
         cell_1790_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1790_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1790_a_HPC2_and_p_1_in_0__1_, cell_1790_a_HPC2_and_p_1_in_1__0_,
         cell_1790_a_HPC2_and_s_out_0__1_, cell_1790_a_HPC2_and_s_out_1__0_,
         cell_1790_a_HPC2_and_p_0_in_0__1_, cell_1790_a_HPC2_and_p_0_in_1__0_,
         cell_1790_a_HPC2_and_s_in_0__1_, cell_1790_a_HPC2_and_s_in_1__0_,
         cell_1790_a_HPC2_and_z_0__0_, cell_1790_a_HPC2_and_z_1__1_,
         cell_1791_n4, cell_1791_n3, cell_1791_a_HPC2_and_n9,
         cell_1791_a_HPC2_and_n8, cell_1791_a_HPC2_and_n7,
         cell_1791_a_HPC2_and_p_0_out_0__1_,
         cell_1791_a_HPC2_and_p_0_out_1__0_,
         cell_1791_a_HPC2_and_p_1_out_0__1_,
         cell_1791_a_HPC2_and_p_1_out_1__0_,
         cell_1791_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1791_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1791_a_HPC2_and_p_1_in_0__1_, cell_1791_a_HPC2_and_p_1_in_1__0_,
         cell_1791_a_HPC2_and_s_out_0__1_, cell_1791_a_HPC2_and_s_out_1__0_,
         cell_1791_a_HPC2_and_p_0_in_0__1_, cell_1791_a_HPC2_and_p_0_in_1__0_,
         cell_1791_a_HPC2_and_s_in_0__1_, cell_1791_a_HPC2_and_s_in_1__0_,
         cell_1791_a_HPC2_and_z_0__0_, cell_1791_a_HPC2_and_z_1__1_,
         cell_1792_a_HPC2_and_n9, cell_1792_a_HPC2_and_n8,
         cell_1792_a_HPC2_and_n7, cell_1792_a_HPC2_and_p_0_out_0__1_,
         cell_1792_a_HPC2_and_p_0_out_1__0_,
         cell_1792_a_HPC2_and_p_1_out_0__1_,
         cell_1792_a_HPC2_and_p_1_out_1__0_,
         cell_1792_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1792_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1792_a_HPC2_and_p_1_in_0__1_, cell_1792_a_HPC2_and_p_1_in_1__0_,
         cell_1792_a_HPC2_and_s_out_0__1_, cell_1792_a_HPC2_and_s_out_1__0_,
         cell_1792_a_HPC2_and_p_0_in_0__1_, cell_1792_a_HPC2_and_p_0_in_1__0_,
         cell_1792_a_HPC2_and_s_in_0__1_, cell_1792_a_HPC2_and_s_in_1__0_,
         cell_1792_a_HPC2_and_z_0__0_, cell_1792_a_HPC2_and_z_1__1_,
         cell_1793_a_HPC2_and_n9, cell_1793_a_HPC2_and_n8,
         cell_1793_a_HPC2_and_n7, cell_1793_a_HPC2_and_p_0_out_0__1_,
         cell_1793_a_HPC2_and_p_0_out_1__0_,
         cell_1793_a_HPC2_and_p_1_out_0__1_,
         cell_1793_a_HPC2_and_p_1_out_1__0_,
         cell_1793_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1793_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1793_a_HPC2_and_p_1_in_0__1_, cell_1793_a_HPC2_and_p_1_in_1__0_,
         cell_1793_a_HPC2_and_s_out_0__1_, cell_1793_a_HPC2_and_s_out_1__0_,
         cell_1793_a_HPC2_and_p_0_in_0__1_, cell_1793_a_HPC2_and_p_0_in_1__0_,
         cell_1793_a_HPC2_and_s_in_0__1_, cell_1793_a_HPC2_and_s_in_1__0_,
         cell_1793_a_HPC2_and_z_0__0_, cell_1793_a_HPC2_and_z_1__1_,
         cell_1794_a_HPC2_and_n9, cell_1794_a_HPC2_and_n8,
         cell_1794_a_HPC2_and_n7, cell_1794_a_HPC2_and_p_0_out_0__1_,
         cell_1794_a_HPC2_and_p_0_out_1__0_,
         cell_1794_a_HPC2_and_p_1_out_0__1_,
         cell_1794_a_HPC2_and_p_1_out_1__0_,
         cell_1794_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1794_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1794_a_HPC2_and_p_1_in_0__1_, cell_1794_a_HPC2_and_p_1_in_1__0_,
         cell_1794_a_HPC2_and_s_out_0__1_, cell_1794_a_HPC2_and_s_out_1__0_,
         cell_1794_a_HPC2_and_p_0_in_0__1_, cell_1794_a_HPC2_and_p_0_in_1__0_,
         cell_1794_a_HPC2_and_s_in_0__1_, cell_1794_a_HPC2_and_s_in_1__0_,
         cell_1794_a_HPC2_and_z_0__0_, cell_1794_a_HPC2_and_z_1__1_,
         cell_1795_a_HPC2_and_n9, cell_1795_a_HPC2_and_n8,
         cell_1795_a_HPC2_and_n7, cell_1795_a_HPC2_and_p_0_out_0__1_,
         cell_1795_a_HPC2_and_p_0_out_1__0_,
         cell_1795_a_HPC2_and_p_1_out_0__1_,
         cell_1795_a_HPC2_and_p_1_out_1__0_,
         cell_1795_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1795_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1795_a_HPC2_and_p_1_in_0__1_, cell_1795_a_HPC2_and_p_1_in_1__0_,
         cell_1795_a_HPC2_and_s_out_0__1_, cell_1795_a_HPC2_and_s_out_1__0_,
         cell_1795_a_HPC2_and_p_0_in_0__1_, cell_1795_a_HPC2_and_p_0_in_1__0_,
         cell_1795_a_HPC2_and_s_in_0__1_, cell_1795_a_HPC2_and_s_in_1__0_,
         cell_1795_a_HPC2_and_z_0__0_, cell_1795_a_HPC2_and_z_1__1_,
         cell_1796_n4, cell_1796_n3, cell_1796_a_HPC2_and_n9,
         cell_1796_a_HPC2_and_n8, cell_1796_a_HPC2_and_n7,
         cell_1796_a_HPC2_and_p_0_out_0__1_,
         cell_1796_a_HPC2_and_p_0_out_1__0_,
         cell_1796_a_HPC2_and_p_1_out_0__1_,
         cell_1796_a_HPC2_and_p_1_out_1__0_,
         cell_1796_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1796_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1796_a_HPC2_and_p_1_in_0__1_, cell_1796_a_HPC2_and_p_1_in_1__0_,
         cell_1796_a_HPC2_and_s_out_0__1_, cell_1796_a_HPC2_and_s_out_1__0_,
         cell_1796_a_HPC2_and_p_0_in_0__1_, cell_1796_a_HPC2_and_p_0_in_1__0_,
         cell_1796_a_HPC2_and_s_in_0__1_, cell_1796_a_HPC2_and_s_in_1__0_,
         cell_1796_a_HPC2_and_z_0__0_, cell_1796_a_HPC2_and_z_1__1_,
         cell_1797_a_HPC2_and_n9, cell_1797_a_HPC2_and_n8,
         cell_1797_a_HPC2_and_n7, cell_1797_a_HPC2_and_p_0_out_0__1_,
         cell_1797_a_HPC2_and_p_0_out_1__0_,
         cell_1797_a_HPC2_and_p_1_out_0__1_,
         cell_1797_a_HPC2_and_p_1_out_1__0_,
         cell_1797_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1797_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1797_a_HPC2_and_p_1_in_0__1_, cell_1797_a_HPC2_and_p_1_in_1__0_,
         cell_1797_a_HPC2_and_s_out_0__1_, cell_1797_a_HPC2_and_s_out_1__0_,
         cell_1797_a_HPC2_and_p_0_in_0__1_, cell_1797_a_HPC2_and_p_0_in_1__0_,
         cell_1797_a_HPC2_and_s_in_0__1_, cell_1797_a_HPC2_and_s_in_1__0_,
         cell_1797_a_HPC2_and_z_0__0_, cell_1797_a_HPC2_and_z_1__1_,
         cell_1798_a_HPC2_and_n9, cell_1798_a_HPC2_and_n8,
         cell_1798_a_HPC2_and_n7, cell_1798_a_HPC2_and_p_0_out_0__1_,
         cell_1798_a_HPC2_and_p_0_out_1__0_,
         cell_1798_a_HPC2_and_p_1_out_0__1_,
         cell_1798_a_HPC2_and_p_1_out_1__0_,
         cell_1798_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1798_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1798_a_HPC2_and_p_1_in_0__1_, cell_1798_a_HPC2_and_p_1_in_1__0_,
         cell_1798_a_HPC2_and_s_out_0__1_, cell_1798_a_HPC2_and_s_out_1__0_,
         cell_1798_a_HPC2_and_p_0_in_0__1_, cell_1798_a_HPC2_and_p_0_in_1__0_,
         cell_1798_a_HPC2_and_s_in_0__1_, cell_1798_a_HPC2_and_s_in_1__0_,
         cell_1798_a_HPC2_and_z_0__0_, cell_1798_a_HPC2_and_z_1__1_,
         cell_1799_a_HPC2_and_n9, cell_1799_a_HPC2_and_n8,
         cell_1799_a_HPC2_and_n7, cell_1799_a_HPC2_and_p_0_out_0__1_,
         cell_1799_a_HPC2_and_p_0_out_1__0_,
         cell_1799_a_HPC2_and_p_1_out_0__1_,
         cell_1799_a_HPC2_and_p_1_out_1__0_,
         cell_1799_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1799_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1799_a_HPC2_and_p_1_in_0__1_, cell_1799_a_HPC2_and_p_1_in_1__0_,
         cell_1799_a_HPC2_and_s_out_0__1_, cell_1799_a_HPC2_and_s_out_1__0_,
         cell_1799_a_HPC2_and_p_0_in_0__1_, cell_1799_a_HPC2_and_p_0_in_1__0_,
         cell_1799_a_HPC2_and_s_in_0__1_, cell_1799_a_HPC2_and_s_in_1__0_,
         cell_1799_a_HPC2_and_z_0__0_, cell_1799_a_HPC2_and_z_1__1_,
         cell_1800_a_HPC2_and_n9, cell_1800_a_HPC2_and_n8,
         cell_1800_a_HPC2_and_n7, cell_1800_a_HPC2_and_p_0_out_0__1_,
         cell_1800_a_HPC2_and_p_0_out_1__0_,
         cell_1800_a_HPC2_and_p_1_out_0__1_,
         cell_1800_a_HPC2_and_p_1_out_1__0_,
         cell_1800_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1800_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1800_a_HPC2_and_p_1_in_0__1_, cell_1800_a_HPC2_and_p_1_in_1__0_,
         cell_1800_a_HPC2_and_s_out_0__1_, cell_1800_a_HPC2_and_s_out_1__0_,
         cell_1800_a_HPC2_and_p_0_in_0__1_, cell_1800_a_HPC2_and_p_0_in_1__0_,
         cell_1800_a_HPC2_and_s_in_0__1_, cell_1800_a_HPC2_and_s_in_1__0_,
         cell_1800_a_HPC2_and_z_0__0_, cell_1800_a_HPC2_and_z_1__1_,
         cell_1801_a_HPC2_and_n9, cell_1801_a_HPC2_and_n8,
         cell_1801_a_HPC2_and_n7, cell_1801_a_HPC2_and_p_0_out_0__1_,
         cell_1801_a_HPC2_and_p_0_out_1__0_,
         cell_1801_a_HPC2_and_p_1_out_0__1_,
         cell_1801_a_HPC2_and_p_1_out_1__0_,
         cell_1801_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1801_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1801_a_HPC2_and_p_1_in_0__1_, cell_1801_a_HPC2_and_p_1_in_1__0_,
         cell_1801_a_HPC2_and_s_out_0__1_, cell_1801_a_HPC2_and_s_out_1__0_,
         cell_1801_a_HPC2_and_p_0_in_0__1_, cell_1801_a_HPC2_and_p_0_in_1__0_,
         cell_1801_a_HPC2_and_s_in_0__1_, cell_1801_a_HPC2_and_s_in_1__0_,
         cell_1801_a_HPC2_and_z_0__0_, cell_1801_a_HPC2_and_z_1__1_,
         cell_1802_a_HPC2_and_n9, cell_1802_a_HPC2_and_n8,
         cell_1802_a_HPC2_and_n7, cell_1802_a_HPC2_and_p_0_out_0__1_,
         cell_1802_a_HPC2_and_p_0_out_1__0_,
         cell_1802_a_HPC2_and_p_1_out_0__1_,
         cell_1802_a_HPC2_and_p_1_out_1__0_,
         cell_1802_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1802_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1802_a_HPC2_and_p_1_in_0__1_, cell_1802_a_HPC2_and_p_1_in_1__0_,
         cell_1802_a_HPC2_and_s_out_0__1_, cell_1802_a_HPC2_and_s_out_1__0_,
         cell_1802_a_HPC2_and_p_0_in_0__1_, cell_1802_a_HPC2_and_p_0_in_1__0_,
         cell_1802_a_HPC2_and_s_in_0__1_, cell_1802_a_HPC2_and_s_in_1__0_,
         cell_1802_a_HPC2_and_z_0__0_, cell_1802_a_HPC2_and_z_1__1_,
         cell_1803_a_HPC2_and_n9, cell_1803_a_HPC2_and_n8,
         cell_1803_a_HPC2_and_n7, cell_1803_a_HPC2_and_p_0_out_0__1_,
         cell_1803_a_HPC2_and_p_0_out_1__0_,
         cell_1803_a_HPC2_and_p_1_out_0__1_,
         cell_1803_a_HPC2_and_p_1_out_1__0_,
         cell_1803_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1803_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1803_a_HPC2_and_p_1_in_0__1_, cell_1803_a_HPC2_and_p_1_in_1__0_,
         cell_1803_a_HPC2_and_s_out_0__1_, cell_1803_a_HPC2_and_s_out_1__0_,
         cell_1803_a_HPC2_and_p_0_in_0__1_, cell_1803_a_HPC2_and_p_0_in_1__0_,
         cell_1803_a_HPC2_and_s_in_0__1_, cell_1803_a_HPC2_and_s_in_1__0_,
         cell_1803_a_HPC2_and_z_0__0_, cell_1803_a_HPC2_and_z_1__1_,
         cell_1804_a_HPC2_and_n9, cell_1804_a_HPC2_and_n8,
         cell_1804_a_HPC2_and_n7, cell_1804_a_HPC2_and_p_0_out_0__1_,
         cell_1804_a_HPC2_and_p_0_out_1__0_,
         cell_1804_a_HPC2_and_p_1_out_0__1_,
         cell_1804_a_HPC2_and_p_1_out_1__0_,
         cell_1804_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1804_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1804_a_HPC2_and_p_1_in_0__1_, cell_1804_a_HPC2_and_p_1_in_1__0_,
         cell_1804_a_HPC2_and_s_out_0__1_, cell_1804_a_HPC2_and_s_out_1__0_,
         cell_1804_a_HPC2_and_p_0_in_0__1_, cell_1804_a_HPC2_and_p_0_in_1__0_,
         cell_1804_a_HPC2_and_s_in_0__1_, cell_1804_a_HPC2_and_s_in_1__0_,
         cell_1804_a_HPC2_and_z_0__0_, cell_1804_a_HPC2_and_z_1__1_,
         cell_1805_a_HPC2_and_n9, cell_1805_a_HPC2_and_n8,
         cell_1805_a_HPC2_and_n7, cell_1805_a_HPC2_and_p_0_out_0__1_,
         cell_1805_a_HPC2_and_p_0_out_1__0_,
         cell_1805_a_HPC2_and_p_1_out_0__1_,
         cell_1805_a_HPC2_and_p_1_out_1__0_,
         cell_1805_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1805_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1805_a_HPC2_and_p_1_in_0__1_, cell_1805_a_HPC2_and_p_1_in_1__0_,
         cell_1805_a_HPC2_and_s_out_0__1_, cell_1805_a_HPC2_and_s_out_1__0_,
         cell_1805_a_HPC2_and_p_0_in_0__1_, cell_1805_a_HPC2_and_p_0_in_1__0_,
         cell_1805_a_HPC2_and_s_in_0__1_, cell_1805_a_HPC2_and_s_in_1__0_,
         cell_1805_a_HPC2_and_z_0__0_, cell_1805_a_HPC2_and_z_1__1_,
         cell_1806_a_HPC2_and_n9, cell_1806_a_HPC2_and_n8,
         cell_1806_a_HPC2_and_n7, cell_1806_a_HPC2_and_p_0_out_0__1_,
         cell_1806_a_HPC2_and_p_0_out_1__0_,
         cell_1806_a_HPC2_and_p_1_out_0__1_,
         cell_1806_a_HPC2_and_p_1_out_1__0_,
         cell_1806_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1806_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1806_a_HPC2_and_p_1_in_0__1_, cell_1806_a_HPC2_and_p_1_in_1__0_,
         cell_1806_a_HPC2_and_s_out_0__1_, cell_1806_a_HPC2_and_s_out_1__0_,
         cell_1806_a_HPC2_and_p_0_in_0__1_, cell_1806_a_HPC2_and_p_0_in_1__0_,
         cell_1806_a_HPC2_and_s_in_0__1_, cell_1806_a_HPC2_and_s_in_1__0_,
         cell_1806_a_HPC2_and_z_0__0_, cell_1806_a_HPC2_and_z_1__1_,
         cell_1807_n4, cell_1807_n3, cell_1807_a_HPC2_and_n9,
         cell_1807_a_HPC2_and_n8, cell_1807_a_HPC2_and_n7,
         cell_1807_a_HPC2_and_p_0_out_0__1_,
         cell_1807_a_HPC2_and_p_0_out_1__0_,
         cell_1807_a_HPC2_and_p_1_out_0__1_,
         cell_1807_a_HPC2_and_p_1_out_1__0_,
         cell_1807_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1807_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1807_a_HPC2_and_p_1_in_0__1_, cell_1807_a_HPC2_and_p_1_in_1__0_,
         cell_1807_a_HPC2_and_s_out_0__1_, cell_1807_a_HPC2_and_s_out_1__0_,
         cell_1807_a_HPC2_and_p_0_in_0__1_, cell_1807_a_HPC2_and_p_0_in_1__0_,
         cell_1807_a_HPC2_and_s_in_0__1_, cell_1807_a_HPC2_and_s_in_1__0_,
         cell_1807_a_HPC2_and_z_0__0_, cell_1807_a_HPC2_and_z_1__1_,
         cell_1808_a_HPC2_and_n9, cell_1808_a_HPC2_and_n8,
         cell_1808_a_HPC2_and_n7, cell_1808_a_HPC2_and_p_0_out_0__1_,
         cell_1808_a_HPC2_and_p_0_out_1__0_,
         cell_1808_a_HPC2_and_p_1_out_0__1_,
         cell_1808_a_HPC2_and_p_1_out_1__0_,
         cell_1808_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1808_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1808_a_HPC2_and_p_1_in_0__1_, cell_1808_a_HPC2_and_p_1_in_1__0_,
         cell_1808_a_HPC2_and_s_out_0__1_, cell_1808_a_HPC2_and_s_out_1__0_,
         cell_1808_a_HPC2_and_p_0_in_0__1_, cell_1808_a_HPC2_and_p_0_in_1__0_,
         cell_1808_a_HPC2_and_s_in_0__1_, cell_1808_a_HPC2_and_s_in_1__0_,
         cell_1808_a_HPC2_and_z_0__0_, cell_1808_a_HPC2_and_z_1__1_,
         cell_1809_a_HPC2_and_n9, cell_1809_a_HPC2_and_n8,
         cell_1809_a_HPC2_and_n7, cell_1809_a_HPC2_and_p_0_out_0__1_,
         cell_1809_a_HPC2_and_p_0_out_1__0_,
         cell_1809_a_HPC2_and_p_1_out_0__1_,
         cell_1809_a_HPC2_and_p_1_out_1__0_,
         cell_1809_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1809_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1809_a_HPC2_and_p_1_in_0__1_, cell_1809_a_HPC2_and_p_1_in_1__0_,
         cell_1809_a_HPC2_and_s_out_0__1_, cell_1809_a_HPC2_and_s_out_1__0_,
         cell_1809_a_HPC2_and_p_0_in_0__1_, cell_1809_a_HPC2_and_p_0_in_1__0_,
         cell_1809_a_HPC2_and_s_in_0__1_, cell_1809_a_HPC2_and_s_in_1__0_,
         cell_1809_a_HPC2_and_z_0__0_, cell_1809_a_HPC2_and_z_1__1_,
         cell_1810_a_HPC2_and_n9, cell_1810_a_HPC2_and_n8,
         cell_1810_a_HPC2_and_n7, cell_1810_a_HPC2_and_p_0_out_0__1_,
         cell_1810_a_HPC2_and_p_0_out_1__0_,
         cell_1810_a_HPC2_and_p_1_out_0__1_,
         cell_1810_a_HPC2_and_p_1_out_1__0_,
         cell_1810_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1810_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1810_a_HPC2_and_p_1_in_0__1_, cell_1810_a_HPC2_and_p_1_in_1__0_,
         cell_1810_a_HPC2_and_s_out_0__1_, cell_1810_a_HPC2_and_s_out_1__0_,
         cell_1810_a_HPC2_and_p_0_in_0__1_, cell_1810_a_HPC2_and_p_0_in_1__0_,
         cell_1810_a_HPC2_and_s_in_0__1_, cell_1810_a_HPC2_and_s_in_1__0_,
         cell_1810_a_HPC2_and_z_0__0_, cell_1810_a_HPC2_and_z_1__1_,
         cell_1811_a_HPC2_and_n9, cell_1811_a_HPC2_and_n8,
         cell_1811_a_HPC2_and_n7, cell_1811_a_HPC2_and_p_0_out_0__1_,
         cell_1811_a_HPC2_and_p_0_out_1__0_,
         cell_1811_a_HPC2_and_p_1_out_0__1_,
         cell_1811_a_HPC2_and_p_1_out_1__0_,
         cell_1811_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1811_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1811_a_HPC2_and_p_1_in_0__1_, cell_1811_a_HPC2_and_p_1_in_1__0_,
         cell_1811_a_HPC2_and_s_out_0__1_, cell_1811_a_HPC2_and_s_out_1__0_,
         cell_1811_a_HPC2_and_p_0_in_0__1_, cell_1811_a_HPC2_and_p_0_in_1__0_,
         cell_1811_a_HPC2_and_s_in_0__1_, cell_1811_a_HPC2_and_s_in_1__0_,
         cell_1811_a_HPC2_and_z_0__0_, cell_1811_a_HPC2_and_z_1__1_,
         cell_1812_a_HPC2_and_n9, cell_1812_a_HPC2_and_n8,
         cell_1812_a_HPC2_and_n7, cell_1812_a_HPC2_and_p_0_out_0__1_,
         cell_1812_a_HPC2_and_p_0_out_1__0_,
         cell_1812_a_HPC2_and_p_1_out_0__1_,
         cell_1812_a_HPC2_and_p_1_out_1__0_,
         cell_1812_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1812_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1812_a_HPC2_and_p_1_in_0__1_, cell_1812_a_HPC2_and_p_1_in_1__0_,
         cell_1812_a_HPC2_and_s_out_0__1_, cell_1812_a_HPC2_and_s_out_1__0_,
         cell_1812_a_HPC2_and_p_0_in_0__1_, cell_1812_a_HPC2_and_p_0_in_1__0_,
         cell_1812_a_HPC2_and_s_in_0__1_, cell_1812_a_HPC2_and_s_in_1__0_,
         cell_1812_a_HPC2_and_z_0__0_, cell_1812_a_HPC2_and_z_1__1_,
         cell_1813_a_HPC2_and_n9, cell_1813_a_HPC2_and_n8,
         cell_1813_a_HPC2_and_n7, cell_1813_a_HPC2_and_p_0_out_0__1_,
         cell_1813_a_HPC2_and_p_0_out_1__0_,
         cell_1813_a_HPC2_and_p_1_out_0__1_,
         cell_1813_a_HPC2_and_p_1_out_1__0_,
         cell_1813_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1813_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1813_a_HPC2_and_p_1_in_0__1_, cell_1813_a_HPC2_and_p_1_in_1__0_,
         cell_1813_a_HPC2_and_s_out_0__1_, cell_1813_a_HPC2_and_s_out_1__0_,
         cell_1813_a_HPC2_and_p_0_in_0__1_, cell_1813_a_HPC2_and_p_0_in_1__0_,
         cell_1813_a_HPC2_and_s_in_0__1_, cell_1813_a_HPC2_and_s_in_1__0_,
         cell_1813_a_HPC2_and_z_0__0_, cell_1813_a_HPC2_and_z_1__1_,
         cell_1814_a_HPC2_and_n9, cell_1814_a_HPC2_and_n8,
         cell_1814_a_HPC2_and_n7, cell_1814_a_HPC2_and_p_0_out_0__1_,
         cell_1814_a_HPC2_and_p_0_out_1__0_,
         cell_1814_a_HPC2_and_p_1_out_0__1_,
         cell_1814_a_HPC2_and_p_1_out_1__0_,
         cell_1814_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1814_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1814_a_HPC2_and_p_1_in_0__1_, cell_1814_a_HPC2_and_p_1_in_1__0_,
         cell_1814_a_HPC2_and_s_out_0__1_, cell_1814_a_HPC2_and_s_out_1__0_,
         cell_1814_a_HPC2_and_p_0_in_0__1_, cell_1814_a_HPC2_and_p_0_in_1__0_,
         cell_1814_a_HPC2_and_s_in_0__1_, cell_1814_a_HPC2_and_s_in_1__0_,
         cell_1814_a_HPC2_and_z_0__0_, cell_1814_a_HPC2_and_z_1__1_,
         cell_1815_a_HPC2_and_n9, cell_1815_a_HPC2_and_n8,
         cell_1815_a_HPC2_and_n7, cell_1815_a_HPC2_and_p_0_out_0__1_,
         cell_1815_a_HPC2_and_p_0_out_1__0_,
         cell_1815_a_HPC2_and_p_1_out_0__1_,
         cell_1815_a_HPC2_and_p_1_out_1__0_,
         cell_1815_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1815_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1815_a_HPC2_and_p_1_in_0__1_, cell_1815_a_HPC2_and_p_1_in_1__0_,
         cell_1815_a_HPC2_and_s_out_0__1_, cell_1815_a_HPC2_and_s_out_1__0_,
         cell_1815_a_HPC2_and_p_0_in_0__1_, cell_1815_a_HPC2_and_p_0_in_1__0_,
         cell_1815_a_HPC2_and_s_in_0__1_, cell_1815_a_HPC2_and_s_in_1__0_,
         cell_1815_a_HPC2_and_z_0__0_, cell_1815_a_HPC2_and_z_1__1_,
         cell_1816_a_HPC2_and_n9, cell_1816_a_HPC2_and_n8,
         cell_1816_a_HPC2_and_n7, cell_1816_a_HPC2_and_p_0_out_0__1_,
         cell_1816_a_HPC2_and_p_0_out_1__0_,
         cell_1816_a_HPC2_and_p_1_out_0__1_,
         cell_1816_a_HPC2_and_p_1_out_1__0_,
         cell_1816_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1816_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1816_a_HPC2_and_p_1_in_0__1_, cell_1816_a_HPC2_and_p_1_in_1__0_,
         cell_1816_a_HPC2_and_s_out_0__1_, cell_1816_a_HPC2_and_s_out_1__0_,
         cell_1816_a_HPC2_and_p_0_in_0__1_, cell_1816_a_HPC2_and_p_0_in_1__0_,
         cell_1816_a_HPC2_and_s_in_0__1_, cell_1816_a_HPC2_and_s_in_1__0_,
         cell_1816_a_HPC2_and_z_0__0_, cell_1816_a_HPC2_and_z_1__1_,
         cell_1817_a_HPC2_and_n9, cell_1817_a_HPC2_and_n8,
         cell_1817_a_HPC2_and_n7, cell_1817_a_HPC2_and_p_0_out_0__1_,
         cell_1817_a_HPC2_and_p_0_out_1__0_,
         cell_1817_a_HPC2_and_p_1_out_0__1_,
         cell_1817_a_HPC2_and_p_1_out_1__0_,
         cell_1817_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1817_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1817_a_HPC2_and_p_1_in_0__1_, cell_1817_a_HPC2_and_p_1_in_1__0_,
         cell_1817_a_HPC2_and_s_out_0__1_, cell_1817_a_HPC2_and_s_out_1__0_,
         cell_1817_a_HPC2_and_p_0_in_0__1_, cell_1817_a_HPC2_and_p_0_in_1__0_,
         cell_1817_a_HPC2_and_s_in_0__1_, cell_1817_a_HPC2_and_s_in_1__0_,
         cell_1817_a_HPC2_and_z_0__0_, cell_1817_a_HPC2_and_z_1__1_,
         cell_1818_a_HPC2_and_n9, cell_1818_a_HPC2_and_n8,
         cell_1818_a_HPC2_and_n7, cell_1818_a_HPC2_and_p_0_out_0__1_,
         cell_1818_a_HPC2_and_p_0_out_1__0_,
         cell_1818_a_HPC2_and_p_1_out_0__1_,
         cell_1818_a_HPC2_and_p_1_out_1__0_,
         cell_1818_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1818_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1818_a_HPC2_and_p_1_in_0__1_, cell_1818_a_HPC2_and_p_1_in_1__0_,
         cell_1818_a_HPC2_and_s_out_0__1_, cell_1818_a_HPC2_and_s_out_1__0_,
         cell_1818_a_HPC2_and_p_0_in_0__1_, cell_1818_a_HPC2_and_p_0_in_1__0_,
         cell_1818_a_HPC2_and_s_in_0__1_, cell_1818_a_HPC2_and_s_in_1__0_,
         cell_1818_a_HPC2_and_z_0__0_, cell_1818_a_HPC2_and_z_1__1_,
         cell_1819_a_HPC2_and_n9, cell_1819_a_HPC2_and_n8,
         cell_1819_a_HPC2_and_n7, cell_1819_a_HPC2_and_p_0_out_0__1_,
         cell_1819_a_HPC2_and_p_0_out_1__0_,
         cell_1819_a_HPC2_and_p_1_out_0__1_,
         cell_1819_a_HPC2_and_p_1_out_1__0_,
         cell_1819_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1819_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1819_a_HPC2_and_p_1_in_0__1_, cell_1819_a_HPC2_and_p_1_in_1__0_,
         cell_1819_a_HPC2_and_s_out_0__1_, cell_1819_a_HPC2_and_s_out_1__0_,
         cell_1819_a_HPC2_and_p_0_in_0__1_, cell_1819_a_HPC2_and_p_0_in_1__0_,
         cell_1819_a_HPC2_and_s_in_0__1_, cell_1819_a_HPC2_and_s_in_1__0_,
         cell_1819_a_HPC2_and_z_0__0_, cell_1819_a_HPC2_and_z_1__1_,
         cell_1820_a_HPC2_and_n9, cell_1820_a_HPC2_and_n8,
         cell_1820_a_HPC2_and_n7, cell_1820_a_HPC2_and_p_0_out_0__1_,
         cell_1820_a_HPC2_and_p_0_out_1__0_,
         cell_1820_a_HPC2_and_p_1_out_0__1_,
         cell_1820_a_HPC2_and_p_1_out_1__0_,
         cell_1820_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1820_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1820_a_HPC2_and_p_1_in_0__1_, cell_1820_a_HPC2_and_p_1_in_1__0_,
         cell_1820_a_HPC2_and_s_out_0__1_, cell_1820_a_HPC2_and_s_out_1__0_,
         cell_1820_a_HPC2_and_p_0_in_0__1_, cell_1820_a_HPC2_and_p_0_in_1__0_,
         cell_1820_a_HPC2_and_s_in_0__1_, cell_1820_a_HPC2_and_s_in_1__0_,
         cell_1820_a_HPC2_and_z_0__0_, cell_1820_a_HPC2_and_z_1__1_,
         cell_1821_a_HPC2_and_n9, cell_1821_a_HPC2_and_n8,
         cell_1821_a_HPC2_and_n7, cell_1821_a_HPC2_and_p_0_out_0__1_,
         cell_1821_a_HPC2_and_p_0_out_1__0_,
         cell_1821_a_HPC2_and_p_1_out_0__1_,
         cell_1821_a_HPC2_and_p_1_out_1__0_,
         cell_1821_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1821_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1821_a_HPC2_and_p_1_in_0__1_, cell_1821_a_HPC2_and_p_1_in_1__0_,
         cell_1821_a_HPC2_and_s_out_0__1_, cell_1821_a_HPC2_and_s_out_1__0_,
         cell_1821_a_HPC2_and_p_0_in_0__1_, cell_1821_a_HPC2_and_p_0_in_1__0_,
         cell_1821_a_HPC2_and_s_in_0__1_, cell_1821_a_HPC2_and_s_in_1__0_,
         cell_1821_a_HPC2_and_z_0__0_, cell_1821_a_HPC2_and_z_1__1_,
         cell_1822_a_HPC2_and_n9, cell_1822_a_HPC2_and_n8,
         cell_1822_a_HPC2_and_n7, cell_1822_a_HPC2_and_p_0_out_0__1_,
         cell_1822_a_HPC2_and_p_0_out_1__0_,
         cell_1822_a_HPC2_and_p_1_out_0__1_,
         cell_1822_a_HPC2_and_p_1_out_1__0_,
         cell_1822_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1822_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1822_a_HPC2_and_p_1_in_0__1_, cell_1822_a_HPC2_and_p_1_in_1__0_,
         cell_1822_a_HPC2_and_s_out_0__1_, cell_1822_a_HPC2_and_s_out_1__0_,
         cell_1822_a_HPC2_and_p_0_in_0__1_, cell_1822_a_HPC2_and_p_0_in_1__0_,
         cell_1822_a_HPC2_and_s_in_0__1_, cell_1822_a_HPC2_and_s_in_1__0_,
         cell_1822_a_HPC2_and_z_0__0_, cell_1822_a_HPC2_and_z_1__1_,
         cell_1823_a_HPC2_and_n9, cell_1823_a_HPC2_and_n8,
         cell_1823_a_HPC2_and_n7, cell_1823_a_HPC2_and_p_0_out_0__1_,
         cell_1823_a_HPC2_and_p_0_out_1__0_,
         cell_1823_a_HPC2_and_p_1_out_0__1_,
         cell_1823_a_HPC2_and_p_1_out_1__0_,
         cell_1823_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1823_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1823_a_HPC2_and_p_1_in_0__1_, cell_1823_a_HPC2_and_p_1_in_1__0_,
         cell_1823_a_HPC2_and_s_out_0__1_, cell_1823_a_HPC2_and_s_out_1__0_,
         cell_1823_a_HPC2_and_p_0_in_0__1_, cell_1823_a_HPC2_and_p_0_in_1__0_,
         cell_1823_a_HPC2_and_s_in_0__1_, cell_1823_a_HPC2_and_s_in_1__0_,
         cell_1823_a_HPC2_and_z_0__0_, cell_1823_a_HPC2_and_z_1__1_,
         cell_1824_n4, cell_1824_n3, cell_1824_a_HPC2_and_n9,
         cell_1824_a_HPC2_and_n8, cell_1824_a_HPC2_and_n7,
         cell_1824_a_HPC2_and_p_0_out_0__1_,
         cell_1824_a_HPC2_and_p_0_out_1__0_,
         cell_1824_a_HPC2_and_p_1_out_0__1_,
         cell_1824_a_HPC2_and_p_1_out_1__0_,
         cell_1824_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1824_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1824_a_HPC2_and_p_1_in_0__1_, cell_1824_a_HPC2_and_p_1_in_1__0_,
         cell_1824_a_HPC2_and_s_out_0__1_, cell_1824_a_HPC2_and_s_out_1__0_,
         cell_1824_a_HPC2_and_p_0_in_0__1_, cell_1824_a_HPC2_and_p_0_in_1__0_,
         cell_1824_a_HPC2_and_s_in_0__1_, cell_1824_a_HPC2_and_s_in_1__0_,
         cell_1824_a_HPC2_and_z_0__0_, cell_1824_a_HPC2_and_z_1__1_,
         cell_1825_a_HPC2_and_n9, cell_1825_a_HPC2_and_n8,
         cell_1825_a_HPC2_and_n7, cell_1825_a_HPC2_and_p_0_out_0__1_,
         cell_1825_a_HPC2_and_p_0_out_1__0_,
         cell_1825_a_HPC2_and_p_1_out_0__1_,
         cell_1825_a_HPC2_and_p_1_out_1__0_,
         cell_1825_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1825_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1825_a_HPC2_and_p_1_in_0__1_, cell_1825_a_HPC2_and_p_1_in_1__0_,
         cell_1825_a_HPC2_and_s_out_0__1_, cell_1825_a_HPC2_and_s_out_1__0_,
         cell_1825_a_HPC2_and_p_0_in_0__1_, cell_1825_a_HPC2_and_p_0_in_1__0_,
         cell_1825_a_HPC2_and_s_in_0__1_, cell_1825_a_HPC2_and_s_in_1__0_,
         cell_1825_a_HPC2_and_z_0__0_, cell_1825_a_HPC2_and_z_1__1_,
         cell_1826_a_HPC2_and_n9, cell_1826_a_HPC2_and_n8,
         cell_1826_a_HPC2_and_n7, cell_1826_a_HPC2_and_p_0_out_0__1_,
         cell_1826_a_HPC2_and_p_0_out_1__0_,
         cell_1826_a_HPC2_and_p_1_out_0__1_,
         cell_1826_a_HPC2_and_p_1_out_1__0_,
         cell_1826_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1826_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1826_a_HPC2_and_p_1_in_0__1_, cell_1826_a_HPC2_and_p_1_in_1__0_,
         cell_1826_a_HPC2_and_s_out_0__1_, cell_1826_a_HPC2_and_s_out_1__0_,
         cell_1826_a_HPC2_and_p_0_in_0__1_, cell_1826_a_HPC2_and_p_0_in_1__0_,
         cell_1826_a_HPC2_and_s_in_0__1_, cell_1826_a_HPC2_and_s_in_1__0_,
         cell_1826_a_HPC2_and_z_0__0_, cell_1826_a_HPC2_and_z_1__1_,
         cell_1827_a_HPC2_and_n9, cell_1827_a_HPC2_and_n8,
         cell_1827_a_HPC2_and_n7, cell_1827_a_HPC2_and_p_0_out_0__1_,
         cell_1827_a_HPC2_and_p_0_out_1__0_,
         cell_1827_a_HPC2_and_p_1_out_0__1_,
         cell_1827_a_HPC2_and_p_1_out_1__0_,
         cell_1827_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1827_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1827_a_HPC2_and_p_1_in_0__1_, cell_1827_a_HPC2_and_p_1_in_1__0_,
         cell_1827_a_HPC2_and_s_out_0__1_, cell_1827_a_HPC2_and_s_out_1__0_,
         cell_1827_a_HPC2_and_p_0_in_0__1_, cell_1827_a_HPC2_and_p_0_in_1__0_,
         cell_1827_a_HPC2_and_s_in_0__1_, cell_1827_a_HPC2_and_s_in_1__0_,
         cell_1827_a_HPC2_and_z_0__0_, cell_1827_a_HPC2_and_z_1__1_,
         cell_1828_a_HPC2_and_n9, cell_1828_a_HPC2_and_n8,
         cell_1828_a_HPC2_and_n7, cell_1828_a_HPC2_and_p_0_out_0__1_,
         cell_1828_a_HPC2_and_p_0_out_1__0_,
         cell_1828_a_HPC2_and_p_1_out_0__1_,
         cell_1828_a_HPC2_and_p_1_out_1__0_,
         cell_1828_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1828_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1828_a_HPC2_and_p_1_in_0__1_, cell_1828_a_HPC2_and_p_1_in_1__0_,
         cell_1828_a_HPC2_and_s_out_0__1_, cell_1828_a_HPC2_and_s_out_1__0_,
         cell_1828_a_HPC2_and_p_0_in_0__1_, cell_1828_a_HPC2_and_p_0_in_1__0_,
         cell_1828_a_HPC2_and_s_in_0__1_, cell_1828_a_HPC2_and_s_in_1__0_,
         cell_1828_a_HPC2_and_z_0__0_, cell_1828_a_HPC2_and_z_1__1_,
         cell_1829_a_HPC2_and_n9, cell_1829_a_HPC2_and_n8,
         cell_1829_a_HPC2_and_n7, cell_1829_a_HPC2_and_p_0_out_0__1_,
         cell_1829_a_HPC2_and_p_0_out_1__0_,
         cell_1829_a_HPC2_and_p_1_out_0__1_,
         cell_1829_a_HPC2_and_p_1_out_1__0_,
         cell_1829_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1829_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1829_a_HPC2_and_p_1_in_0__1_, cell_1829_a_HPC2_and_p_1_in_1__0_,
         cell_1829_a_HPC2_and_s_out_0__1_, cell_1829_a_HPC2_and_s_out_1__0_,
         cell_1829_a_HPC2_and_p_0_in_0__1_, cell_1829_a_HPC2_and_p_0_in_1__0_,
         cell_1829_a_HPC2_and_s_in_0__1_, cell_1829_a_HPC2_and_s_in_1__0_,
         cell_1829_a_HPC2_and_z_0__0_, cell_1829_a_HPC2_and_z_1__1_,
         cell_1830_a_HPC2_and_n9, cell_1830_a_HPC2_and_n8,
         cell_1830_a_HPC2_and_n7, cell_1830_a_HPC2_and_p_0_out_0__1_,
         cell_1830_a_HPC2_and_p_0_out_1__0_,
         cell_1830_a_HPC2_and_p_1_out_0__1_,
         cell_1830_a_HPC2_and_p_1_out_1__0_,
         cell_1830_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1830_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1830_a_HPC2_and_p_1_in_0__1_, cell_1830_a_HPC2_and_p_1_in_1__0_,
         cell_1830_a_HPC2_and_s_out_0__1_, cell_1830_a_HPC2_and_s_out_1__0_,
         cell_1830_a_HPC2_and_p_0_in_0__1_, cell_1830_a_HPC2_and_p_0_in_1__0_,
         cell_1830_a_HPC2_and_s_in_0__1_, cell_1830_a_HPC2_and_s_in_1__0_,
         cell_1830_a_HPC2_and_z_0__0_, cell_1830_a_HPC2_and_z_1__1_,
         cell_1831_a_HPC2_and_n9, cell_1831_a_HPC2_and_n8,
         cell_1831_a_HPC2_and_n7, cell_1831_a_HPC2_and_p_0_out_0__1_,
         cell_1831_a_HPC2_and_p_0_out_1__0_,
         cell_1831_a_HPC2_and_p_1_out_0__1_,
         cell_1831_a_HPC2_and_p_1_out_1__0_,
         cell_1831_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1831_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1831_a_HPC2_and_p_1_in_0__1_, cell_1831_a_HPC2_and_p_1_in_1__0_,
         cell_1831_a_HPC2_and_s_out_0__1_, cell_1831_a_HPC2_and_s_out_1__0_,
         cell_1831_a_HPC2_and_p_0_in_0__1_, cell_1831_a_HPC2_and_p_0_in_1__0_,
         cell_1831_a_HPC2_and_s_in_0__1_, cell_1831_a_HPC2_and_s_in_1__0_,
         cell_1831_a_HPC2_and_z_0__0_, cell_1831_a_HPC2_and_z_1__1_,
         cell_1832_a_HPC2_and_n9, cell_1832_a_HPC2_and_n8,
         cell_1832_a_HPC2_and_n7, cell_1832_a_HPC2_and_p_0_out_0__1_,
         cell_1832_a_HPC2_and_p_0_out_1__0_,
         cell_1832_a_HPC2_and_p_1_out_0__1_,
         cell_1832_a_HPC2_and_p_1_out_1__0_,
         cell_1832_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1832_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1832_a_HPC2_and_p_1_in_0__1_, cell_1832_a_HPC2_and_p_1_in_1__0_,
         cell_1832_a_HPC2_and_s_out_0__1_, cell_1832_a_HPC2_and_s_out_1__0_,
         cell_1832_a_HPC2_and_p_0_in_0__1_, cell_1832_a_HPC2_and_p_0_in_1__0_,
         cell_1832_a_HPC2_and_s_in_0__1_, cell_1832_a_HPC2_and_s_in_1__0_,
         cell_1832_a_HPC2_and_z_0__0_, cell_1832_a_HPC2_and_z_1__1_,
         cell_1833_a_HPC2_and_n9, cell_1833_a_HPC2_and_n8,
         cell_1833_a_HPC2_and_n7, cell_1833_a_HPC2_and_p_0_out_0__1_,
         cell_1833_a_HPC2_and_p_0_out_1__0_,
         cell_1833_a_HPC2_and_p_1_out_0__1_,
         cell_1833_a_HPC2_and_p_1_out_1__0_,
         cell_1833_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1833_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1833_a_HPC2_and_p_1_in_0__1_, cell_1833_a_HPC2_and_p_1_in_1__0_,
         cell_1833_a_HPC2_and_s_out_0__1_, cell_1833_a_HPC2_and_s_out_1__0_,
         cell_1833_a_HPC2_and_p_0_in_0__1_, cell_1833_a_HPC2_and_p_0_in_1__0_,
         cell_1833_a_HPC2_and_s_in_0__1_, cell_1833_a_HPC2_and_s_in_1__0_,
         cell_1833_a_HPC2_and_z_0__0_, cell_1833_a_HPC2_and_z_1__1_,
         cell_1834_a_HPC2_and_n9, cell_1834_a_HPC2_and_n8,
         cell_1834_a_HPC2_and_n7, cell_1834_a_HPC2_and_p_0_out_0__1_,
         cell_1834_a_HPC2_and_p_0_out_1__0_,
         cell_1834_a_HPC2_and_p_1_out_0__1_,
         cell_1834_a_HPC2_and_p_1_out_1__0_,
         cell_1834_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1834_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1834_a_HPC2_and_p_1_in_0__1_, cell_1834_a_HPC2_and_p_1_in_1__0_,
         cell_1834_a_HPC2_and_s_out_0__1_, cell_1834_a_HPC2_and_s_out_1__0_,
         cell_1834_a_HPC2_and_p_0_in_0__1_, cell_1834_a_HPC2_and_p_0_in_1__0_,
         cell_1834_a_HPC2_and_s_in_0__1_, cell_1834_a_HPC2_and_s_in_1__0_,
         cell_1834_a_HPC2_and_z_0__0_, cell_1834_a_HPC2_and_z_1__1_,
         cell_1835_a_HPC2_and_n9, cell_1835_a_HPC2_and_n8,
         cell_1835_a_HPC2_and_n7, cell_1835_a_HPC2_and_p_0_out_0__1_,
         cell_1835_a_HPC2_and_p_0_out_1__0_,
         cell_1835_a_HPC2_and_p_1_out_0__1_,
         cell_1835_a_HPC2_and_p_1_out_1__0_,
         cell_1835_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1835_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1835_a_HPC2_and_p_1_in_0__1_, cell_1835_a_HPC2_and_p_1_in_1__0_,
         cell_1835_a_HPC2_and_s_out_0__1_, cell_1835_a_HPC2_and_s_out_1__0_,
         cell_1835_a_HPC2_and_p_0_in_0__1_, cell_1835_a_HPC2_and_p_0_in_1__0_,
         cell_1835_a_HPC2_and_s_in_0__1_, cell_1835_a_HPC2_and_s_in_1__0_,
         cell_1835_a_HPC2_and_z_0__0_, cell_1835_a_HPC2_and_z_1__1_,
         cell_1836_a_HPC2_and_n9, cell_1836_a_HPC2_and_n8,
         cell_1836_a_HPC2_and_n7, cell_1836_a_HPC2_and_p_0_out_0__1_,
         cell_1836_a_HPC2_and_p_0_out_1__0_,
         cell_1836_a_HPC2_and_p_1_out_0__1_,
         cell_1836_a_HPC2_and_p_1_out_1__0_,
         cell_1836_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1836_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1836_a_HPC2_and_p_1_in_0__1_, cell_1836_a_HPC2_and_p_1_in_1__0_,
         cell_1836_a_HPC2_and_s_out_0__1_, cell_1836_a_HPC2_and_s_out_1__0_,
         cell_1836_a_HPC2_and_p_0_in_0__1_, cell_1836_a_HPC2_and_p_0_in_1__0_,
         cell_1836_a_HPC2_and_s_in_0__1_, cell_1836_a_HPC2_and_s_in_1__0_,
         cell_1836_a_HPC2_and_z_0__0_, cell_1836_a_HPC2_and_z_1__1_,
         cell_1837_a_HPC2_and_n9, cell_1837_a_HPC2_and_n8,
         cell_1837_a_HPC2_and_n7, cell_1837_a_HPC2_and_p_0_out_0__1_,
         cell_1837_a_HPC2_and_p_0_out_1__0_,
         cell_1837_a_HPC2_and_p_1_out_0__1_,
         cell_1837_a_HPC2_and_p_1_out_1__0_,
         cell_1837_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1837_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1837_a_HPC2_and_p_1_in_0__1_, cell_1837_a_HPC2_and_p_1_in_1__0_,
         cell_1837_a_HPC2_and_s_out_0__1_, cell_1837_a_HPC2_and_s_out_1__0_,
         cell_1837_a_HPC2_and_p_0_in_0__1_, cell_1837_a_HPC2_and_p_0_in_1__0_,
         cell_1837_a_HPC2_and_s_in_0__1_, cell_1837_a_HPC2_and_s_in_1__0_,
         cell_1837_a_HPC2_and_z_0__0_, cell_1837_a_HPC2_and_z_1__1_,
         cell_1838_a_HPC2_and_n9, cell_1838_a_HPC2_and_n8,
         cell_1838_a_HPC2_and_n7, cell_1838_a_HPC2_and_p_0_out_0__1_,
         cell_1838_a_HPC2_and_p_0_out_1__0_,
         cell_1838_a_HPC2_and_p_1_out_0__1_,
         cell_1838_a_HPC2_and_p_1_out_1__0_,
         cell_1838_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1838_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1838_a_HPC2_and_p_1_in_0__1_, cell_1838_a_HPC2_and_p_1_in_1__0_,
         cell_1838_a_HPC2_and_s_out_0__1_, cell_1838_a_HPC2_and_s_out_1__0_,
         cell_1838_a_HPC2_and_p_0_in_0__1_, cell_1838_a_HPC2_and_p_0_in_1__0_,
         cell_1838_a_HPC2_and_s_in_0__1_, cell_1838_a_HPC2_and_s_in_1__0_,
         cell_1838_a_HPC2_and_z_0__0_, cell_1838_a_HPC2_and_z_1__1_,
         cell_1839_a_HPC2_and_n9, cell_1839_a_HPC2_and_n8,
         cell_1839_a_HPC2_and_n7, cell_1839_a_HPC2_and_p_0_out_0__1_,
         cell_1839_a_HPC2_and_p_0_out_1__0_,
         cell_1839_a_HPC2_and_p_1_out_0__1_,
         cell_1839_a_HPC2_and_p_1_out_1__0_,
         cell_1839_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1839_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1839_a_HPC2_and_p_1_in_0__1_, cell_1839_a_HPC2_and_p_1_in_1__0_,
         cell_1839_a_HPC2_and_s_out_0__1_, cell_1839_a_HPC2_and_s_out_1__0_,
         cell_1839_a_HPC2_and_p_0_in_0__1_, cell_1839_a_HPC2_and_p_0_in_1__0_,
         cell_1839_a_HPC2_and_s_in_0__1_, cell_1839_a_HPC2_and_s_in_1__0_,
         cell_1839_a_HPC2_and_z_0__0_, cell_1839_a_HPC2_and_z_1__1_,
         cell_1840_a_HPC2_and_n9, cell_1840_a_HPC2_and_n8,
         cell_1840_a_HPC2_and_n7, cell_1840_a_HPC2_and_p_0_out_0__1_,
         cell_1840_a_HPC2_and_p_0_out_1__0_,
         cell_1840_a_HPC2_and_p_1_out_0__1_,
         cell_1840_a_HPC2_and_p_1_out_1__0_,
         cell_1840_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1840_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1840_a_HPC2_and_p_1_in_0__1_, cell_1840_a_HPC2_and_p_1_in_1__0_,
         cell_1840_a_HPC2_and_s_out_0__1_, cell_1840_a_HPC2_and_s_out_1__0_,
         cell_1840_a_HPC2_and_p_0_in_0__1_, cell_1840_a_HPC2_and_p_0_in_1__0_,
         cell_1840_a_HPC2_and_s_in_0__1_, cell_1840_a_HPC2_and_s_in_1__0_,
         cell_1840_a_HPC2_and_z_0__0_, cell_1840_a_HPC2_and_z_1__1_,
         cell_1841_a_HPC2_and_n9, cell_1841_a_HPC2_and_n8,
         cell_1841_a_HPC2_and_n7, cell_1841_a_HPC2_and_p_0_out_0__1_,
         cell_1841_a_HPC2_and_p_0_out_1__0_,
         cell_1841_a_HPC2_and_p_1_out_0__1_,
         cell_1841_a_HPC2_and_p_1_out_1__0_,
         cell_1841_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1841_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1841_a_HPC2_and_p_1_in_0__1_, cell_1841_a_HPC2_and_p_1_in_1__0_,
         cell_1841_a_HPC2_and_s_out_0__1_, cell_1841_a_HPC2_and_s_out_1__0_,
         cell_1841_a_HPC2_and_p_0_in_0__1_, cell_1841_a_HPC2_and_p_0_in_1__0_,
         cell_1841_a_HPC2_and_s_in_0__1_, cell_1841_a_HPC2_and_s_in_1__0_,
         cell_1841_a_HPC2_and_z_0__0_, cell_1841_a_HPC2_and_z_1__1_,
         cell_1842_a_HPC2_and_n9, cell_1842_a_HPC2_and_n8,
         cell_1842_a_HPC2_and_n7, cell_1842_a_HPC2_and_p_0_out_0__1_,
         cell_1842_a_HPC2_and_p_0_out_1__0_,
         cell_1842_a_HPC2_and_p_1_out_0__1_,
         cell_1842_a_HPC2_and_p_1_out_1__0_,
         cell_1842_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1842_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1842_a_HPC2_and_p_1_in_0__1_, cell_1842_a_HPC2_and_p_1_in_1__0_,
         cell_1842_a_HPC2_and_s_out_0__1_, cell_1842_a_HPC2_and_s_out_1__0_,
         cell_1842_a_HPC2_and_p_0_in_0__1_, cell_1842_a_HPC2_and_p_0_in_1__0_,
         cell_1842_a_HPC2_and_s_in_0__1_, cell_1842_a_HPC2_and_s_in_1__0_,
         cell_1842_a_HPC2_and_z_0__0_, cell_1842_a_HPC2_and_z_1__1_,
         cell_1843_a_HPC2_and_n9, cell_1843_a_HPC2_and_n8,
         cell_1843_a_HPC2_and_n7, cell_1843_a_HPC2_and_p_0_out_0__1_,
         cell_1843_a_HPC2_and_p_0_out_1__0_,
         cell_1843_a_HPC2_and_p_1_out_0__1_,
         cell_1843_a_HPC2_and_p_1_out_1__0_,
         cell_1843_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1843_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1843_a_HPC2_and_p_1_in_0__1_, cell_1843_a_HPC2_and_p_1_in_1__0_,
         cell_1843_a_HPC2_and_s_out_0__1_, cell_1843_a_HPC2_and_s_out_1__0_,
         cell_1843_a_HPC2_and_p_0_in_0__1_, cell_1843_a_HPC2_and_p_0_in_1__0_,
         cell_1843_a_HPC2_and_s_in_0__1_, cell_1843_a_HPC2_and_s_in_1__0_,
         cell_1843_a_HPC2_and_z_0__0_, cell_1843_a_HPC2_and_z_1__1_,
         cell_1844_a_HPC2_and_n9, cell_1844_a_HPC2_and_n8,
         cell_1844_a_HPC2_and_n7, cell_1844_a_HPC2_and_p_0_out_0__1_,
         cell_1844_a_HPC2_and_p_0_out_1__0_,
         cell_1844_a_HPC2_and_p_1_out_0__1_,
         cell_1844_a_HPC2_and_p_1_out_1__0_,
         cell_1844_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1844_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1844_a_HPC2_and_p_1_in_0__1_, cell_1844_a_HPC2_and_p_1_in_1__0_,
         cell_1844_a_HPC2_and_s_out_0__1_, cell_1844_a_HPC2_and_s_out_1__0_,
         cell_1844_a_HPC2_and_p_0_in_0__1_, cell_1844_a_HPC2_and_p_0_in_1__0_,
         cell_1844_a_HPC2_and_s_in_0__1_, cell_1844_a_HPC2_and_s_in_1__0_,
         cell_1844_a_HPC2_and_z_0__0_, cell_1844_a_HPC2_and_z_1__1_,
         cell_1845_a_HPC2_and_n9, cell_1845_a_HPC2_and_n8,
         cell_1845_a_HPC2_and_n7, cell_1845_a_HPC2_and_p_0_out_0__1_,
         cell_1845_a_HPC2_and_p_0_out_1__0_,
         cell_1845_a_HPC2_and_p_1_out_0__1_,
         cell_1845_a_HPC2_and_p_1_out_1__0_,
         cell_1845_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1845_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1845_a_HPC2_and_p_1_in_0__1_, cell_1845_a_HPC2_and_p_1_in_1__0_,
         cell_1845_a_HPC2_and_s_out_0__1_, cell_1845_a_HPC2_and_s_out_1__0_,
         cell_1845_a_HPC2_and_p_0_in_0__1_, cell_1845_a_HPC2_and_p_0_in_1__0_,
         cell_1845_a_HPC2_and_s_in_0__1_, cell_1845_a_HPC2_and_s_in_1__0_,
         cell_1845_a_HPC2_and_z_0__0_, cell_1845_a_HPC2_and_z_1__1_,
         cell_1846_a_HPC2_and_n9, cell_1846_a_HPC2_and_n8,
         cell_1846_a_HPC2_and_n7, cell_1846_a_HPC2_and_p_0_out_0__1_,
         cell_1846_a_HPC2_and_p_0_out_1__0_,
         cell_1846_a_HPC2_and_p_1_out_0__1_,
         cell_1846_a_HPC2_and_p_1_out_1__0_,
         cell_1846_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1846_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1846_a_HPC2_and_p_1_in_0__1_, cell_1846_a_HPC2_and_p_1_in_1__0_,
         cell_1846_a_HPC2_and_s_out_0__1_, cell_1846_a_HPC2_and_s_out_1__0_,
         cell_1846_a_HPC2_and_p_0_in_0__1_, cell_1846_a_HPC2_and_p_0_in_1__0_,
         cell_1846_a_HPC2_and_s_in_0__1_, cell_1846_a_HPC2_and_s_in_1__0_,
         cell_1846_a_HPC2_and_z_0__0_, cell_1846_a_HPC2_and_z_1__1_,
         cell_1847_a_HPC2_and_n9, cell_1847_a_HPC2_and_n8,
         cell_1847_a_HPC2_and_n7, cell_1847_a_HPC2_and_p_0_out_0__1_,
         cell_1847_a_HPC2_and_p_0_out_1__0_,
         cell_1847_a_HPC2_and_p_1_out_0__1_,
         cell_1847_a_HPC2_and_p_1_out_1__0_,
         cell_1847_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1847_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1847_a_HPC2_and_p_1_in_0__1_, cell_1847_a_HPC2_and_p_1_in_1__0_,
         cell_1847_a_HPC2_and_s_out_0__1_, cell_1847_a_HPC2_and_s_out_1__0_,
         cell_1847_a_HPC2_and_p_0_in_0__1_, cell_1847_a_HPC2_and_p_0_in_1__0_,
         cell_1847_a_HPC2_and_s_in_0__1_, cell_1847_a_HPC2_and_s_in_1__0_,
         cell_1847_a_HPC2_and_z_0__0_, cell_1847_a_HPC2_and_z_1__1_,
         cell_1848_a_HPC2_and_n9, cell_1848_a_HPC2_and_n8,
         cell_1848_a_HPC2_and_n7, cell_1848_a_HPC2_and_p_0_out_0__1_,
         cell_1848_a_HPC2_and_p_0_out_1__0_,
         cell_1848_a_HPC2_and_p_1_out_0__1_,
         cell_1848_a_HPC2_and_p_1_out_1__0_,
         cell_1848_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1848_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1848_a_HPC2_and_p_1_in_0__1_, cell_1848_a_HPC2_and_p_1_in_1__0_,
         cell_1848_a_HPC2_and_s_out_0__1_, cell_1848_a_HPC2_and_s_out_1__0_,
         cell_1848_a_HPC2_and_p_0_in_0__1_, cell_1848_a_HPC2_and_p_0_in_1__0_,
         cell_1848_a_HPC2_and_s_in_0__1_, cell_1848_a_HPC2_and_s_in_1__0_,
         cell_1848_a_HPC2_and_z_0__0_, cell_1848_a_HPC2_and_z_1__1_,
         cell_1849_a_HPC2_and_n9, cell_1849_a_HPC2_and_n8,
         cell_1849_a_HPC2_and_n7, cell_1849_a_HPC2_and_p_0_out_0__1_,
         cell_1849_a_HPC2_and_p_0_out_1__0_,
         cell_1849_a_HPC2_and_p_1_out_0__1_,
         cell_1849_a_HPC2_and_p_1_out_1__0_,
         cell_1849_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1849_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1849_a_HPC2_and_p_1_in_0__1_, cell_1849_a_HPC2_and_p_1_in_1__0_,
         cell_1849_a_HPC2_and_s_out_0__1_, cell_1849_a_HPC2_and_s_out_1__0_,
         cell_1849_a_HPC2_and_p_0_in_0__1_, cell_1849_a_HPC2_and_p_0_in_1__0_,
         cell_1849_a_HPC2_and_s_in_0__1_, cell_1849_a_HPC2_and_s_in_1__0_,
         cell_1849_a_HPC2_and_z_0__0_, cell_1849_a_HPC2_and_z_1__1_,
         cell_1850_a_HPC2_and_n9, cell_1850_a_HPC2_and_n8,
         cell_1850_a_HPC2_and_n7, cell_1850_a_HPC2_and_p_0_out_0__1_,
         cell_1850_a_HPC2_and_p_0_out_1__0_,
         cell_1850_a_HPC2_and_p_1_out_0__1_,
         cell_1850_a_HPC2_and_p_1_out_1__0_,
         cell_1850_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1850_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1850_a_HPC2_and_p_1_in_0__1_, cell_1850_a_HPC2_and_p_1_in_1__0_,
         cell_1850_a_HPC2_and_s_out_0__1_, cell_1850_a_HPC2_and_s_out_1__0_,
         cell_1850_a_HPC2_and_p_0_in_0__1_, cell_1850_a_HPC2_and_p_0_in_1__0_,
         cell_1850_a_HPC2_and_s_in_0__1_, cell_1850_a_HPC2_and_s_in_1__0_,
         cell_1850_a_HPC2_and_z_0__0_, cell_1850_a_HPC2_and_z_1__1_,
         cell_1851_a_HPC2_and_n9, cell_1851_a_HPC2_and_n8,
         cell_1851_a_HPC2_and_n7, cell_1851_a_HPC2_and_p_0_out_0__1_,
         cell_1851_a_HPC2_and_p_0_out_1__0_,
         cell_1851_a_HPC2_and_p_1_out_0__1_,
         cell_1851_a_HPC2_and_p_1_out_1__0_,
         cell_1851_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1851_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1851_a_HPC2_and_p_1_in_0__1_, cell_1851_a_HPC2_and_p_1_in_1__0_,
         cell_1851_a_HPC2_and_s_out_0__1_, cell_1851_a_HPC2_and_s_out_1__0_,
         cell_1851_a_HPC2_and_p_0_in_0__1_, cell_1851_a_HPC2_and_p_0_in_1__0_,
         cell_1851_a_HPC2_and_s_in_0__1_, cell_1851_a_HPC2_and_s_in_1__0_,
         cell_1851_a_HPC2_and_z_0__0_, cell_1851_a_HPC2_and_z_1__1_,
         cell_1852_a_HPC2_and_n9, cell_1852_a_HPC2_and_n8,
         cell_1852_a_HPC2_and_n7, cell_1852_a_HPC2_and_p_0_out_0__1_,
         cell_1852_a_HPC2_and_p_0_out_1__0_,
         cell_1852_a_HPC2_and_p_1_out_0__1_,
         cell_1852_a_HPC2_and_p_1_out_1__0_,
         cell_1852_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1852_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1852_a_HPC2_and_p_1_in_0__1_, cell_1852_a_HPC2_and_p_1_in_1__0_,
         cell_1852_a_HPC2_and_s_out_0__1_, cell_1852_a_HPC2_and_s_out_1__0_,
         cell_1852_a_HPC2_and_p_0_in_0__1_, cell_1852_a_HPC2_and_p_0_in_1__0_,
         cell_1852_a_HPC2_and_s_in_0__1_, cell_1852_a_HPC2_and_s_in_1__0_,
         cell_1852_a_HPC2_and_z_0__0_, cell_1852_a_HPC2_and_z_1__1_,
         cell_1853_a_HPC2_and_n9, cell_1853_a_HPC2_and_n8,
         cell_1853_a_HPC2_and_n7, cell_1853_a_HPC2_and_p_0_out_0__1_,
         cell_1853_a_HPC2_and_p_0_out_1__0_,
         cell_1853_a_HPC2_and_p_1_out_0__1_,
         cell_1853_a_HPC2_and_p_1_out_1__0_,
         cell_1853_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1853_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1853_a_HPC2_and_p_1_in_0__1_, cell_1853_a_HPC2_and_p_1_in_1__0_,
         cell_1853_a_HPC2_and_s_out_0__1_, cell_1853_a_HPC2_and_s_out_1__0_,
         cell_1853_a_HPC2_and_p_0_in_0__1_, cell_1853_a_HPC2_and_p_0_in_1__0_,
         cell_1853_a_HPC2_and_s_in_0__1_, cell_1853_a_HPC2_and_s_in_1__0_,
         cell_1853_a_HPC2_and_z_0__0_, cell_1853_a_HPC2_and_z_1__1_,
         cell_1854_a_HPC2_and_n9, cell_1854_a_HPC2_and_n8,
         cell_1854_a_HPC2_and_n7, cell_1854_a_HPC2_and_p_0_out_0__1_,
         cell_1854_a_HPC2_and_p_0_out_1__0_,
         cell_1854_a_HPC2_and_p_1_out_0__1_,
         cell_1854_a_HPC2_and_p_1_out_1__0_,
         cell_1854_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1854_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1854_a_HPC2_and_p_1_in_0__1_, cell_1854_a_HPC2_and_p_1_in_1__0_,
         cell_1854_a_HPC2_and_s_out_0__1_, cell_1854_a_HPC2_and_s_out_1__0_,
         cell_1854_a_HPC2_and_p_0_in_0__1_, cell_1854_a_HPC2_and_p_0_in_1__0_,
         cell_1854_a_HPC2_and_s_in_0__1_, cell_1854_a_HPC2_and_s_in_1__0_,
         cell_1854_a_HPC2_and_z_0__0_, cell_1854_a_HPC2_and_z_1__1_,
         cell_1855_a_HPC2_and_n9, cell_1855_a_HPC2_and_n8,
         cell_1855_a_HPC2_and_n7, cell_1855_a_HPC2_and_p_0_out_0__1_,
         cell_1855_a_HPC2_and_p_0_out_1__0_,
         cell_1855_a_HPC2_and_p_1_out_0__1_,
         cell_1855_a_HPC2_and_p_1_out_1__0_,
         cell_1855_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1855_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1855_a_HPC2_and_p_1_in_0__1_, cell_1855_a_HPC2_and_p_1_in_1__0_,
         cell_1855_a_HPC2_and_s_out_0__1_, cell_1855_a_HPC2_and_s_out_1__0_,
         cell_1855_a_HPC2_and_p_0_in_0__1_, cell_1855_a_HPC2_and_p_0_in_1__0_,
         cell_1855_a_HPC2_and_s_in_0__1_, cell_1855_a_HPC2_and_s_in_1__0_,
         cell_1855_a_HPC2_and_z_0__0_, cell_1855_a_HPC2_and_z_1__1_,
         cell_1856_a_HPC2_and_n9, cell_1856_a_HPC2_and_n8,
         cell_1856_a_HPC2_and_n7, cell_1856_a_HPC2_and_p_0_out_0__1_,
         cell_1856_a_HPC2_and_p_0_out_1__0_,
         cell_1856_a_HPC2_and_p_1_out_0__1_,
         cell_1856_a_HPC2_and_p_1_out_1__0_,
         cell_1856_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1856_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1856_a_HPC2_and_p_1_in_0__1_, cell_1856_a_HPC2_and_p_1_in_1__0_,
         cell_1856_a_HPC2_and_s_out_0__1_, cell_1856_a_HPC2_and_s_out_1__0_,
         cell_1856_a_HPC2_and_p_0_in_0__1_, cell_1856_a_HPC2_and_p_0_in_1__0_,
         cell_1856_a_HPC2_and_s_in_0__1_, cell_1856_a_HPC2_and_s_in_1__0_,
         cell_1856_a_HPC2_and_z_0__0_, cell_1856_a_HPC2_and_z_1__1_,
         cell_1857_a_HPC2_and_n9, cell_1857_a_HPC2_and_n8,
         cell_1857_a_HPC2_and_n7, cell_1857_a_HPC2_and_p_0_out_0__1_,
         cell_1857_a_HPC2_and_p_0_out_1__0_,
         cell_1857_a_HPC2_and_p_1_out_0__1_,
         cell_1857_a_HPC2_and_p_1_out_1__0_,
         cell_1857_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1857_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1857_a_HPC2_and_p_1_in_0__1_, cell_1857_a_HPC2_and_p_1_in_1__0_,
         cell_1857_a_HPC2_and_s_out_0__1_, cell_1857_a_HPC2_and_s_out_1__0_,
         cell_1857_a_HPC2_and_p_0_in_0__1_, cell_1857_a_HPC2_and_p_0_in_1__0_,
         cell_1857_a_HPC2_and_s_in_0__1_, cell_1857_a_HPC2_and_s_in_1__0_,
         cell_1857_a_HPC2_and_z_0__0_, cell_1857_a_HPC2_and_z_1__1_,
         cell_1858_a_HPC2_and_n9, cell_1858_a_HPC2_and_n8,
         cell_1858_a_HPC2_and_n7, cell_1858_a_HPC2_and_p_0_out_0__1_,
         cell_1858_a_HPC2_and_p_0_out_1__0_,
         cell_1858_a_HPC2_and_p_1_out_0__1_,
         cell_1858_a_HPC2_and_p_1_out_1__0_,
         cell_1858_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1858_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1858_a_HPC2_and_p_1_in_0__1_, cell_1858_a_HPC2_and_p_1_in_1__0_,
         cell_1858_a_HPC2_and_s_out_0__1_, cell_1858_a_HPC2_and_s_out_1__0_,
         cell_1858_a_HPC2_and_p_0_in_0__1_, cell_1858_a_HPC2_and_p_0_in_1__0_,
         cell_1858_a_HPC2_and_s_in_0__1_, cell_1858_a_HPC2_and_s_in_1__0_,
         cell_1858_a_HPC2_and_z_0__0_, cell_1858_a_HPC2_and_z_1__1_,
         cell_1859_a_HPC2_and_n9, cell_1859_a_HPC2_and_n8,
         cell_1859_a_HPC2_and_n7, cell_1859_a_HPC2_and_p_0_out_0__1_,
         cell_1859_a_HPC2_and_p_0_out_1__0_,
         cell_1859_a_HPC2_and_p_1_out_0__1_,
         cell_1859_a_HPC2_and_p_1_out_1__0_,
         cell_1859_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1859_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1859_a_HPC2_and_p_1_in_0__1_, cell_1859_a_HPC2_and_p_1_in_1__0_,
         cell_1859_a_HPC2_and_s_out_0__1_, cell_1859_a_HPC2_and_s_out_1__0_,
         cell_1859_a_HPC2_and_p_0_in_0__1_, cell_1859_a_HPC2_and_p_0_in_1__0_,
         cell_1859_a_HPC2_and_s_in_0__1_, cell_1859_a_HPC2_and_s_in_1__0_,
         cell_1859_a_HPC2_and_z_0__0_, cell_1859_a_HPC2_and_z_1__1_,
         cell_1860_a_HPC2_and_n9, cell_1860_a_HPC2_and_n8,
         cell_1860_a_HPC2_and_n7, cell_1860_a_HPC2_and_p_0_out_0__1_,
         cell_1860_a_HPC2_and_p_0_out_1__0_,
         cell_1860_a_HPC2_and_p_1_out_0__1_,
         cell_1860_a_HPC2_and_p_1_out_1__0_,
         cell_1860_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1860_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1860_a_HPC2_and_p_1_in_0__1_, cell_1860_a_HPC2_and_p_1_in_1__0_,
         cell_1860_a_HPC2_and_s_out_0__1_, cell_1860_a_HPC2_and_s_out_1__0_,
         cell_1860_a_HPC2_and_p_0_in_0__1_, cell_1860_a_HPC2_and_p_0_in_1__0_,
         cell_1860_a_HPC2_and_s_in_0__1_, cell_1860_a_HPC2_and_s_in_1__0_,
         cell_1860_a_HPC2_and_z_0__0_, cell_1860_a_HPC2_and_z_1__1_,
         cell_1861_a_HPC2_and_n9, cell_1861_a_HPC2_and_n8,
         cell_1861_a_HPC2_and_n7, cell_1861_a_HPC2_and_p_0_out_0__1_,
         cell_1861_a_HPC2_and_p_0_out_1__0_,
         cell_1861_a_HPC2_and_p_1_out_0__1_,
         cell_1861_a_HPC2_and_p_1_out_1__0_,
         cell_1861_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1861_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1861_a_HPC2_and_p_1_in_0__1_, cell_1861_a_HPC2_and_p_1_in_1__0_,
         cell_1861_a_HPC2_and_s_out_0__1_, cell_1861_a_HPC2_and_s_out_1__0_,
         cell_1861_a_HPC2_and_p_0_in_0__1_, cell_1861_a_HPC2_and_p_0_in_1__0_,
         cell_1861_a_HPC2_and_s_in_0__1_, cell_1861_a_HPC2_and_s_in_1__0_,
         cell_1861_a_HPC2_and_z_0__0_, cell_1861_a_HPC2_and_z_1__1_,
         cell_1862_a_HPC2_and_n9, cell_1862_a_HPC2_and_n8,
         cell_1862_a_HPC2_and_n7, cell_1862_a_HPC2_and_p_0_out_0__1_,
         cell_1862_a_HPC2_and_p_0_out_1__0_,
         cell_1862_a_HPC2_and_p_1_out_0__1_,
         cell_1862_a_HPC2_and_p_1_out_1__0_,
         cell_1862_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1862_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1862_a_HPC2_and_p_1_in_0__1_, cell_1862_a_HPC2_and_p_1_in_1__0_,
         cell_1862_a_HPC2_and_s_out_0__1_, cell_1862_a_HPC2_and_s_out_1__0_,
         cell_1862_a_HPC2_and_p_0_in_0__1_, cell_1862_a_HPC2_and_p_0_in_1__0_,
         cell_1862_a_HPC2_and_s_in_0__1_, cell_1862_a_HPC2_and_s_in_1__0_,
         cell_1862_a_HPC2_and_z_0__0_, cell_1862_a_HPC2_and_z_1__1_,
         cell_1863_a_HPC2_and_n9, cell_1863_a_HPC2_and_n8,
         cell_1863_a_HPC2_and_n7, cell_1863_a_HPC2_and_p_0_out_0__1_,
         cell_1863_a_HPC2_and_p_0_out_1__0_,
         cell_1863_a_HPC2_and_p_1_out_0__1_,
         cell_1863_a_HPC2_and_p_1_out_1__0_,
         cell_1863_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1863_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1863_a_HPC2_and_p_1_in_0__1_, cell_1863_a_HPC2_and_p_1_in_1__0_,
         cell_1863_a_HPC2_and_s_out_0__1_, cell_1863_a_HPC2_and_s_out_1__0_,
         cell_1863_a_HPC2_and_p_0_in_0__1_, cell_1863_a_HPC2_and_p_0_in_1__0_,
         cell_1863_a_HPC2_and_s_in_0__1_, cell_1863_a_HPC2_and_s_in_1__0_,
         cell_1863_a_HPC2_and_z_0__0_, cell_1863_a_HPC2_and_z_1__1_,
         cell_1864_a_HPC2_and_n9, cell_1864_a_HPC2_and_n8,
         cell_1864_a_HPC2_and_n7, cell_1864_a_HPC2_and_p_0_out_0__1_,
         cell_1864_a_HPC2_and_p_0_out_1__0_,
         cell_1864_a_HPC2_and_p_1_out_0__1_,
         cell_1864_a_HPC2_and_p_1_out_1__0_,
         cell_1864_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1864_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1864_a_HPC2_and_p_1_in_0__1_, cell_1864_a_HPC2_and_p_1_in_1__0_,
         cell_1864_a_HPC2_and_s_out_0__1_, cell_1864_a_HPC2_and_s_out_1__0_,
         cell_1864_a_HPC2_and_p_0_in_0__1_, cell_1864_a_HPC2_and_p_0_in_1__0_,
         cell_1864_a_HPC2_and_s_in_0__1_, cell_1864_a_HPC2_and_s_in_1__0_,
         cell_1864_a_HPC2_and_z_0__0_, cell_1864_a_HPC2_and_z_1__1_,
         cell_1865_a_HPC2_and_n9, cell_1865_a_HPC2_and_n8,
         cell_1865_a_HPC2_and_n7, cell_1865_a_HPC2_and_p_0_out_0__1_,
         cell_1865_a_HPC2_and_p_0_out_1__0_,
         cell_1865_a_HPC2_and_p_1_out_0__1_,
         cell_1865_a_HPC2_and_p_1_out_1__0_,
         cell_1865_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1865_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1865_a_HPC2_and_p_1_in_0__1_, cell_1865_a_HPC2_and_p_1_in_1__0_,
         cell_1865_a_HPC2_and_s_out_0__1_, cell_1865_a_HPC2_and_s_out_1__0_,
         cell_1865_a_HPC2_and_p_0_in_0__1_, cell_1865_a_HPC2_and_p_0_in_1__0_,
         cell_1865_a_HPC2_and_s_in_0__1_, cell_1865_a_HPC2_and_s_in_1__0_,
         cell_1865_a_HPC2_and_z_0__0_, cell_1865_a_HPC2_and_z_1__1_,
         cell_1866_a_HPC2_and_n9, cell_1866_a_HPC2_and_n8,
         cell_1866_a_HPC2_and_n7, cell_1866_a_HPC2_and_p_0_out_0__1_,
         cell_1866_a_HPC2_and_p_0_out_1__0_,
         cell_1866_a_HPC2_and_p_1_out_0__1_,
         cell_1866_a_HPC2_and_p_1_out_1__0_,
         cell_1866_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1866_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1866_a_HPC2_and_p_1_in_0__1_, cell_1866_a_HPC2_and_p_1_in_1__0_,
         cell_1866_a_HPC2_and_s_out_0__1_, cell_1866_a_HPC2_and_s_out_1__0_,
         cell_1866_a_HPC2_and_p_0_in_0__1_, cell_1866_a_HPC2_and_p_0_in_1__0_,
         cell_1866_a_HPC2_and_s_in_0__1_, cell_1866_a_HPC2_and_s_in_1__0_,
         cell_1866_a_HPC2_and_z_0__0_, cell_1866_a_HPC2_and_z_1__1_,
         cell_1867_a_HPC2_and_n9, cell_1867_a_HPC2_and_n8,
         cell_1867_a_HPC2_and_n7, cell_1867_a_HPC2_and_p_0_out_0__1_,
         cell_1867_a_HPC2_and_p_0_out_1__0_,
         cell_1867_a_HPC2_and_p_1_out_0__1_,
         cell_1867_a_HPC2_and_p_1_out_1__0_,
         cell_1867_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1867_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1867_a_HPC2_and_p_1_in_0__1_, cell_1867_a_HPC2_and_p_1_in_1__0_,
         cell_1867_a_HPC2_and_s_out_0__1_, cell_1867_a_HPC2_and_s_out_1__0_,
         cell_1867_a_HPC2_and_p_0_in_0__1_, cell_1867_a_HPC2_and_p_0_in_1__0_,
         cell_1867_a_HPC2_and_s_in_0__1_, cell_1867_a_HPC2_and_s_in_1__0_,
         cell_1867_a_HPC2_and_z_0__0_, cell_1867_a_HPC2_and_z_1__1_,
         cell_1868_a_HPC2_and_n9, cell_1868_a_HPC2_and_n8,
         cell_1868_a_HPC2_and_n7, cell_1868_a_HPC2_and_p_0_out_0__1_,
         cell_1868_a_HPC2_and_p_0_out_1__0_,
         cell_1868_a_HPC2_and_p_1_out_0__1_,
         cell_1868_a_HPC2_and_p_1_out_1__0_,
         cell_1868_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1868_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1868_a_HPC2_and_p_1_in_0__1_, cell_1868_a_HPC2_and_p_1_in_1__0_,
         cell_1868_a_HPC2_and_s_out_0__1_, cell_1868_a_HPC2_and_s_out_1__0_,
         cell_1868_a_HPC2_and_p_0_in_0__1_, cell_1868_a_HPC2_and_p_0_in_1__0_,
         cell_1868_a_HPC2_and_s_in_0__1_, cell_1868_a_HPC2_and_s_in_1__0_,
         cell_1868_a_HPC2_and_z_0__0_, cell_1868_a_HPC2_and_z_1__1_,
         cell_1869_a_HPC2_and_n9, cell_1869_a_HPC2_and_n8,
         cell_1869_a_HPC2_and_n7, cell_1869_a_HPC2_and_p_0_out_0__1_,
         cell_1869_a_HPC2_and_p_0_out_1__0_,
         cell_1869_a_HPC2_and_p_1_out_0__1_,
         cell_1869_a_HPC2_and_p_1_out_1__0_,
         cell_1869_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1869_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1869_a_HPC2_and_p_1_in_0__1_, cell_1869_a_HPC2_and_p_1_in_1__0_,
         cell_1869_a_HPC2_and_s_out_0__1_, cell_1869_a_HPC2_and_s_out_1__0_,
         cell_1869_a_HPC2_and_p_0_in_0__1_, cell_1869_a_HPC2_and_p_0_in_1__0_,
         cell_1869_a_HPC2_and_s_in_0__1_, cell_1869_a_HPC2_and_s_in_1__0_,
         cell_1869_a_HPC2_and_z_0__0_, cell_1869_a_HPC2_and_z_1__1_,
         cell_1870_a_HPC2_and_n9, cell_1870_a_HPC2_and_n8,
         cell_1870_a_HPC2_and_n7, cell_1870_a_HPC2_and_p_0_out_0__1_,
         cell_1870_a_HPC2_and_p_0_out_1__0_,
         cell_1870_a_HPC2_and_p_1_out_0__1_,
         cell_1870_a_HPC2_and_p_1_out_1__0_,
         cell_1870_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1870_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1870_a_HPC2_and_p_1_in_0__1_, cell_1870_a_HPC2_and_p_1_in_1__0_,
         cell_1870_a_HPC2_and_s_out_0__1_, cell_1870_a_HPC2_and_s_out_1__0_,
         cell_1870_a_HPC2_and_p_0_in_0__1_, cell_1870_a_HPC2_and_p_0_in_1__0_,
         cell_1870_a_HPC2_and_s_in_0__1_, cell_1870_a_HPC2_and_s_in_1__0_,
         cell_1870_a_HPC2_and_z_0__0_, cell_1870_a_HPC2_and_z_1__1_,
         cell_1871_a_HPC2_and_n9, cell_1871_a_HPC2_and_n8,
         cell_1871_a_HPC2_and_n7, cell_1871_a_HPC2_and_p_0_out_0__1_,
         cell_1871_a_HPC2_and_p_0_out_1__0_,
         cell_1871_a_HPC2_and_p_1_out_0__1_,
         cell_1871_a_HPC2_and_p_1_out_1__0_,
         cell_1871_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1871_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1871_a_HPC2_and_p_1_in_0__1_, cell_1871_a_HPC2_and_p_1_in_1__0_,
         cell_1871_a_HPC2_and_s_out_0__1_, cell_1871_a_HPC2_and_s_out_1__0_,
         cell_1871_a_HPC2_and_p_0_in_0__1_, cell_1871_a_HPC2_and_p_0_in_1__0_,
         cell_1871_a_HPC2_and_s_in_0__1_, cell_1871_a_HPC2_and_s_in_1__0_,
         cell_1871_a_HPC2_and_z_0__0_, cell_1871_a_HPC2_and_z_1__1_,
         cell_1872_a_HPC2_and_n9, cell_1872_a_HPC2_and_n8,
         cell_1872_a_HPC2_and_n7, cell_1872_a_HPC2_and_p_0_out_0__1_,
         cell_1872_a_HPC2_and_p_0_out_1__0_,
         cell_1872_a_HPC2_and_p_1_out_0__1_,
         cell_1872_a_HPC2_and_p_1_out_1__0_,
         cell_1872_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1872_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1872_a_HPC2_and_p_1_in_0__1_, cell_1872_a_HPC2_and_p_1_in_1__0_,
         cell_1872_a_HPC2_and_s_out_0__1_, cell_1872_a_HPC2_and_s_out_1__0_,
         cell_1872_a_HPC2_and_p_0_in_0__1_, cell_1872_a_HPC2_and_p_0_in_1__0_,
         cell_1872_a_HPC2_and_s_in_0__1_, cell_1872_a_HPC2_and_s_in_1__0_,
         cell_1872_a_HPC2_and_z_0__0_, cell_1872_a_HPC2_and_z_1__1_,
         cell_1873_a_HPC2_and_n9, cell_1873_a_HPC2_and_n8,
         cell_1873_a_HPC2_and_n7, cell_1873_a_HPC2_and_p_0_out_0__1_,
         cell_1873_a_HPC2_and_p_0_out_1__0_,
         cell_1873_a_HPC2_and_p_1_out_0__1_,
         cell_1873_a_HPC2_and_p_1_out_1__0_,
         cell_1873_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1873_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1873_a_HPC2_and_p_1_in_0__1_, cell_1873_a_HPC2_and_p_1_in_1__0_,
         cell_1873_a_HPC2_and_s_out_0__1_, cell_1873_a_HPC2_and_s_out_1__0_,
         cell_1873_a_HPC2_and_p_0_in_0__1_, cell_1873_a_HPC2_and_p_0_in_1__0_,
         cell_1873_a_HPC2_and_s_in_0__1_, cell_1873_a_HPC2_and_s_in_1__0_,
         cell_1873_a_HPC2_and_z_0__0_, cell_1873_a_HPC2_and_z_1__1_,
         cell_1874_a_HPC2_and_n9, cell_1874_a_HPC2_and_n8,
         cell_1874_a_HPC2_and_n7, cell_1874_a_HPC2_and_p_0_out_0__1_,
         cell_1874_a_HPC2_and_p_0_out_1__0_,
         cell_1874_a_HPC2_and_p_1_out_0__1_,
         cell_1874_a_HPC2_and_p_1_out_1__0_,
         cell_1874_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1874_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1874_a_HPC2_and_p_1_in_0__1_, cell_1874_a_HPC2_and_p_1_in_1__0_,
         cell_1874_a_HPC2_and_s_out_0__1_, cell_1874_a_HPC2_and_s_out_1__0_,
         cell_1874_a_HPC2_and_p_0_in_0__1_, cell_1874_a_HPC2_and_p_0_in_1__0_,
         cell_1874_a_HPC2_and_s_in_0__1_, cell_1874_a_HPC2_and_s_in_1__0_,
         cell_1874_a_HPC2_and_z_0__0_, cell_1874_a_HPC2_and_z_1__1_,
         cell_1875_a_HPC2_and_n9, cell_1875_a_HPC2_and_n8,
         cell_1875_a_HPC2_and_n7, cell_1875_a_HPC2_and_p_0_out_0__1_,
         cell_1875_a_HPC2_and_p_0_out_1__0_,
         cell_1875_a_HPC2_and_p_1_out_0__1_,
         cell_1875_a_HPC2_and_p_1_out_1__0_,
         cell_1875_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1875_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1875_a_HPC2_and_p_1_in_0__1_, cell_1875_a_HPC2_and_p_1_in_1__0_,
         cell_1875_a_HPC2_and_s_out_0__1_, cell_1875_a_HPC2_and_s_out_1__0_,
         cell_1875_a_HPC2_and_p_0_in_0__1_, cell_1875_a_HPC2_and_p_0_in_1__0_,
         cell_1875_a_HPC2_and_s_in_0__1_, cell_1875_a_HPC2_and_s_in_1__0_,
         cell_1875_a_HPC2_and_z_0__0_, cell_1875_a_HPC2_and_z_1__1_,
         cell_1876_a_HPC2_and_n9, cell_1876_a_HPC2_and_n8,
         cell_1876_a_HPC2_and_n7, cell_1876_a_HPC2_and_p_0_out_0__1_,
         cell_1876_a_HPC2_and_p_0_out_1__0_,
         cell_1876_a_HPC2_and_p_1_out_0__1_,
         cell_1876_a_HPC2_and_p_1_out_1__0_,
         cell_1876_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1876_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1876_a_HPC2_and_p_1_in_0__1_, cell_1876_a_HPC2_and_p_1_in_1__0_,
         cell_1876_a_HPC2_and_s_out_0__1_, cell_1876_a_HPC2_and_s_out_1__0_,
         cell_1876_a_HPC2_and_p_0_in_0__1_, cell_1876_a_HPC2_and_p_0_in_1__0_,
         cell_1876_a_HPC2_and_s_in_0__1_, cell_1876_a_HPC2_and_s_in_1__0_,
         cell_1876_a_HPC2_and_z_0__0_, cell_1876_a_HPC2_and_z_1__1_,
         cell_1877_a_HPC2_and_n9, cell_1877_a_HPC2_and_n8,
         cell_1877_a_HPC2_and_n7, cell_1877_a_HPC2_and_p_0_out_0__1_,
         cell_1877_a_HPC2_and_p_0_out_1__0_,
         cell_1877_a_HPC2_and_p_1_out_0__1_,
         cell_1877_a_HPC2_and_p_1_out_1__0_,
         cell_1877_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1877_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1877_a_HPC2_and_p_1_in_0__1_, cell_1877_a_HPC2_and_p_1_in_1__0_,
         cell_1877_a_HPC2_and_s_out_0__1_, cell_1877_a_HPC2_and_s_out_1__0_,
         cell_1877_a_HPC2_and_p_0_in_0__1_, cell_1877_a_HPC2_and_p_0_in_1__0_,
         cell_1877_a_HPC2_and_s_in_0__1_, cell_1877_a_HPC2_and_s_in_1__0_,
         cell_1877_a_HPC2_and_z_0__0_, cell_1877_a_HPC2_and_z_1__1_,
         cell_1878_a_HPC2_and_n9, cell_1878_a_HPC2_and_n8,
         cell_1878_a_HPC2_and_n7, cell_1878_a_HPC2_and_p_0_out_0__1_,
         cell_1878_a_HPC2_and_p_0_out_1__0_,
         cell_1878_a_HPC2_and_p_1_out_0__1_,
         cell_1878_a_HPC2_and_p_1_out_1__0_,
         cell_1878_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1878_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1878_a_HPC2_and_p_1_in_0__1_, cell_1878_a_HPC2_and_p_1_in_1__0_,
         cell_1878_a_HPC2_and_s_out_0__1_, cell_1878_a_HPC2_and_s_out_1__0_,
         cell_1878_a_HPC2_and_p_0_in_0__1_, cell_1878_a_HPC2_and_p_0_in_1__0_,
         cell_1878_a_HPC2_and_s_in_0__1_, cell_1878_a_HPC2_and_s_in_1__0_,
         cell_1878_a_HPC2_and_z_0__0_, cell_1878_a_HPC2_and_z_1__1_,
         cell_1879_a_HPC2_and_n9, cell_1879_a_HPC2_and_n8,
         cell_1879_a_HPC2_and_n7, cell_1879_a_HPC2_and_p_0_out_0__1_,
         cell_1879_a_HPC2_and_p_0_out_1__0_,
         cell_1879_a_HPC2_and_p_1_out_0__1_,
         cell_1879_a_HPC2_and_p_1_out_1__0_,
         cell_1879_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1879_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1879_a_HPC2_and_p_1_in_0__1_, cell_1879_a_HPC2_and_p_1_in_1__0_,
         cell_1879_a_HPC2_and_s_out_0__1_, cell_1879_a_HPC2_and_s_out_1__0_,
         cell_1879_a_HPC2_and_p_0_in_0__1_, cell_1879_a_HPC2_and_p_0_in_1__0_,
         cell_1879_a_HPC2_and_s_in_0__1_, cell_1879_a_HPC2_and_s_in_1__0_,
         cell_1879_a_HPC2_and_z_0__0_, cell_1879_a_HPC2_and_z_1__1_,
         cell_1880_a_HPC2_and_n9, cell_1880_a_HPC2_and_n8,
         cell_1880_a_HPC2_and_n7, cell_1880_a_HPC2_and_p_0_out_0__1_,
         cell_1880_a_HPC2_and_p_0_out_1__0_,
         cell_1880_a_HPC2_and_p_1_out_0__1_,
         cell_1880_a_HPC2_and_p_1_out_1__0_,
         cell_1880_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1880_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1880_a_HPC2_and_p_1_in_0__1_, cell_1880_a_HPC2_and_p_1_in_1__0_,
         cell_1880_a_HPC2_and_s_out_0__1_, cell_1880_a_HPC2_and_s_out_1__0_,
         cell_1880_a_HPC2_and_p_0_in_0__1_, cell_1880_a_HPC2_and_p_0_in_1__0_,
         cell_1880_a_HPC2_and_s_in_0__1_, cell_1880_a_HPC2_and_s_in_1__0_,
         cell_1880_a_HPC2_and_z_0__0_, cell_1880_a_HPC2_and_z_1__1_,
         cell_1881_a_HPC2_and_n9, cell_1881_a_HPC2_and_n8,
         cell_1881_a_HPC2_and_n7, cell_1881_a_HPC2_and_p_0_out_0__1_,
         cell_1881_a_HPC2_and_p_0_out_1__0_,
         cell_1881_a_HPC2_and_p_1_out_0__1_,
         cell_1881_a_HPC2_and_p_1_out_1__0_,
         cell_1881_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1881_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1881_a_HPC2_and_p_1_in_0__1_, cell_1881_a_HPC2_and_p_1_in_1__0_,
         cell_1881_a_HPC2_and_s_out_0__1_, cell_1881_a_HPC2_and_s_out_1__0_,
         cell_1881_a_HPC2_and_p_0_in_0__1_, cell_1881_a_HPC2_and_p_0_in_1__0_,
         cell_1881_a_HPC2_and_s_in_0__1_, cell_1881_a_HPC2_and_s_in_1__0_,
         cell_1881_a_HPC2_and_z_0__0_, cell_1881_a_HPC2_and_z_1__1_,
         cell_1882_a_HPC2_and_n9, cell_1882_a_HPC2_and_n8,
         cell_1882_a_HPC2_and_n7, cell_1882_a_HPC2_and_p_0_out_0__1_,
         cell_1882_a_HPC2_and_p_0_out_1__0_,
         cell_1882_a_HPC2_and_p_1_out_0__1_,
         cell_1882_a_HPC2_and_p_1_out_1__0_,
         cell_1882_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1882_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1882_a_HPC2_and_p_1_in_0__1_, cell_1882_a_HPC2_and_p_1_in_1__0_,
         cell_1882_a_HPC2_and_s_out_0__1_, cell_1882_a_HPC2_and_s_out_1__0_,
         cell_1882_a_HPC2_and_p_0_in_0__1_, cell_1882_a_HPC2_and_p_0_in_1__0_,
         cell_1882_a_HPC2_and_s_in_0__1_, cell_1882_a_HPC2_and_s_in_1__0_,
         cell_1882_a_HPC2_and_z_0__0_, cell_1882_a_HPC2_and_z_1__1_,
         cell_1883_a_HPC2_and_n9, cell_1883_a_HPC2_and_n8,
         cell_1883_a_HPC2_and_n7, cell_1883_a_HPC2_and_p_0_out_0__1_,
         cell_1883_a_HPC2_and_p_0_out_1__0_,
         cell_1883_a_HPC2_and_p_1_out_0__1_,
         cell_1883_a_HPC2_and_p_1_out_1__0_,
         cell_1883_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1883_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1883_a_HPC2_and_p_1_in_0__1_, cell_1883_a_HPC2_and_p_1_in_1__0_,
         cell_1883_a_HPC2_and_s_out_0__1_, cell_1883_a_HPC2_and_s_out_1__0_,
         cell_1883_a_HPC2_and_p_0_in_0__1_, cell_1883_a_HPC2_and_p_0_in_1__0_,
         cell_1883_a_HPC2_and_s_in_0__1_, cell_1883_a_HPC2_and_s_in_1__0_,
         cell_1883_a_HPC2_and_z_0__0_, cell_1883_a_HPC2_and_z_1__1_,
         cell_1884_a_HPC2_and_n9, cell_1884_a_HPC2_and_n8,
         cell_1884_a_HPC2_and_n7, cell_1884_a_HPC2_and_p_0_out_0__1_,
         cell_1884_a_HPC2_and_p_0_out_1__0_,
         cell_1884_a_HPC2_and_p_1_out_0__1_,
         cell_1884_a_HPC2_and_p_1_out_1__0_,
         cell_1884_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1884_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1884_a_HPC2_and_p_1_in_0__1_, cell_1884_a_HPC2_and_p_1_in_1__0_,
         cell_1884_a_HPC2_and_s_out_0__1_, cell_1884_a_HPC2_and_s_out_1__0_,
         cell_1884_a_HPC2_and_p_0_in_0__1_, cell_1884_a_HPC2_and_p_0_in_1__0_,
         cell_1884_a_HPC2_and_s_in_0__1_, cell_1884_a_HPC2_and_s_in_1__0_,
         cell_1884_a_HPC2_and_z_0__0_, cell_1884_a_HPC2_and_z_1__1_,
         cell_1885_a_HPC2_and_n9, cell_1885_a_HPC2_and_n8,
         cell_1885_a_HPC2_and_n7, cell_1885_a_HPC2_and_p_0_out_0__1_,
         cell_1885_a_HPC2_and_p_0_out_1__0_,
         cell_1885_a_HPC2_and_p_1_out_0__1_,
         cell_1885_a_HPC2_and_p_1_out_1__0_,
         cell_1885_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1885_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1885_a_HPC2_and_p_1_in_0__1_, cell_1885_a_HPC2_and_p_1_in_1__0_,
         cell_1885_a_HPC2_and_s_out_0__1_, cell_1885_a_HPC2_and_s_out_1__0_,
         cell_1885_a_HPC2_and_p_0_in_0__1_, cell_1885_a_HPC2_and_p_0_in_1__0_,
         cell_1885_a_HPC2_and_s_in_0__1_, cell_1885_a_HPC2_and_s_in_1__0_,
         cell_1885_a_HPC2_and_z_0__0_, cell_1885_a_HPC2_and_z_1__1_,
         cell_1886_a_HPC2_and_n9, cell_1886_a_HPC2_and_n8,
         cell_1886_a_HPC2_and_n7, cell_1886_a_HPC2_and_p_0_out_0__1_,
         cell_1886_a_HPC2_and_p_0_out_1__0_,
         cell_1886_a_HPC2_and_p_1_out_0__1_,
         cell_1886_a_HPC2_and_p_1_out_1__0_,
         cell_1886_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1886_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1886_a_HPC2_and_p_1_in_0__1_, cell_1886_a_HPC2_and_p_1_in_1__0_,
         cell_1886_a_HPC2_and_s_out_0__1_, cell_1886_a_HPC2_and_s_out_1__0_,
         cell_1886_a_HPC2_and_p_0_in_0__1_, cell_1886_a_HPC2_and_p_0_in_1__0_,
         cell_1886_a_HPC2_and_s_in_0__1_, cell_1886_a_HPC2_and_s_in_1__0_,
         cell_1886_a_HPC2_and_z_0__0_, cell_1886_a_HPC2_and_z_1__1_,
         cell_1887_a_HPC2_and_n9, cell_1887_a_HPC2_and_n8,
         cell_1887_a_HPC2_and_n7, cell_1887_a_HPC2_and_p_0_out_0__1_,
         cell_1887_a_HPC2_and_p_0_out_1__0_,
         cell_1887_a_HPC2_and_p_1_out_0__1_,
         cell_1887_a_HPC2_and_p_1_out_1__0_,
         cell_1887_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1887_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1887_a_HPC2_and_p_1_in_0__1_, cell_1887_a_HPC2_and_p_1_in_1__0_,
         cell_1887_a_HPC2_and_s_out_0__1_, cell_1887_a_HPC2_and_s_out_1__0_,
         cell_1887_a_HPC2_and_p_0_in_0__1_, cell_1887_a_HPC2_and_p_0_in_1__0_,
         cell_1887_a_HPC2_and_s_in_0__1_, cell_1887_a_HPC2_and_s_in_1__0_,
         cell_1887_a_HPC2_and_z_0__0_, cell_1887_a_HPC2_and_z_1__1_,
         cell_1888_a_HPC2_and_n9, cell_1888_a_HPC2_and_n8,
         cell_1888_a_HPC2_and_n7, cell_1888_a_HPC2_and_p_0_out_0__1_,
         cell_1888_a_HPC2_and_p_0_out_1__0_,
         cell_1888_a_HPC2_and_p_1_out_0__1_,
         cell_1888_a_HPC2_and_p_1_out_1__0_,
         cell_1888_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1888_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1888_a_HPC2_and_p_1_in_0__1_, cell_1888_a_HPC2_and_p_1_in_1__0_,
         cell_1888_a_HPC2_and_s_out_0__1_, cell_1888_a_HPC2_and_s_out_1__0_,
         cell_1888_a_HPC2_and_p_0_in_0__1_, cell_1888_a_HPC2_and_p_0_in_1__0_,
         cell_1888_a_HPC2_and_s_in_0__1_, cell_1888_a_HPC2_and_s_in_1__0_,
         cell_1888_a_HPC2_and_z_0__0_, cell_1888_a_HPC2_and_z_1__1_,
         cell_1889_a_HPC2_and_n9, cell_1889_a_HPC2_and_n8,
         cell_1889_a_HPC2_and_n7, cell_1889_a_HPC2_and_p_0_out_0__1_,
         cell_1889_a_HPC2_and_p_0_out_1__0_,
         cell_1889_a_HPC2_and_p_1_out_0__1_,
         cell_1889_a_HPC2_and_p_1_out_1__0_,
         cell_1889_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1889_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1889_a_HPC2_and_p_1_in_0__1_, cell_1889_a_HPC2_and_p_1_in_1__0_,
         cell_1889_a_HPC2_and_s_out_0__1_, cell_1889_a_HPC2_and_s_out_1__0_,
         cell_1889_a_HPC2_and_p_0_in_0__1_, cell_1889_a_HPC2_and_p_0_in_1__0_,
         cell_1889_a_HPC2_and_s_in_0__1_, cell_1889_a_HPC2_and_s_in_1__0_,
         cell_1889_a_HPC2_and_z_0__0_, cell_1889_a_HPC2_and_z_1__1_,
         cell_1890_a_HPC2_and_n9, cell_1890_a_HPC2_and_n8,
         cell_1890_a_HPC2_and_n7, cell_1890_a_HPC2_and_p_0_out_0__1_,
         cell_1890_a_HPC2_and_p_0_out_1__0_,
         cell_1890_a_HPC2_and_p_1_out_0__1_,
         cell_1890_a_HPC2_and_p_1_out_1__0_,
         cell_1890_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1890_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1890_a_HPC2_and_p_1_in_0__1_, cell_1890_a_HPC2_and_p_1_in_1__0_,
         cell_1890_a_HPC2_and_s_out_0__1_, cell_1890_a_HPC2_and_s_out_1__0_,
         cell_1890_a_HPC2_and_p_0_in_0__1_, cell_1890_a_HPC2_and_p_0_in_1__0_,
         cell_1890_a_HPC2_and_s_in_0__1_, cell_1890_a_HPC2_and_s_in_1__0_,
         cell_1890_a_HPC2_and_z_0__0_, cell_1890_a_HPC2_and_z_1__1_,
         cell_1891_a_HPC2_and_n9, cell_1891_a_HPC2_and_n8,
         cell_1891_a_HPC2_and_n7, cell_1891_a_HPC2_and_p_0_out_0__1_,
         cell_1891_a_HPC2_and_p_0_out_1__0_,
         cell_1891_a_HPC2_and_p_1_out_0__1_,
         cell_1891_a_HPC2_and_p_1_out_1__0_,
         cell_1891_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1891_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1891_a_HPC2_and_p_1_in_0__1_, cell_1891_a_HPC2_and_p_1_in_1__0_,
         cell_1891_a_HPC2_and_s_out_0__1_, cell_1891_a_HPC2_and_s_out_1__0_,
         cell_1891_a_HPC2_and_p_0_in_0__1_, cell_1891_a_HPC2_and_p_0_in_1__0_,
         cell_1891_a_HPC2_and_s_in_0__1_, cell_1891_a_HPC2_and_s_in_1__0_,
         cell_1891_a_HPC2_and_z_0__0_, cell_1891_a_HPC2_and_z_1__1_,
         cell_1892_a_HPC2_and_n9, cell_1892_a_HPC2_and_n8,
         cell_1892_a_HPC2_and_n7, cell_1892_a_HPC2_and_p_0_out_0__1_,
         cell_1892_a_HPC2_and_p_0_out_1__0_,
         cell_1892_a_HPC2_and_p_1_out_0__1_,
         cell_1892_a_HPC2_and_p_1_out_1__0_,
         cell_1892_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1892_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1892_a_HPC2_and_p_1_in_0__1_, cell_1892_a_HPC2_and_p_1_in_1__0_,
         cell_1892_a_HPC2_and_s_out_0__1_, cell_1892_a_HPC2_and_s_out_1__0_,
         cell_1892_a_HPC2_and_p_0_in_0__1_, cell_1892_a_HPC2_and_p_0_in_1__0_,
         cell_1892_a_HPC2_and_s_in_0__1_, cell_1892_a_HPC2_and_s_in_1__0_,
         cell_1892_a_HPC2_and_z_0__0_, cell_1892_a_HPC2_and_z_1__1_,
         cell_1893_a_HPC2_and_n9, cell_1893_a_HPC2_and_n8,
         cell_1893_a_HPC2_and_n7, cell_1893_a_HPC2_and_p_0_out_0__1_,
         cell_1893_a_HPC2_and_p_0_out_1__0_,
         cell_1893_a_HPC2_and_p_1_out_0__1_,
         cell_1893_a_HPC2_and_p_1_out_1__0_,
         cell_1893_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1893_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1893_a_HPC2_and_p_1_in_0__1_, cell_1893_a_HPC2_and_p_1_in_1__0_,
         cell_1893_a_HPC2_and_s_out_0__1_, cell_1893_a_HPC2_and_s_out_1__0_,
         cell_1893_a_HPC2_and_p_0_in_0__1_, cell_1893_a_HPC2_and_p_0_in_1__0_,
         cell_1893_a_HPC2_and_s_in_0__1_, cell_1893_a_HPC2_and_s_in_1__0_,
         cell_1893_a_HPC2_and_z_0__0_, cell_1893_a_HPC2_and_z_1__1_,
         cell_1894_a_HPC2_and_n9, cell_1894_a_HPC2_and_n8,
         cell_1894_a_HPC2_and_n7, cell_1894_a_HPC2_and_p_0_out_0__1_,
         cell_1894_a_HPC2_and_p_0_out_1__0_,
         cell_1894_a_HPC2_and_p_1_out_0__1_,
         cell_1894_a_HPC2_and_p_1_out_1__0_,
         cell_1894_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1894_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1894_a_HPC2_and_p_1_in_0__1_, cell_1894_a_HPC2_and_p_1_in_1__0_,
         cell_1894_a_HPC2_and_s_out_0__1_, cell_1894_a_HPC2_and_s_out_1__0_,
         cell_1894_a_HPC2_and_p_0_in_0__1_, cell_1894_a_HPC2_and_p_0_in_1__0_,
         cell_1894_a_HPC2_and_s_in_0__1_, cell_1894_a_HPC2_and_s_in_1__0_,
         cell_1894_a_HPC2_and_z_0__0_, cell_1894_a_HPC2_and_z_1__1_,
         cell_1895_a_HPC2_and_n9, cell_1895_a_HPC2_and_n8,
         cell_1895_a_HPC2_and_n7, cell_1895_a_HPC2_and_p_0_out_0__1_,
         cell_1895_a_HPC2_and_p_0_out_1__0_,
         cell_1895_a_HPC2_and_p_1_out_0__1_,
         cell_1895_a_HPC2_and_p_1_out_1__0_,
         cell_1895_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1895_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1895_a_HPC2_and_p_1_in_0__1_, cell_1895_a_HPC2_and_p_1_in_1__0_,
         cell_1895_a_HPC2_and_s_out_0__1_, cell_1895_a_HPC2_and_s_out_1__0_,
         cell_1895_a_HPC2_and_p_0_in_0__1_, cell_1895_a_HPC2_and_p_0_in_1__0_,
         cell_1895_a_HPC2_and_s_in_0__1_, cell_1895_a_HPC2_and_s_in_1__0_,
         cell_1895_a_HPC2_and_z_0__0_, cell_1895_a_HPC2_and_z_1__1_,
         cell_1896_a_HPC2_and_n9, cell_1896_a_HPC2_and_n8,
         cell_1896_a_HPC2_and_n7, cell_1896_a_HPC2_and_p_0_out_0__1_,
         cell_1896_a_HPC2_and_p_0_out_1__0_,
         cell_1896_a_HPC2_and_p_1_out_0__1_,
         cell_1896_a_HPC2_and_p_1_out_1__0_,
         cell_1896_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1896_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1896_a_HPC2_and_p_1_in_0__1_, cell_1896_a_HPC2_and_p_1_in_1__0_,
         cell_1896_a_HPC2_and_s_out_0__1_, cell_1896_a_HPC2_and_s_out_1__0_,
         cell_1896_a_HPC2_and_p_0_in_0__1_, cell_1896_a_HPC2_and_p_0_in_1__0_,
         cell_1896_a_HPC2_and_s_in_0__1_, cell_1896_a_HPC2_and_s_in_1__0_,
         cell_1896_a_HPC2_and_z_0__0_, cell_1896_a_HPC2_and_z_1__1_,
         cell_1897_a_HPC2_and_n9, cell_1897_a_HPC2_and_n8,
         cell_1897_a_HPC2_and_n7, cell_1897_a_HPC2_and_p_0_out_0__1_,
         cell_1897_a_HPC2_and_p_0_out_1__0_,
         cell_1897_a_HPC2_and_p_1_out_0__1_,
         cell_1897_a_HPC2_and_p_1_out_1__0_,
         cell_1897_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1897_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1897_a_HPC2_and_p_1_in_0__1_, cell_1897_a_HPC2_and_p_1_in_1__0_,
         cell_1897_a_HPC2_and_s_out_0__1_, cell_1897_a_HPC2_and_s_out_1__0_,
         cell_1897_a_HPC2_and_p_0_in_0__1_, cell_1897_a_HPC2_and_p_0_in_1__0_,
         cell_1897_a_HPC2_and_s_in_0__1_, cell_1897_a_HPC2_and_s_in_1__0_,
         cell_1897_a_HPC2_and_z_0__0_, cell_1897_a_HPC2_and_z_1__1_,
         cell_1898_a_HPC2_and_n9, cell_1898_a_HPC2_and_n8,
         cell_1898_a_HPC2_and_n7, cell_1898_a_HPC2_and_p_0_out_0__1_,
         cell_1898_a_HPC2_and_p_0_out_1__0_,
         cell_1898_a_HPC2_and_p_1_out_0__1_,
         cell_1898_a_HPC2_and_p_1_out_1__0_,
         cell_1898_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1898_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1898_a_HPC2_and_p_1_in_0__1_, cell_1898_a_HPC2_and_p_1_in_1__0_,
         cell_1898_a_HPC2_and_s_out_0__1_, cell_1898_a_HPC2_and_s_out_1__0_,
         cell_1898_a_HPC2_and_p_0_in_0__1_, cell_1898_a_HPC2_and_p_0_in_1__0_,
         cell_1898_a_HPC2_and_s_in_0__1_, cell_1898_a_HPC2_and_s_in_1__0_,
         cell_1898_a_HPC2_and_z_0__0_, cell_1898_a_HPC2_and_z_1__1_,
         cell_1899_a_HPC2_and_n9, cell_1899_a_HPC2_and_n8,
         cell_1899_a_HPC2_and_n7, cell_1899_a_HPC2_and_p_0_out_0__1_,
         cell_1899_a_HPC2_and_p_0_out_1__0_,
         cell_1899_a_HPC2_and_p_1_out_0__1_,
         cell_1899_a_HPC2_and_p_1_out_1__0_,
         cell_1899_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1899_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1899_a_HPC2_and_p_1_in_0__1_, cell_1899_a_HPC2_and_p_1_in_1__0_,
         cell_1899_a_HPC2_and_s_out_0__1_, cell_1899_a_HPC2_and_s_out_1__0_,
         cell_1899_a_HPC2_and_p_0_in_0__1_, cell_1899_a_HPC2_and_p_0_in_1__0_,
         cell_1899_a_HPC2_and_s_in_0__1_, cell_1899_a_HPC2_and_s_in_1__0_,
         cell_1899_a_HPC2_and_z_0__0_, cell_1899_a_HPC2_and_z_1__1_,
         cell_1900_a_HPC2_and_n9, cell_1900_a_HPC2_and_n8,
         cell_1900_a_HPC2_and_n7, cell_1900_a_HPC2_and_p_0_out_0__1_,
         cell_1900_a_HPC2_and_p_0_out_1__0_,
         cell_1900_a_HPC2_and_p_1_out_0__1_,
         cell_1900_a_HPC2_and_p_1_out_1__0_,
         cell_1900_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1900_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1900_a_HPC2_and_p_1_in_0__1_, cell_1900_a_HPC2_and_p_1_in_1__0_,
         cell_1900_a_HPC2_and_s_out_0__1_, cell_1900_a_HPC2_and_s_out_1__0_,
         cell_1900_a_HPC2_and_p_0_in_0__1_, cell_1900_a_HPC2_and_p_0_in_1__0_,
         cell_1900_a_HPC2_and_s_in_0__1_, cell_1900_a_HPC2_and_s_in_1__0_,
         cell_1900_a_HPC2_and_z_0__0_, cell_1900_a_HPC2_and_z_1__1_,
         cell_1901_a_HPC2_and_n9, cell_1901_a_HPC2_and_n8,
         cell_1901_a_HPC2_and_n7, cell_1901_a_HPC2_and_p_0_out_0__1_,
         cell_1901_a_HPC2_and_p_0_out_1__0_,
         cell_1901_a_HPC2_and_p_1_out_0__1_,
         cell_1901_a_HPC2_and_p_1_out_1__0_,
         cell_1901_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1901_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1901_a_HPC2_and_p_1_in_0__1_, cell_1901_a_HPC2_and_p_1_in_1__0_,
         cell_1901_a_HPC2_and_s_out_0__1_, cell_1901_a_HPC2_and_s_out_1__0_,
         cell_1901_a_HPC2_and_p_0_in_0__1_, cell_1901_a_HPC2_and_p_0_in_1__0_,
         cell_1901_a_HPC2_and_s_in_0__1_, cell_1901_a_HPC2_and_s_in_1__0_,
         cell_1901_a_HPC2_and_z_0__0_, cell_1901_a_HPC2_and_z_1__1_,
         cell_1902_a_HPC2_and_n9, cell_1902_a_HPC2_and_n8,
         cell_1902_a_HPC2_and_n7, cell_1902_a_HPC2_and_p_0_out_0__1_,
         cell_1902_a_HPC2_and_p_0_out_1__0_,
         cell_1902_a_HPC2_and_p_1_out_0__1_,
         cell_1902_a_HPC2_and_p_1_out_1__0_,
         cell_1902_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1902_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1902_a_HPC2_and_p_1_in_0__1_, cell_1902_a_HPC2_and_p_1_in_1__0_,
         cell_1902_a_HPC2_and_s_out_0__1_, cell_1902_a_HPC2_and_s_out_1__0_,
         cell_1902_a_HPC2_and_p_0_in_0__1_, cell_1902_a_HPC2_and_p_0_in_1__0_,
         cell_1902_a_HPC2_and_s_in_0__1_, cell_1902_a_HPC2_and_s_in_1__0_,
         cell_1902_a_HPC2_and_z_0__0_, cell_1902_a_HPC2_and_z_1__1_,
         cell_1903_a_HPC2_and_n9, cell_1903_a_HPC2_and_n8,
         cell_1903_a_HPC2_and_n7, cell_1903_a_HPC2_and_p_0_out_0__1_,
         cell_1903_a_HPC2_and_p_0_out_1__0_,
         cell_1903_a_HPC2_and_p_1_out_0__1_,
         cell_1903_a_HPC2_and_p_1_out_1__0_,
         cell_1903_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1903_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1903_a_HPC2_and_p_1_in_0__1_, cell_1903_a_HPC2_and_p_1_in_1__0_,
         cell_1903_a_HPC2_and_s_out_0__1_, cell_1903_a_HPC2_and_s_out_1__0_,
         cell_1903_a_HPC2_and_p_0_in_0__1_, cell_1903_a_HPC2_and_p_0_in_1__0_,
         cell_1903_a_HPC2_and_s_in_0__1_, cell_1903_a_HPC2_and_s_in_1__0_,
         cell_1903_a_HPC2_and_z_0__0_, cell_1903_a_HPC2_and_z_1__1_,
         cell_1904_a_HPC2_and_n9, cell_1904_a_HPC2_and_n8,
         cell_1904_a_HPC2_and_n7, cell_1904_a_HPC2_and_p_0_out_0__1_,
         cell_1904_a_HPC2_and_p_0_out_1__0_,
         cell_1904_a_HPC2_and_p_1_out_0__1_,
         cell_1904_a_HPC2_and_p_1_out_1__0_,
         cell_1904_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1904_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1904_a_HPC2_and_p_1_in_0__1_, cell_1904_a_HPC2_and_p_1_in_1__0_,
         cell_1904_a_HPC2_and_s_out_0__1_, cell_1904_a_HPC2_and_s_out_1__0_,
         cell_1904_a_HPC2_and_p_0_in_0__1_, cell_1904_a_HPC2_and_p_0_in_1__0_,
         cell_1904_a_HPC2_and_s_in_0__1_, cell_1904_a_HPC2_and_s_in_1__0_,
         cell_1904_a_HPC2_and_z_0__0_, cell_1904_a_HPC2_and_z_1__1_,
         cell_1905_a_HPC2_and_n9, cell_1905_a_HPC2_and_n8,
         cell_1905_a_HPC2_and_n7, cell_1905_a_HPC2_and_p_0_out_0__1_,
         cell_1905_a_HPC2_and_p_0_out_1__0_,
         cell_1905_a_HPC2_and_p_1_out_0__1_,
         cell_1905_a_HPC2_and_p_1_out_1__0_,
         cell_1905_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1905_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1905_a_HPC2_and_p_1_in_0__1_, cell_1905_a_HPC2_and_p_1_in_1__0_,
         cell_1905_a_HPC2_and_s_out_0__1_, cell_1905_a_HPC2_and_s_out_1__0_,
         cell_1905_a_HPC2_and_p_0_in_0__1_, cell_1905_a_HPC2_and_p_0_in_1__0_,
         cell_1905_a_HPC2_and_s_in_0__1_, cell_1905_a_HPC2_and_s_in_1__0_,
         cell_1905_a_HPC2_and_z_0__0_, cell_1905_a_HPC2_and_z_1__1_,
         cell_1906_a_HPC2_and_n9, cell_1906_a_HPC2_and_n8,
         cell_1906_a_HPC2_and_n7, cell_1906_a_HPC2_and_p_0_out_0__1_,
         cell_1906_a_HPC2_and_p_0_out_1__0_,
         cell_1906_a_HPC2_and_p_1_out_0__1_,
         cell_1906_a_HPC2_and_p_1_out_1__0_,
         cell_1906_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1906_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1906_a_HPC2_and_p_1_in_0__1_, cell_1906_a_HPC2_and_p_1_in_1__0_,
         cell_1906_a_HPC2_and_s_out_0__1_, cell_1906_a_HPC2_and_s_out_1__0_,
         cell_1906_a_HPC2_and_p_0_in_0__1_, cell_1906_a_HPC2_and_p_0_in_1__0_,
         cell_1906_a_HPC2_and_s_in_0__1_, cell_1906_a_HPC2_and_s_in_1__0_,
         cell_1906_a_HPC2_and_z_0__0_, cell_1906_a_HPC2_and_z_1__1_,
         cell_1907_a_HPC2_and_n9, cell_1907_a_HPC2_and_n8,
         cell_1907_a_HPC2_and_n7, cell_1907_a_HPC2_and_p_0_out_0__1_,
         cell_1907_a_HPC2_and_p_0_out_1__0_,
         cell_1907_a_HPC2_and_p_1_out_0__1_,
         cell_1907_a_HPC2_and_p_1_out_1__0_,
         cell_1907_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1907_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1907_a_HPC2_and_p_1_in_0__1_, cell_1907_a_HPC2_and_p_1_in_1__0_,
         cell_1907_a_HPC2_and_s_out_0__1_, cell_1907_a_HPC2_and_s_out_1__0_,
         cell_1907_a_HPC2_and_p_0_in_0__1_, cell_1907_a_HPC2_and_p_0_in_1__0_,
         cell_1907_a_HPC2_and_s_in_0__1_, cell_1907_a_HPC2_and_s_in_1__0_,
         cell_1907_a_HPC2_and_z_0__0_, cell_1907_a_HPC2_and_z_1__1_,
         cell_1908_a_HPC2_and_n9, cell_1908_a_HPC2_and_n8,
         cell_1908_a_HPC2_and_n7, cell_1908_a_HPC2_and_p_0_out_0__1_,
         cell_1908_a_HPC2_and_p_0_out_1__0_,
         cell_1908_a_HPC2_and_p_1_out_0__1_,
         cell_1908_a_HPC2_and_p_1_out_1__0_,
         cell_1908_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1908_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1908_a_HPC2_and_p_1_in_0__1_, cell_1908_a_HPC2_and_p_1_in_1__0_,
         cell_1908_a_HPC2_and_s_out_0__1_, cell_1908_a_HPC2_and_s_out_1__0_,
         cell_1908_a_HPC2_and_p_0_in_0__1_, cell_1908_a_HPC2_and_p_0_in_1__0_,
         cell_1908_a_HPC2_and_s_in_0__1_, cell_1908_a_HPC2_and_s_in_1__0_,
         cell_1908_a_HPC2_and_z_0__0_, cell_1908_a_HPC2_and_z_1__1_,
         cell_1909_a_HPC2_and_n9, cell_1909_a_HPC2_and_n8,
         cell_1909_a_HPC2_and_n7, cell_1909_a_HPC2_and_p_0_out_0__1_,
         cell_1909_a_HPC2_and_p_0_out_1__0_,
         cell_1909_a_HPC2_and_p_1_out_0__1_,
         cell_1909_a_HPC2_and_p_1_out_1__0_,
         cell_1909_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1909_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1909_a_HPC2_and_p_1_in_0__1_, cell_1909_a_HPC2_and_p_1_in_1__0_,
         cell_1909_a_HPC2_and_s_out_0__1_, cell_1909_a_HPC2_and_s_out_1__0_,
         cell_1909_a_HPC2_and_p_0_in_0__1_, cell_1909_a_HPC2_and_p_0_in_1__0_,
         cell_1909_a_HPC2_and_s_in_0__1_, cell_1909_a_HPC2_and_s_in_1__0_,
         cell_1909_a_HPC2_and_z_0__0_, cell_1909_a_HPC2_and_z_1__1_,
         cell_1910_a_HPC2_and_n9, cell_1910_a_HPC2_and_n8,
         cell_1910_a_HPC2_and_n7, cell_1910_a_HPC2_and_p_0_out_0__1_,
         cell_1910_a_HPC2_and_p_0_out_1__0_,
         cell_1910_a_HPC2_and_p_1_out_0__1_,
         cell_1910_a_HPC2_and_p_1_out_1__0_,
         cell_1910_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1910_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1910_a_HPC2_and_p_1_in_0__1_, cell_1910_a_HPC2_and_p_1_in_1__0_,
         cell_1910_a_HPC2_and_s_out_0__1_, cell_1910_a_HPC2_and_s_out_1__0_,
         cell_1910_a_HPC2_and_p_0_in_0__1_, cell_1910_a_HPC2_and_p_0_in_1__0_,
         cell_1910_a_HPC2_and_s_in_0__1_, cell_1910_a_HPC2_and_s_in_1__0_,
         cell_1910_a_HPC2_and_z_0__0_, cell_1910_a_HPC2_and_z_1__1_,
         cell_1911_a_HPC2_and_n9, cell_1911_a_HPC2_and_n8,
         cell_1911_a_HPC2_and_n7, cell_1911_a_HPC2_and_p_0_out_0__1_,
         cell_1911_a_HPC2_and_p_0_out_1__0_,
         cell_1911_a_HPC2_and_p_1_out_0__1_,
         cell_1911_a_HPC2_and_p_1_out_1__0_,
         cell_1911_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1911_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1911_a_HPC2_and_p_1_in_0__1_, cell_1911_a_HPC2_and_p_1_in_1__0_,
         cell_1911_a_HPC2_and_s_out_0__1_, cell_1911_a_HPC2_and_s_out_1__0_,
         cell_1911_a_HPC2_and_p_0_in_0__1_, cell_1911_a_HPC2_and_p_0_in_1__0_,
         cell_1911_a_HPC2_and_s_in_0__1_, cell_1911_a_HPC2_and_s_in_1__0_,
         cell_1911_a_HPC2_and_z_0__0_, cell_1911_a_HPC2_and_z_1__1_,
         cell_1912_a_HPC2_and_n9, cell_1912_a_HPC2_and_n8,
         cell_1912_a_HPC2_and_n7, cell_1912_a_HPC2_and_p_0_out_0__1_,
         cell_1912_a_HPC2_and_p_0_out_1__0_,
         cell_1912_a_HPC2_and_p_1_out_0__1_,
         cell_1912_a_HPC2_and_p_1_out_1__0_,
         cell_1912_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1912_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1912_a_HPC2_and_p_1_in_0__1_, cell_1912_a_HPC2_and_p_1_in_1__0_,
         cell_1912_a_HPC2_and_s_out_0__1_, cell_1912_a_HPC2_and_s_out_1__0_,
         cell_1912_a_HPC2_and_p_0_in_0__1_, cell_1912_a_HPC2_and_p_0_in_1__0_,
         cell_1912_a_HPC2_and_s_in_0__1_, cell_1912_a_HPC2_and_s_in_1__0_,
         cell_1912_a_HPC2_and_z_0__0_, cell_1912_a_HPC2_and_z_1__1_,
         cell_1913_a_HPC2_and_n9, cell_1913_a_HPC2_and_n8,
         cell_1913_a_HPC2_and_n7, cell_1913_a_HPC2_and_p_0_out_0__1_,
         cell_1913_a_HPC2_and_p_0_out_1__0_,
         cell_1913_a_HPC2_and_p_1_out_0__1_,
         cell_1913_a_HPC2_and_p_1_out_1__0_,
         cell_1913_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1913_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1913_a_HPC2_and_p_1_in_0__1_, cell_1913_a_HPC2_and_p_1_in_1__0_,
         cell_1913_a_HPC2_and_s_out_0__1_, cell_1913_a_HPC2_and_s_out_1__0_,
         cell_1913_a_HPC2_and_p_0_in_0__1_, cell_1913_a_HPC2_and_p_0_in_1__0_,
         cell_1913_a_HPC2_and_s_in_0__1_, cell_1913_a_HPC2_and_s_in_1__0_,
         cell_1913_a_HPC2_and_z_0__0_, cell_1913_a_HPC2_and_z_1__1_,
         cell_1914_a_HPC2_and_n9, cell_1914_a_HPC2_and_n8,
         cell_1914_a_HPC2_and_n7, cell_1914_a_HPC2_and_p_0_out_0__1_,
         cell_1914_a_HPC2_and_p_0_out_1__0_,
         cell_1914_a_HPC2_and_p_1_out_0__1_,
         cell_1914_a_HPC2_and_p_1_out_1__0_,
         cell_1914_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1914_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1914_a_HPC2_and_p_1_in_0__1_, cell_1914_a_HPC2_and_p_1_in_1__0_,
         cell_1914_a_HPC2_and_s_out_0__1_, cell_1914_a_HPC2_and_s_out_1__0_,
         cell_1914_a_HPC2_and_p_0_in_0__1_, cell_1914_a_HPC2_and_p_0_in_1__0_,
         cell_1914_a_HPC2_and_s_in_0__1_, cell_1914_a_HPC2_and_s_in_1__0_,
         cell_1914_a_HPC2_and_z_0__0_, cell_1914_a_HPC2_and_z_1__1_,
         cell_1915_a_HPC2_and_n9, cell_1915_a_HPC2_and_n8,
         cell_1915_a_HPC2_and_n7, cell_1915_a_HPC2_and_p_0_out_0__1_,
         cell_1915_a_HPC2_and_p_0_out_1__0_,
         cell_1915_a_HPC2_and_p_1_out_0__1_,
         cell_1915_a_HPC2_and_p_1_out_1__0_,
         cell_1915_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1915_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1915_a_HPC2_and_p_1_in_0__1_, cell_1915_a_HPC2_and_p_1_in_1__0_,
         cell_1915_a_HPC2_and_s_out_0__1_, cell_1915_a_HPC2_and_s_out_1__0_,
         cell_1915_a_HPC2_and_p_0_in_0__1_, cell_1915_a_HPC2_and_p_0_in_1__0_,
         cell_1915_a_HPC2_and_s_in_0__1_, cell_1915_a_HPC2_and_s_in_1__0_,
         cell_1915_a_HPC2_and_z_0__0_, cell_1915_a_HPC2_and_z_1__1_,
         cell_1916_a_HPC2_and_n9, cell_1916_a_HPC2_and_n8,
         cell_1916_a_HPC2_and_n7, cell_1916_a_HPC2_and_p_0_out_0__1_,
         cell_1916_a_HPC2_and_p_0_out_1__0_,
         cell_1916_a_HPC2_and_p_1_out_0__1_,
         cell_1916_a_HPC2_and_p_1_out_1__0_,
         cell_1916_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1916_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1916_a_HPC2_and_p_1_in_0__1_, cell_1916_a_HPC2_and_p_1_in_1__0_,
         cell_1916_a_HPC2_and_s_out_0__1_, cell_1916_a_HPC2_and_s_out_1__0_,
         cell_1916_a_HPC2_and_p_0_in_0__1_, cell_1916_a_HPC2_and_p_0_in_1__0_,
         cell_1916_a_HPC2_and_s_in_0__1_, cell_1916_a_HPC2_and_s_in_1__0_,
         cell_1916_a_HPC2_and_z_0__0_, cell_1916_a_HPC2_and_z_1__1_,
         cell_1917_a_HPC2_and_n9, cell_1917_a_HPC2_and_n8,
         cell_1917_a_HPC2_and_n7, cell_1917_a_HPC2_and_p_0_out_0__1_,
         cell_1917_a_HPC2_and_p_0_out_1__0_,
         cell_1917_a_HPC2_and_p_1_out_0__1_,
         cell_1917_a_HPC2_and_p_1_out_1__0_,
         cell_1917_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1917_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1917_a_HPC2_and_p_1_in_0__1_, cell_1917_a_HPC2_and_p_1_in_1__0_,
         cell_1917_a_HPC2_and_s_out_0__1_, cell_1917_a_HPC2_and_s_out_1__0_,
         cell_1917_a_HPC2_and_p_0_in_0__1_, cell_1917_a_HPC2_and_p_0_in_1__0_,
         cell_1917_a_HPC2_and_s_in_0__1_, cell_1917_a_HPC2_and_s_in_1__0_,
         cell_1917_a_HPC2_and_z_0__0_, cell_1917_a_HPC2_and_z_1__1_,
         cell_1918_a_HPC2_and_n9, cell_1918_a_HPC2_and_n8,
         cell_1918_a_HPC2_and_n7, cell_1918_a_HPC2_and_p_0_out_0__1_,
         cell_1918_a_HPC2_and_p_0_out_1__0_,
         cell_1918_a_HPC2_and_p_1_out_0__1_,
         cell_1918_a_HPC2_and_p_1_out_1__0_,
         cell_1918_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1918_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1918_a_HPC2_and_p_1_in_0__1_, cell_1918_a_HPC2_and_p_1_in_1__0_,
         cell_1918_a_HPC2_and_s_out_0__1_, cell_1918_a_HPC2_and_s_out_1__0_,
         cell_1918_a_HPC2_and_p_0_in_0__1_, cell_1918_a_HPC2_and_p_0_in_1__0_,
         cell_1918_a_HPC2_and_s_in_0__1_, cell_1918_a_HPC2_and_s_in_1__0_,
         cell_1918_a_HPC2_and_z_0__0_, cell_1918_a_HPC2_and_z_1__1_,
         cell_1919_a_HPC2_and_n9, cell_1919_a_HPC2_and_n8,
         cell_1919_a_HPC2_and_n7, cell_1919_a_HPC2_and_p_0_out_0__1_,
         cell_1919_a_HPC2_and_p_0_out_1__0_,
         cell_1919_a_HPC2_and_p_1_out_0__1_,
         cell_1919_a_HPC2_and_p_1_out_1__0_,
         cell_1919_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1919_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1919_a_HPC2_and_p_1_in_0__1_, cell_1919_a_HPC2_and_p_1_in_1__0_,
         cell_1919_a_HPC2_and_s_out_0__1_, cell_1919_a_HPC2_and_s_out_1__0_,
         cell_1919_a_HPC2_and_p_0_in_0__1_, cell_1919_a_HPC2_and_p_0_in_1__0_,
         cell_1919_a_HPC2_and_s_in_0__1_, cell_1919_a_HPC2_and_s_in_1__0_,
         cell_1919_a_HPC2_and_z_0__0_, cell_1919_a_HPC2_and_z_1__1_,
         cell_1920_a_HPC2_and_n9, cell_1920_a_HPC2_and_n8,
         cell_1920_a_HPC2_and_n7, cell_1920_a_HPC2_and_p_0_out_0__1_,
         cell_1920_a_HPC2_and_p_0_out_1__0_,
         cell_1920_a_HPC2_and_p_1_out_0__1_,
         cell_1920_a_HPC2_and_p_1_out_1__0_,
         cell_1920_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1920_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1920_a_HPC2_and_p_1_in_0__1_, cell_1920_a_HPC2_and_p_1_in_1__0_,
         cell_1920_a_HPC2_and_s_out_0__1_, cell_1920_a_HPC2_and_s_out_1__0_,
         cell_1920_a_HPC2_and_p_0_in_0__1_, cell_1920_a_HPC2_and_p_0_in_1__0_,
         cell_1920_a_HPC2_and_s_in_0__1_, cell_1920_a_HPC2_and_s_in_1__0_,
         cell_1920_a_HPC2_and_z_0__0_, cell_1920_a_HPC2_and_z_1__1_,
         cell_1921_a_HPC2_and_n9, cell_1921_a_HPC2_and_n8,
         cell_1921_a_HPC2_and_n7, cell_1921_a_HPC2_and_p_0_out_0__1_,
         cell_1921_a_HPC2_and_p_0_out_1__0_,
         cell_1921_a_HPC2_and_p_1_out_0__1_,
         cell_1921_a_HPC2_and_p_1_out_1__0_,
         cell_1921_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1921_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1921_a_HPC2_and_p_1_in_0__1_, cell_1921_a_HPC2_and_p_1_in_1__0_,
         cell_1921_a_HPC2_and_s_out_0__1_, cell_1921_a_HPC2_and_s_out_1__0_,
         cell_1921_a_HPC2_and_p_0_in_0__1_, cell_1921_a_HPC2_and_p_0_in_1__0_,
         cell_1921_a_HPC2_and_s_in_0__1_, cell_1921_a_HPC2_and_s_in_1__0_,
         cell_1921_a_HPC2_and_z_0__0_, cell_1921_a_HPC2_and_z_1__1_,
         cell_1922_a_HPC2_and_n9, cell_1922_a_HPC2_and_n8,
         cell_1922_a_HPC2_and_n7, cell_1922_a_HPC2_and_p_0_out_0__1_,
         cell_1922_a_HPC2_and_p_0_out_1__0_,
         cell_1922_a_HPC2_and_p_1_out_0__1_,
         cell_1922_a_HPC2_and_p_1_out_1__0_,
         cell_1922_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1922_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1922_a_HPC2_and_p_1_in_0__1_, cell_1922_a_HPC2_and_p_1_in_1__0_,
         cell_1922_a_HPC2_and_s_out_0__1_, cell_1922_a_HPC2_and_s_out_1__0_,
         cell_1922_a_HPC2_and_p_0_in_0__1_, cell_1922_a_HPC2_and_p_0_in_1__0_,
         cell_1922_a_HPC2_and_s_in_0__1_, cell_1922_a_HPC2_and_s_in_1__0_,
         cell_1922_a_HPC2_and_z_0__0_, cell_1922_a_HPC2_and_z_1__1_,
         cell_1923_a_HPC2_and_n9, cell_1923_a_HPC2_and_n8,
         cell_1923_a_HPC2_and_n7, cell_1923_a_HPC2_and_p_0_out_0__1_,
         cell_1923_a_HPC2_and_p_0_out_1__0_,
         cell_1923_a_HPC2_and_p_1_out_0__1_,
         cell_1923_a_HPC2_and_p_1_out_1__0_,
         cell_1923_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1923_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1923_a_HPC2_and_p_1_in_0__1_, cell_1923_a_HPC2_and_p_1_in_1__0_,
         cell_1923_a_HPC2_and_s_out_0__1_, cell_1923_a_HPC2_and_s_out_1__0_,
         cell_1923_a_HPC2_and_p_0_in_0__1_, cell_1923_a_HPC2_and_p_0_in_1__0_,
         cell_1923_a_HPC2_and_s_in_0__1_, cell_1923_a_HPC2_and_s_in_1__0_,
         cell_1923_a_HPC2_and_z_0__0_, cell_1923_a_HPC2_and_z_1__1_,
         cell_1924_a_HPC2_and_n9, cell_1924_a_HPC2_and_n8,
         cell_1924_a_HPC2_and_n7, cell_1924_a_HPC2_and_p_0_out_0__1_,
         cell_1924_a_HPC2_and_p_0_out_1__0_,
         cell_1924_a_HPC2_and_p_1_out_0__1_,
         cell_1924_a_HPC2_and_p_1_out_1__0_,
         cell_1924_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1924_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1924_a_HPC2_and_p_1_in_0__1_, cell_1924_a_HPC2_and_p_1_in_1__0_,
         cell_1924_a_HPC2_and_s_out_0__1_, cell_1924_a_HPC2_and_s_out_1__0_,
         cell_1924_a_HPC2_and_p_0_in_0__1_, cell_1924_a_HPC2_and_p_0_in_1__0_,
         cell_1924_a_HPC2_and_s_in_0__1_, cell_1924_a_HPC2_and_s_in_1__0_,
         cell_1924_a_HPC2_and_z_0__0_, cell_1924_a_HPC2_and_z_1__1_,
         cell_1925_a_HPC2_and_n9, cell_1925_a_HPC2_and_n8,
         cell_1925_a_HPC2_and_n7, cell_1925_a_HPC2_and_p_0_out_0__1_,
         cell_1925_a_HPC2_and_p_0_out_1__0_,
         cell_1925_a_HPC2_and_p_1_out_0__1_,
         cell_1925_a_HPC2_and_p_1_out_1__0_,
         cell_1925_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1925_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1925_a_HPC2_and_p_1_in_0__1_, cell_1925_a_HPC2_and_p_1_in_1__0_,
         cell_1925_a_HPC2_and_s_out_0__1_, cell_1925_a_HPC2_and_s_out_1__0_,
         cell_1925_a_HPC2_and_p_0_in_0__1_, cell_1925_a_HPC2_and_p_0_in_1__0_,
         cell_1925_a_HPC2_and_s_in_0__1_, cell_1925_a_HPC2_and_s_in_1__0_,
         cell_1925_a_HPC2_and_z_0__0_, cell_1925_a_HPC2_and_z_1__1_,
         cell_1926_a_HPC2_and_n9, cell_1926_a_HPC2_and_n8,
         cell_1926_a_HPC2_and_n7, cell_1926_a_HPC2_and_p_0_out_0__1_,
         cell_1926_a_HPC2_and_p_0_out_1__0_,
         cell_1926_a_HPC2_and_p_1_out_0__1_,
         cell_1926_a_HPC2_and_p_1_out_1__0_,
         cell_1926_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1926_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1926_a_HPC2_and_p_1_in_0__1_, cell_1926_a_HPC2_and_p_1_in_1__0_,
         cell_1926_a_HPC2_and_s_out_0__1_, cell_1926_a_HPC2_and_s_out_1__0_,
         cell_1926_a_HPC2_and_p_0_in_0__1_, cell_1926_a_HPC2_and_p_0_in_1__0_,
         cell_1926_a_HPC2_and_s_in_0__1_, cell_1926_a_HPC2_and_s_in_1__0_,
         cell_1926_a_HPC2_and_z_0__0_, cell_1926_a_HPC2_and_z_1__1_,
         cell_1927_a_HPC2_and_n9, cell_1927_a_HPC2_and_n8,
         cell_1927_a_HPC2_and_n7, cell_1927_a_HPC2_and_p_0_out_0__1_,
         cell_1927_a_HPC2_and_p_0_out_1__0_,
         cell_1927_a_HPC2_and_p_1_out_0__1_,
         cell_1927_a_HPC2_and_p_1_out_1__0_,
         cell_1927_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1927_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1927_a_HPC2_and_p_1_in_0__1_, cell_1927_a_HPC2_and_p_1_in_1__0_,
         cell_1927_a_HPC2_and_s_out_0__1_, cell_1927_a_HPC2_and_s_out_1__0_,
         cell_1927_a_HPC2_and_p_0_in_0__1_, cell_1927_a_HPC2_and_p_0_in_1__0_,
         cell_1927_a_HPC2_and_s_in_0__1_, cell_1927_a_HPC2_and_s_in_1__0_,
         cell_1927_a_HPC2_and_z_0__0_, cell_1927_a_HPC2_and_z_1__1_,
         cell_1928_a_HPC2_and_n9, cell_1928_a_HPC2_and_n8,
         cell_1928_a_HPC2_and_n7, cell_1928_a_HPC2_and_p_0_out_0__1_,
         cell_1928_a_HPC2_and_p_0_out_1__0_,
         cell_1928_a_HPC2_and_p_1_out_0__1_,
         cell_1928_a_HPC2_and_p_1_out_1__0_,
         cell_1928_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1928_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1928_a_HPC2_and_p_1_in_0__1_, cell_1928_a_HPC2_and_p_1_in_1__0_,
         cell_1928_a_HPC2_and_s_out_0__1_, cell_1928_a_HPC2_and_s_out_1__0_,
         cell_1928_a_HPC2_and_p_0_in_0__1_, cell_1928_a_HPC2_and_p_0_in_1__0_,
         cell_1928_a_HPC2_and_s_in_0__1_, cell_1928_a_HPC2_and_s_in_1__0_,
         cell_1928_a_HPC2_and_z_0__0_, cell_1928_a_HPC2_and_z_1__1_,
         cell_1929_a_HPC2_and_n9, cell_1929_a_HPC2_and_n8,
         cell_1929_a_HPC2_and_n7, cell_1929_a_HPC2_and_p_0_out_0__1_,
         cell_1929_a_HPC2_and_p_0_out_1__0_,
         cell_1929_a_HPC2_and_p_1_out_0__1_,
         cell_1929_a_HPC2_and_p_1_out_1__0_,
         cell_1929_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1929_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1929_a_HPC2_and_p_1_in_0__1_, cell_1929_a_HPC2_and_p_1_in_1__0_,
         cell_1929_a_HPC2_and_s_out_0__1_, cell_1929_a_HPC2_and_s_out_1__0_,
         cell_1929_a_HPC2_and_p_0_in_0__1_, cell_1929_a_HPC2_and_p_0_in_1__0_,
         cell_1929_a_HPC2_and_s_in_0__1_, cell_1929_a_HPC2_and_s_in_1__0_,
         cell_1929_a_HPC2_and_z_0__0_, cell_1929_a_HPC2_and_z_1__1_,
         cell_1930_a_HPC2_and_n9, cell_1930_a_HPC2_and_n8,
         cell_1930_a_HPC2_and_n7, cell_1930_a_HPC2_and_p_0_out_0__1_,
         cell_1930_a_HPC2_and_p_0_out_1__0_,
         cell_1930_a_HPC2_and_p_1_out_0__1_,
         cell_1930_a_HPC2_and_p_1_out_1__0_,
         cell_1930_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1930_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1930_a_HPC2_and_p_1_in_0__1_, cell_1930_a_HPC2_and_p_1_in_1__0_,
         cell_1930_a_HPC2_and_s_out_0__1_, cell_1930_a_HPC2_and_s_out_1__0_,
         cell_1930_a_HPC2_and_p_0_in_0__1_, cell_1930_a_HPC2_and_p_0_in_1__0_,
         cell_1930_a_HPC2_and_s_in_0__1_, cell_1930_a_HPC2_and_s_in_1__0_,
         cell_1930_a_HPC2_and_z_0__0_, cell_1930_a_HPC2_and_z_1__1_,
         cell_1931_a_HPC2_and_n9, cell_1931_a_HPC2_and_n8,
         cell_1931_a_HPC2_and_n7, cell_1931_a_HPC2_and_p_0_out_0__1_,
         cell_1931_a_HPC2_and_p_0_out_1__0_,
         cell_1931_a_HPC2_and_p_1_out_0__1_,
         cell_1931_a_HPC2_and_p_1_out_1__0_,
         cell_1931_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1931_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1931_a_HPC2_and_p_1_in_0__1_, cell_1931_a_HPC2_and_p_1_in_1__0_,
         cell_1931_a_HPC2_and_s_out_0__1_, cell_1931_a_HPC2_and_s_out_1__0_,
         cell_1931_a_HPC2_and_p_0_in_0__1_, cell_1931_a_HPC2_and_p_0_in_1__0_,
         cell_1931_a_HPC2_and_s_in_0__1_, cell_1931_a_HPC2_and_s_in_1__0_,
         cell_1931_a_HPC2_and_z_0__0_, cell_1931_a_HPC2_and_z_1__1_,
         cell_1932_a_HPC2_and_n9, cell_1932_a_HPC2_and_n8,
         cell_1932_a_HPC2_and_n7, cell_1932_a_HPC2_and_p_0_out_0__1_,
         cell_1932_a_HPC2_and_p_0_out_1__0_,
         cell_1932_a_HPC2_and_p_1_out_0__1_,
         cell_1932_a_HPC2_and_p_1_out_1__0_,
         cell_1932_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1932_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1932_a_HPC2_and_p_1_in_0__1_, cell_1932_a_HPC2_and_p_1_in_1__0_,
         cell_1932_a_HPC2_and_s_out_0__1_, cell_1932_a_HPC2_and_s_out_1__0_,
         cell_1932_a_HPC2_and_p_0_in_0__1_, cell_1932_a_HPC2_and_p_0_in_1__0_,
         cell_1932_a_HPC2_and_s_in_0__1_, cell_1932_a_HPC2_and_s_in_1__0_,
         cell_1932_a_HPC2_and_z_0__0_, cell_1932_a_HPC2_and_z_1__1_,
         cell_1933_a_HPC2_and_n9, cell_1933_a_HPC2_and_n8,
         cell_1933_a_HPC2_and_n7, cell_1933_a_HPC2_and_p_0_out_0__1_,
         cell_1933_a_HPC2_and_p_0_out_1__0_,
         cell_1933_a_HPC2_and_p_1_out_0__1_,
         cell_1933_a_HPC2_and_p_1_out_1__0_,
         cell_1933_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1933_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1933_a_HPC2_and_p_1_in_0__1_, cell_1933_a_HPC2_and_p_1_in_1__0_,
         cell_1933_a_HPC2_and_s_out_0__1_, cell_1933_a_HPC2_and_s_out_1__0_,
         cell_1933_a_HPC2_and_p_0_in_0__1_, cell_1933_a_HPC2_and_p_0_in_1__0_,
         cell_1933_a_HPC2_and_s_in_0__1_, cell_1933_a_HPC2_and_s_in_1__0_,
         cell_1933_a_HPC2_and_z_0__0_, cell_1933_a_HPC2_and_z_1__1_,
         cell_1934_a_HPC2_and_n9, cell_1934_a_HPC2_and_n8,
         cell_1934_a_HPC2_and_n7, cell_1934_a_HPC2_and_p_0_out_0__1_,
         cell_1934_a_HPC2_and_p_0_out_1__0_,
         cell_1934_a_HPC2_and_p_1_out_0__1_,
         cell_1934_a_HPC2_and_p_1_out_1__0_,
         cell_1934_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1934_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1934_a_HPC2_and_p_1_in_0__1_, cell_1934_a_HPC2_and_p_1_in_1__0_,
         cell_1934_a_HPC2_and_s_out_0__1_, cell_1934_a_HPC2_and_s_out_1__0_,
         cell_1934_a_HPC2_and_p_0_in_0__1_, cell_1934_a_HPC2_and_p_0_in_1__0_,
         cell_1934_a_HPC2_and_s_in_0__1_, cell_1934_a_HPC2_and_s_in_1__0_,
         cell_1934_a_HPC2_and_z_0__0_, cell_1934_a_HPC2_and_z_1__1_,
         cell_1935_a_HPC2_and_n9, cell_1935_a_HPC2_and_n8,
         cell_1935_a_HPC2_and_n7, cell_1935_a_HPC2_and_p_0_out_0__1_,
         cell_1935_a_HPC2_and_p_0_out_1__0_,
         cell_1935_a_HPC2_and_p_1_out_0__1_,
         cell_1935_a_HPC2_and_p_1_out_1__0_,
         cell_1935_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1935_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1935_a_HPC2_and_p_1_in_0__1_, cell_1935_a_HPC2_and_p_1_in_1__0_,
         cell_1935_a_HPC2_and_s_out_0__1_, cell_1935_a_HPC2_and_s_out_1__0_,
         cell_1935_a_HPC2_and_p_0_in_0__1_, cell_1935_a_HPC2_and_p_0_in_1__0_,
         cell_1935_a_HPC2_and_s_in_0__1_, cell_1935_a_HPC2_and_s_in_1__0_,
         cell_1935_a_HPC2_and_z_0__0_, cell_1935_a_HPC2_and_z_1__1_,
         cell_1936_a_HPC2_and_n9, cell_1936_a_HPC2_and_n8,
         cell_1936_a_HPC2_and_n7, cell_1936_a_HPC2_and_p_0_out_0__1_,
         cell_1936_a_HPC2_and_p_0_out_1__0_,
         cell_1936_a_HPC2_and_p_1_out_0__1_,
         cell_1936_a_HPC2_and_p_1_out_1__0_,
         cell_1936_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1936_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1936_a_HPC2_and_p_1_in_0__1_, cell_1936_a_HPC2_and_p_1_in_1__0_,
         cell_1936_a_HPC2_and_s_out_0__1_, cell_1936_a_HPC2_and_s_out_1__0_,
         cell_1936_a_HPC2_and_p_0_in_0__1_, cell_1936_a_HPC2_and_p_0_in_1__0_,
         cell_1936_a_HPC2_and_s_in_0__1_, cell_1936_a_HPC2_and_s_in_1__0_,
         cell_1936_a_HPC2_and_z_0__0_, cell_1936_a_HPC2_and_z_1__1_,
         cell_1937_a_HPC2_and_n9, cell_1937_a_HPC2_and_n8,
         cell_1937_a_HPC2_and_n7, cell_1937_a_HPC2_and_p_0_out_0__1_,
         cell_1937_a_HPC2_and_p_0_out_1__0_,
         cell_1937_a_HPC2_and_p_1_out_0__1_,
         cell_1937_a_HPC2_and_p_1_out_1__0_,
         cell_1937_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1937_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1937_a_HPC2_and_p_1_in_0__1_, cell_1937_a_HPC2_and_p_1_in_1__0_,
         cell_1937_a_HPC2_and_s_out_0__1_, cell_1937_a_HPC2_and_s_out_1__0_,
         cell_1937_a_HPC2_and_p_0_in_0__1_, cell_1937_a_HPC2_and_p_0_in_1__0_,
         cell_1937_a_HPC2_and_s_in_0__1_, cell_1937_a_HPC2_and_s_in_1__0_,
         cell_1937_a_HPC2_and_z_0__0_, cell_1937_a_HPC2_and_z_1__1_,
         cell_1938_a_HPC2_and_n9, cell_1938_a_HPC2_and_n8,
         cell_1938_a_HPC2_and_n7, cell_1938_a_HPC2_and_p_0_out_0__1_,
         cell_1938_a_HPC2_and_p_0_out_1__0_,
         cell_1938_a_HPC2_and_p_1_out_0__1_,
         cell_1938_a_HPC2_and_p_1_out_1__0_,
         cell_1938_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1938_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1938_a_HPC2_and_p_1_in_0__1_, cell_1938_a_HPC2_and_p_1_in_1__0_,
         cell_1938_a_HPC2_and_s_out_0__1_, cell_1938_a_HPC2_and_s_out_1__0_,
         cell_1938_a_HPC2_and_p_0_in_0__1_, cell_1938_a_HPC2_and_p_0_in_1__0_,
         cell_1938_a_HPC2_and_s_in_0__1_, cell_1938_a_HPC2_and_s_in_1__0_,
         cell_1938_a_HPC2_and_z_0__0_, cell_1938_a_HPC2_and_z_1__1_,
         cell_1939_a_HPC2_and_n9, cell_1939_a_HPC2_and_n8,
         cell_1939_a_HPC2_and_n7, cell_1939_a_HPC2_and_p_0_out_0__1_,
         cell_1939_a_HPC2_and_p_0_out_1__0_,
         cell_1939_a_HPC2_and_p_1_out_0__1_,
         cell_1939_a_HPC2_and_p_1_out_1__0_,
         cell_1939_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1939_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1939_a_HPC2_and_p_1_in_0__1_, cell_1939_a_HPC2_and_p_1_in_1__0_,
         cell_1939_a_HPC2_and_s_out_0__1_, cell_1939_a_HPC2_and_s_out_1__0_,
         cell_1939_a_HPC2_and_p_0_in_0__1_, cell_1939_a_HPC2_and_p_0_in_1__0_,
         cell_1939_a_HPC2_and_s_in_0__1_, cell_1939_a_HPC2_and_s_in_1__0_,
         cell_1939_a_HPC2_and_z_0__0_, cell_1939_a_HPC2_and_z_1__1_,
         cell_1940_a_HPC2_and_n9, cell_1940_a_HPC2_and_n8,
         cell_1940_a_HPC2_and_n7, cell_1940_a_HPC2_and_p_0_out_0__1_,
         cell_1940_a_HPC2_and_p_0_out_1__0_,
         cell_1940_a_HPC2_and_p_1_out_0__1_,
         cell_1940_a_HPC2_and_p_1_out_1__0_,
         cell_1940_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1940_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1940_a_HPC2_and_p_1_in_0__1_, cell_1940_a_HPC2_and_p_1_in_1__0_,
         cell_1940_a_HPC2_and_s_out_0__1_, cell_1940_a_HPC2_and_s_out_1__0_,
         cell_1940_a_HPC2_and_p_0_in_0__1_, cell_1940_a_HPC2_and_p_0_in_1__0_,
         cell_1940_a_HPC2_and_s_in_0__1_, cell_1940_a_HPC2_and_s_in_1__0_,
         cell_1940_a_HPC2_and_z_0__0_, cell_1940_a_HPC2_and_z_1__1_,
         cell_1941_a_HPC2_and_n9, cell_1941_a_HPC2_and_n8,
         cell_1941_a_HPC2_and_n7, cell_1941_a_HPC2_and_p_0_out_0__1_,
         cell_1941_a_HPC2_and_p_0_out_1__0_,
         cell_1941_a_HPC2_and_p_1_out_0__1_,
         cell_1941_a_HPC2_and_p_1_out_1__0_,
         cell_1941_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1941_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1941_a_HPC2_and_p_1_in_0__1_, cell_1941_a_HPC2_and_p_1_in_1__0_,
         cell_1941_a_HPC2_and_s_out_0__1_, cell_1941_a_HPC2_and_s_out_1__0_,
         cell_1941_a_HPC2_and_p_0_in_0__1_, cell_1941_a_HPC2_and_p_0_in_1__0_,
         cell_1941_a_HPC2_and_s_in_0__1_, cell_1941_a_HPC2_and_s_in_1__0_,
         cell_1941_a_HPC2_and_z_0__0_, cell_1941_a_HPC2_and_z_1__1_,
         cell_1942_a_HPC2_and_n9, cell_1942_a_HPC2_and_n8,
         cell_1942_a_HPC2_and_n7, cell_1942_a_HPC2_and_p_0_out_0__1_,
         cell_1942_a_HPC2_and_p_0_out_1__0_,
         cell_1942_a_HPC2_and_p_1_out_0__1_,
         cell_1942_a_HPC2_and_p_1_out_1__0_,
         cell_1942_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1942_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1942_a_HPC2_and_p_1_in_0__1_, cell_1942_a_HPC2_and_p_1_in_1__0_,
         cell_1942_a_HPC2_and_s_out_0__1_, cell_1942_a_HPC2_and_s_out_1__0_,
         cell_1942_a_HPC2_and_p_0_in_0__1_, cell_1942_a_HPC2_and_p_0_in_1__0_,
         cell_1942_a_HPC2_and_s_in_0__1_, cell_1942_a_HPC2_and_s_in_1__0_,
         cell_1942_a_HPC2_and_z_0__0_, cell_1942_a_HPC2_and_z_1__1_,
         cell_1943_a_HPC2_and_n9, cell_1943_a_HPC2_and_n8,
         cell_1943_a_HPC2_and_n7, cell_1943_a_HPC2_and_p_0_out_0__1_,
         cell_1943_a_HPC2_and_p_0_out_1__0_,
         cell_1943_a_HPC2_and_p_1_out_0__1_,
         cell_1943_a_HPC2_and_p_1_out_1__0_,
         cell_1943_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1943_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1943_a_HPC2_and_p_1_in_0__1_, cell_1943_a_HPC2_and_p_1_in_1__0_,
         cell_1943_a_HPC2_and_s_out_0__1_, cell_1943_a_HPC2_and_s_out_1__0_,
         cell_1943_a_HPC2_and_p_0_in_0__1_, cell_1943_a_HPC2_and_p_0_in_1__0_,
         cell_1943_a_HPC2_and_s_in_0__1_, cell_1943_a_HPC2_and_s_in_1__0_,
         cell_1943_a_HPC2_and_z_0__0_, cell_1943_a_HPC2_and_z_1__1_,
         cell_1944_a_HPC2_and_n9, cell_1944_a_HPC2_and_n8,
         cell_1944_a_HPC2_and_n7, cell_1944_a_HPC2_and_p_0_out_0__1_,
         cell_1944_a_HPC2_and_p_0_out_1__0_,
         cell_1944_a_HPC2_and_p_1_out_0__1_,
         cell_1944_a_HPC2_and_p_1_out_1__0_,
         cell_1944_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1944_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1944_a_HPC2_and_p_1_in_0__1_, cell_1944_a_HPC2_and_p_1_in_1__0_,
         cell_1944_a_HPC2_and_s_out_0__1_, cell_1944_a_HPC2_and_s_out_1__0_,
         cell_1944_a_HPC2_and_p_0_in_0__1_, cell_1944_a_HPC2_and_p_0_in_1__0_,
         cell_1944_a_HPC2_and_s_in_0__1_, cell_1944_a_HPC2_and_s_in_1__0_,
         cell_1944_a_HPC2_and_z_0__0_, cell_1944_a_HPC2_and_z_1__1_,
         cell_1945_a_HPC2_and_n9, cell_1945_a_HPC2_and_n8,
         cell_1945_a_HPC2_and_n7, cell_1945_a_HPC2_and_p_0_out_0__1_,
         cell_1945_a_HPC2_and_p_0_out_1__0_,
         cell_1945_a_HPC2_and_p_1_out_0__1_,
         cell_1945_a_HPC2_and_p_1_out_1__0_,
         cell_1945_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1945_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1945_a_HPC2_and_p_1_in_0__1_, cell_1945_a_HPC2_and_p_1_in_1__0_,
         cell_1945_a_HPC2_and_s_out_0__1_, cell_1945_a_HPC2_and_s_out_1__0_,
         cell_1945_a_HPC2_and_p_0_in_0__1_, cell_1945_a_HPC2_and_p_0_in_1__0_,
         cell_1945_a_HPC2_and_s_in_0__1_, cell_1945_a_HPC2_and_s_in_1__0_,
         cell_1945_a_HPC2_and_z_0__0_, cell_1945_a_HPC2_and_z_1__1_,
         cell_1946_a_HPC2_and_n9, cell_1946_a_HPC2_and_n8,
         cell_1946_a_HPC2_and_n7, cell_1946_a_HPC2_and_p_0_out_0__1_,
         cell_1946_a_HPC2_and_p_0_out_1__0_,
         cell_1946_a_HPC2_and_p_1_out_0__1_,
         cell_1946_a_HPC2_and_p_1_out_1__0_,
         cell_1946_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1946_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1946_a_HPC2_and_p_1_in_0__1_, cell_1946_a_HPC2_and_p_1_in_1__0_,
         cell_1946_a_HPC2_and_s_out_0__1_, cell_1946_a_HPC2_and_s_out_1__0_,
         cell_1946_a_HPC2_and_p_0_in_0__1_, cell_1946_a_HPC2_and_p_0_in_1__0_,
         cell_1946_a_HPC2_and_s_in_0__1_, cell_1946_a_HPC2_and_s_in_1__0_,
         cell_1946_a_HPC2_and_z_0__0_, cell_1946_a_HPC2_and_z_1__1_,
         cell_1947_a_HPC2_and_n9, cell_1947_a_HPC2_and_n8,
         cell_1947_a_HPC2_and_n7, cell_1947_a_HPC2_and_p_0_out_0__1_,
         cell_1947_a_HPC2_and_p_0_out_1__0_,
         cell_1947_a_HPC2_and_p_1_out_0__1_,
         cell_1947_a_HPC2_and_p_1_out_1__0_,
         cell_1947_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1947_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1947_a_HPC2_and_p_1_in_0__1_, cell_1947_a_HPC2_and_p_1_in_1__0_,
         cell_1947_a_HPC2_and_s_out_0__1_, cell_1947_a_HPC2_and_s_out_1__0_,
         cell_1947_a_HPC2_and_p_0_in_0__1_, cell_1947_a_HPC2_and_p_0_in_1__0_,
         cell_1947_a_HPC2_and_s_in_0__1_, cell_1947_a_HPC2_and_s_in_1__0_,
         cell_1947_a_HPC2_and_z_0__0_, cell_1947_a_HPC2_and_z_1__1_,
         cell_1948_a_HPC2_and_n9, cell_1948_a_HPC2_and_n8,
         cell_1948_a_HPC2_and_n7, cell_1948_a_HPC2_and_p_0_out_0__1_,
         cell_1948_a_HPC2_and_p_0_out_1__0_,
         cell_1948_a_HPC2_and_p_1_out_0__1_,
         cell_1948_a_HPC2_and_p_1_out_1__0_,
         cell_1948_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1948_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1948_a_HPC2_and_p_1_in_0__1_, cell_1948_a_HPC2_and_p_1_in_1__0_,
         cell_1948_a_HPC2_and_s_out_0__1_, cell_1948_a_HPC2_and_s_out_1__0_,
         cell_1948_a_HPC2_and_p_0_in_0__1_, cell_1948_a_HPC2_and_p_0_in_1__0_,
         cell_1948_a_HPC2_and_s_in_0__1_, cell_1948_a_HPC2_and_s_in_1__0_,
         cell_1948_a_HPC2_and_z_0__0_, cell_1948_a_HPC2_and_z_1__1_,
         cell_1949_a_HPC2_and_n9, cell_1949_a_HPC2_and_n8,
         cell_1949_a_HPC2_and_n7, cell_1949_a_HPC2_and_p_0_out_0__1_,
         cell_1949_a_HPC2_and_p_0_out_1__0_,
         cell_1949_a_HPC2_and_p_1_out_0__1_,
         cell_1949_a_HPC2_and_p_1_out_1__0_,
         cell_1949_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1949_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1949_a_HPC2_and_p_1_in_0__1_, cell_1949_a_HPC2_and_p_1_in_1__0_,
         cell_1949_a_HPC2_and_s_out_0__1_, cell_1949_a_HPC2_and_s_out_1__0_,
         cell_1949_a_HPC2_and_p_0_in_0__1_, cell_1949_a_HPC2_and_p_0_in_1__0_,
         cell_1949_a_HPC2_and_s_in_0__1_, cell_1949_a_HPC2_and_s_in_1__0_,
         cell_1949_a_HPC2_and_z_0__0_, cell_1949_a_HPC2_and_z_1__1_,
         cell_1950_a_HPC2_and_n9, cell_1950_a_HPC2_and_n8,
         cell_1950_a_HPC2_and_n7, cell_1950_a_HPC2_and_p_0_out_0__1_,
         cell_1950_a_HPC2_and_p_0_out_1__0_,
         cell_1950_a_HPC2_and_p_1_out_0__1_,
         cell_1950_a_HPC2_and_p_1_out_1__0_,
         cell_1950_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1950_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1950_a_HPC2_and_p_1_in_0__1_, cell_1950_a_HPC2_and_p_1_in_1__0_,
         cell_1950_a_HPC2_and_s_out_0__1_, cell_1950_a_HPC2_and_s_out_1__0_,
         cell_1950_a_HPC2_and_p_0_in_0__1_, cell_1950_a_HPC2_and_p_0_in_1__0_,
         cell_1950_a_HPC2_and_s_in_0__1_, cell_1950_a_HPC2_and_s_in_1__0_,
         cell_1950_a_HPC2_and_z_0__0_, cell_1950_a_HPC2_and_z_1__1_,
         cell_1951_a_HPC2_and_n9, cell_1951_a_HPC2_and_n8,
         cell_1951_a_HPC2_and_n7, cell_1951_a_HPC2_and_p_0_out_0__1_,
         cell_1951_a_HPC2_and_p_0_out_1__0_,
         cell_1951_a_HPC2_and_p_1_out_0__1_,
         cell_1951_a_HPC2_and_p_1_out_1__0_,
         cell_1951_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1951_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1951_a_HPC2_and_p_1_in_0__1_, cell_1951_a_HPC2_and_p_1_in_1__0_,
         cell_1951_a_HPC2_and_s_out_0__1_, cell_1951_a_HPC2_and_s_out_1__0_,
         cell_1951_a_HPC2_and_p_0_in_0__1_, cell_1951_a_HPC2_and_p_0_in_1__0_,
         cell_1951_a_HPC2_and_s_in_0__1_, cell_1951_a_HPC2_and_s_in_1__0_,
         cell_1951_a_HPC2_and_z_0__0_, cell_1951_a_HPC2_and_z_1__1_,
         cell_1952_a_HPC2_and_n9, cell_1952_a_HPC2_and_n8,
         cell_1952_a_HPC2_and_n7, cell_1952_a_HPC2_and_p_0_out_0__1_,
         cell_1952_a_HPC2_and_p_0_out_1__0_,
         cell_1952_a_HPC2_and_p_1_out_0__1_,
         cell_1952_a_HPC2_and_p_1_out_1__0_,
         cell_1952_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1952_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1952_a_HPC2_and_p_1_in_0__1_, cell_1952_a_HPC2_and_p_1_in_1__0_,
         cell_1952_a_HPC2_and_s_out_0__1_, cell_1952_a_HPC2_and_s_out_1__0_,
         cell_1952_a_HPC2_and_p_0_in_0__1_, cell_1952_a_HPC2_and_p_0_in_1__0_,
         cell_1952_a_HPC2_and_s_in_0__1_, cell_1952_a_HPC2_and_s_in_1__0_,
         cell_1952_a_HPC2_and_z_0__0_, cell_1952_a_HPC2_and_z_1__1_,
         cell_1953_a_HPC2_and_n9, cell_1953_a_HPC2_and_n8,
         cell_1953_a_HPC2_and_n7, cell_1953_a_HPC2_and_p_0_out_0__1_,
         cell_1953_a_HPC2_and_p_0_out_1__0_,
         cell_1953_a_HPC2_and_p_1_out_0__1_,
         cell_1953_a_HPC2_and_p_1_out_1__0_,
         cell_1953_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1953_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1953_a_HPC2_and_p_1_in_0__1_, cell_1953_a_HPC2_and_p_1_in_1__0_,
         cell_1953_a_HPC2_and_s_out_0__1_, cell_1953_a_HPC2_and_s_out_1__0_,
         cell_1953_a_HPC2_and_p_0_in_0__1_, cell_1953_a_HPC2_and_p_0_in_1__0_,
         cell_1953_a_HPC2_and_s_in_0__1_, cell_1953_a_HPC2_and_s_in_1__0_,
         cell_1953_a_HPC2_and_z_0__0_, cell_1953_a_HPC2_and_z_1__1_,
         cell_1954_a_HPC2_and_n9, cell_1954_a_HPC2_and_n8,
         cell_1954_a_HPC2_and_n7, cell_1954_a_HPC2_and_p_0_out_0__1_,
         cell_1954_a_HPC2_and_p_0_out_1__0_,
         cell_1954_a_HPC2_and_p_1_out_0__1_,
         cell_1954_a_HPC2_and_p_1_out_1__0_,
         cell_1954_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1954_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1954_a_HPC2_and_p_1_in_0__1_, cell_1954_a_HPC2_and_p_1_in_1__0_,
         cell_1954_a_HPC2_and_s_out_0__1_, cell_1954_a_HPC2_and_s_out_1__0_,
         cell_1954_a_HPC2_and_p_0_in_0__1_, cell_1954_a_HPC2_and_p_0_in_1__0_,
         cell_1954_a_HPC2_and_s_in_0__1_, cell_1954_a_HPC2_and_s_in_1__0_,
         cell_1954_a_HPC2_and_z_0__0_, cell_1954_a_HPC2_and_z_1__1_,
         cell_1955_a_HPC2_and_n9, cell_1955_a_HPC2_and_n8,
         cell_1955_a_HPC2_and_n7, cell_1955_a_HPC2_and_p_0_out_0__1_,
         cell_1955_a_HPC2_and_p_0_out_1__0_,
         cell_1955_a_HPC2_and_p_1_out_0__1_,
         cell_1955_a_HPC2_and_p_1_out_1__0_,
         cell_1955_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1955_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1955_a_HPC2_and_p_1_in_0__1_, cell_1955_a_HPC2_and_p_1_in_1__0_,
         cell_1955_a_HPC2_and_s_out_0__1_, cell_1955_a_HPC2_and_s_out_1__0_,
         cell_1955_a_HPC2_and_p_0_in_0__1_, cell_1955_a_HPC2_and_p_0_in_1__0_,
         cell_1955_a_HPC2_and_s_in_0__1_, cell_1955_a_HPC2_and_s_in_1__0_,
         cell_1955_a_HPC2_and_z_0__0_, cell_1955_a_HPC2_and_z_1__1_,
         cell_1956_a_HPC2_and_n9, cell_1956_a_HPC2_and_n8,
         cell_1956_a_HPC2_and_n7, cell_1956_a_HPC2_and_p_0_out_0__1_,
         cell_1956_a_HPC2_and_p_0_out_1__0_,
         cell_1956_a_HPC2_and_p_1_out_0__1_,
         cell_1956_a_HPC2_and_p_1_out_1__0_,
         cell_1956_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1956_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1956_a_HPC2_and_p_1_in_0__1_, cell_1956_a_HPC2_and_p_1_in_1__0_,
         cell_1956_a_HPC2_and_s_out_0__1_, cell_1956_a_HPC2_and_s_out_1__0_,
         cell_1956_a_HPC2_and_p_0_in_0__1_, cell_1956_a_HPC2_and_p_0_in_1__0_,
         cell_1956_a_HPC2_and_s_in_0__1_, cell_1956_a_HPC2_and_s_in_1__0_,
         cell_1956_a_HPC2_and_z_0__0_, cell_1956_a_HPC2_and_z_1__1_,
         cell_1957_a_HPC2_and_n9, cell_1957_a_HPC2_and_n8,
         cell_1957_a_HPC2_and_n7, cell_1957_a_HPC2_and_p_0_out_0__1_,
         cell_1957_a_HPC2_and_p_0_out_1__0_,
         cell_1957_a_HPC2_and_p_1_out_0__1_,
         cell_1957_a_HPC2_and_p_1_out_1__0_,
         cell_1957_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1957_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1957_a_HPC2_and_p_1_in_0__1_, cell_1957_a_HPC2_and_p_1_in_1__0_,
         cell_1957_a_HPC2_and_s_out_0__1_, cell_1957_a_HPC2_and_s_out_1__0_,
         cell_1957_a_HPC2_and_p_0_in_0__1_, cell_1957_a_HPC2_and_p_0_in_1__0_,
         cell_1957_a_HPC2_and_s_in_0__1_, cell_1957_a_HPC2_and_s_in_1__0_,
         cell_1957_a_HPC2_and_z_0__0_, cell_1957_a_HPC2_and_z_1__1_,
         cell_1958_a_HPC2_and_n9, cell_1958_a_HPC2_and_n8,
         cell_1958_a_HPC2_and_n7, cell_1958_a_HPC2_and_p_0_out_0__1_,
         cell_1958_a_HPC2_and_p_0_out_1__0_,
         cell_1958_a_HPC2_and_p_1_out_0__1_,
         cell_1958_a_HPC2_and_p_1_out_1__0_,
         cell_1958_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1958_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1958_a_HPC2_and_p_1_in_0__1_, cell_1958_a_HPC2_and_p_1_in_1__0_,
         cell_1958_a_HPC2_and_s_out_0__1_, cell_1958_a_HPC2_and_s_out_1__0_,
         cell_1958_a_HPC2_and_p_0_in_0__1_, cell_1958_a_HPC2_and_p_0_in_1__0_,
         cell_1958_a_HPC2_and_s_in_0__1_, cell_1958_a_HPC2_and_s_in_1__0_,
         cell_1958_a_HPC2_and_z_0__0_, cell_1958_a_HPC2_and_z_1__1_,
         cell_1959_a_HPC2_and_n9, cell_1959_a_HPC2_and_n8,
         cell_1959_a_HPC2_and_n7, cell_1959_a_HPC2_and_p_0_out_0__1_,
         cell_1959_a_HPC2_and_p_0_out_1__0_,
         cell_1959_a_HPC2_and_p_1_out_0__1_,
         cell_1959_a_HPC2_and_p_1_out_1__0_,
         cell_1959_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1959_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1959_a_HPC2_and_p_1_in_0__1_, cell_1959_a_HPC2_and_p_1_in_1__0_,
         cell_1959_a_HPC2_and_s_out_0__1_, cell_1959_a_HPC2_and_s_out_1__0_,
         cell_1959_a_HPC2_and_p_0_in_0__1_, cell_1959_a_HPC2_and_p_0_in_1__0_,
         cell_1959_a_HPC2_and_s_in_0__1_, cell_1959_a_HPC2_and_s_in_1__0_,
         cell_1959_a_HPC2_and_z_0__0_, cell_1959_a_HPC2_and_z_1__1_,
         cell_1960_a_HPC2_and_n9, cell_1960_a_HPC2_and_n8,
         cell_1960_a_HPC2_and_n7, cell_1960_a_HPC2_and_p_0_out_0__1_,
         cell_1960_a_HPC2_and_p_0_out_1__0_,
         cell_1960_a_HPC2_and_p_1_out_0__1_,
         cell_1960_a_HPC2_and_p_1_out_1__0_,
         cell_1960_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1960_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1960_a_HPC2_and_p_1_in_0__1_, cell_1960_a_HPC2_and_p_1_in_1__0_,
         cell_1960_a_HPC2_and_s_out_0__1_, cell_1960_a_HPC2_and_s_out_1__0_,
         cell_1960_a_HPC2_and_p_0_in_0__1_, cell_1960_a_HPC2_and_p_0_in_1__0_,
         cell_1960_a_HPC2_and_s_in_0__1_, cell_1960_a_HPC2_and_s_in_1__0_,
         cell_1960_a_HPC2_and_z_0__0_, cell_1960_a_HPC2_and_z_1__1_,
         cell_1961_a_HPC2_and_n9, cell_1961_a_HPC2_and_n8,
         cell_1961_a_HPC2_and_n7, cell_1961_a_HPC2_and_p_0_out_0__1_,
         cell_1961_a_HPC2_and_p_0_out_1__0_,
         cell_1961_a_HPC2_and_p_1_out_0__1_,
         cell_1961_a_HPC2_and_p_1_out_1__0_,
         cell_1961_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1961_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1961_a_HPC2_and_p_1_in_0__1_, cell_1961_a_HPC2_and_p_1_in_1__0_,
         cell_1961_a_HPC2_and_s_out_0__1_, cell_1961_a_HPC2_and_s_out_1__0_,
         cell_1961_a_HPC2_and_p_0_in_0__1_, cell_1961_a_HPC2_and_p_0_in_1__0_,
         cell_1961_a_HPC2_and_s_in_0__1_, cell_1961_a_HPC2_and_s_in_1__0_,
         cell_1961_a_HPC2_and_z_0__0_, cell_1961_a_HPC2_and_z_1__1_,
         cell_1962_a_HPC2_and_n9, cell_1962_a_HPC2_and_n8,
         cell_1962_a_HPC2_and_n7, cell_1962_a_HPC2_and_p_0_out_0__1_,
         cell_1962_a_HPC2_and_p_0_out_1__0_,
         cell_1962_a_HPC2_and_p_1_out_0__1_,
         cell_1962_a_HPC2_and_p_1_out_1__0_,
         cell_1962_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1962_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1962_a_HPC2_and_p_1_in_0__1_, cell_1962_a_HPC2_and_p_1_in_1__0_,
         cell_1962_a_HPC2_and_s_out_0__1_, cell_1962_a_HPC2_and_s_out_1__0_,
         cell_1962_a_HPC2_and_p_0_in_0__1_, cell_1962_a_HPC2_and_p_0_in_1__0_,
         cell_1962_a_HPC2_and_s_in_0__1_, cell_1962_a_HPC2_and_s_in_1__0_,
         cell_1962_a_HPC2_and_z_0__0_, cell_1962_a_HPC2_and_z_1__1_,
         cell_1963_a_HPC2_and_n9, cell_1963_a_HPC2_and_n8,
         cell_1963_a_HPC2_and_n7, cell_1963_a_HPC2_and_p_0_out_0__1_,
         cell_1963_a_HPC2_and_p_0_out_1__0_,
         cell_1963_a_HPC2_and_p_1_out_0__1_,
         cell_1963_a_HPC2_and_p_1_out_1__0_,
         cell_1963_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1963_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1963_a_HPC2_and_p_1_in_0__1_, cell_1963_a_HPC2_and_p_1_in_1__0_,
         cell_1963_a_HPC2_and_s_out_0__1_, cell_1963_a_HPC2_and_s_out_1__0_,
         cell_1963_a_HPC2_and_p_0_in_0__1_, cell_1963_a_HPC2_and_p_0_in_1__0_,
         cell_1963_a_HPC2_and_s_in_0__1_, cell_1963_a_HPC2_and_s_in_1__0_,
         cell_1963_a_HPC2_and_z_0__0_, cell_1963_a_HPC2_and_z_1__1_,
         cell_1964_a_HPC2_and_n9, cell_1964_a_HPC2_and_n8,
         cell_1964_a_HPC2_and_n7, cell_1964_a_HPC2_and_p_0_out_0__1_,
         cell_1964_a_HPC2_and_p_0_out_1__0_,
         cell_1964_a_HPC2_and_p_1_out_0__1_,
         cell_1964_a_HPC2_and_p_1_out_1__0_,
         cell_1964_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1964_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1964_a_HPC2_and_p_1_in_0__1_, cell_1964_a_HPC2_and_p_1_in_1__0_,
         cell_1964_a_HPC2_and_s_out_0__1_, cell_1964_a_HPC2_and_s_out_1__0_,
         cell_1964_a_HPC2_and_p_0_in_0__1_, cell_1964_a_HPC2_and_p_0_in_1__0_,
         cell_1964_a_HPC2_and_s_in_0__1_, cell_1964_a_HPC2_and_s_in_1__0_,
         cell_1964_a_HPC2_and_z_0__0_, cell_1964_a_HPC2_and_z_1__1_,
         cell_1965_a_HPC2_and_n9, cell_1965_a_HPC2_and_n8,
         cell_1965_a_HPC2_and_n7, cell_1965_a_HPC2_and_p_0_out_0__1_,
         cell_1965_a_HPC2_and_p_0_out_1__0_,
         cell_1965_a_HPC2_and_p_1_out_0__1_,
         cell_1965_a_HPC2_and_p_1_out_1__0_,
         cell_1965_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1965_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1965_a_HPC2_and_p_1_in_0__1_, cell_1965_a_HPC2_and_p_1_in_1__0_,
         cell_1965_a_HPC2_and_s_out_0__1_, cell_1965_a_HPC2_and_s_out_1__0_,
         cell_1965_a_HPC2_and_p_0_in_0__1_, cell_1965_a_HPC2_and_p_0_in_1__0_,
         cell_1965_a_HPC2_and_s_in_0__1_, cell_1965_a_HPC2_and_s_in_1__0_,
         cell_1965_a_HPC2_and_z_0__0_, cell_1965_a_HPC2_and_z_1__1_,
         cell_1966_a_HPC2_and_n9, cell_1966_a_HPC2_and_n8,
         cell_1966_a_HPC2_and_n7, cell_1966_a_HPC2_and_p_0_out_0__1_,
         cell_1966_a_HPC2_and_p_0_out_1__0_,
         cell_1966_a_HPC2_and_p_1_out_0__1_,
         cell_1966_a_HPC2_and_p_1_out_1__0_,
         cell_1966_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1966_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1966_a_HPC2_and_p_1_in_0__1_, cell_1966_a_HPC2_and_p_1_in_1__0_,
         cell_1966_a_HPC2_and_s_out_0__1_, cell_1966_a_HPC2_and_s_out_1__0_,
         cell_1966_a_HPC2_and_p_0_in_0__1_, cell_1966_a_HPC2_and_p_0_in_1__0_,
         cell_1966_a_HPC2_and_s_in_0__1_, cell_1966_a_HPC2_and_s_in_1__0_,
         cell_1966_a_HPC2_and_z_0__0_, cell_1966_a_HPC2_and_z_1__1_,
         cell_1967_a_HPC2_and_n9, cell_1967_a_HPC2_and_n8,
         cell_1967_a_HPC2_and_n7, cell_1967_a_HPC2_and_p_0_out_0__1_,
         cell_1967_a_HPC2_and_p_0_out_1__0_,
         cell_1967_a_HPC2_and_p_1_out_0__1_,
         cell_1967_a_HPC2_and_p_1_out_1__0_,
         cell_1967_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1967_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1967_a_HPC2_and_p_1_in_0__1_, cell_1967_a_HPC2_and_p_1_in_1__0_,
         cell_1967_a_HPC2_and_s_out_0__1_, cell_1967_a_HPC2_and_s_out_1__0_,
         cell_1967_a_HPC2_and_p_0_in_0__1_, cell_1967_a_HPC2_and_p_0_in_1__0_,
         cell_1967_a_HPC2_and_s_in_0__1_, cell_1967_a_HPC2_and_s_in_1__0_,
         cell_1967_a_HPC2_and_z_0__0_, cell_1967_a_HPC2_and_z_1__1_,
         cell_1968_a_HPC2_and_n9, cell_1968_a_HPC2_and_n8,
         cell_1968_a_HPC2_and_n7, cell_1968_a_HPC2_and_p_0_out_0__1_,
         cell_1968_a_HPC2_and_p_0_out_1__0_,
         cell_1968_a_HPC2_and_p_1_out_0__1_,
         cell_1968_a_HPC2_and_p_1_out_1__0_,
         cell_1968_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1968_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1968_a_HPC2_and_p_1_in_0__1_, cell_1968_a_HPC2_and_p_1_in_1__0_,
         cell_1968_a_HPC2_and_s_out_0__1_, cell_1968_a_HPC2_and_s_out_1__0_,
         cell_1968_a_HPC2_and_p_0_in_0__1_, cell_1968_a_HPC2_and_p_0_in_1__0_,
         cell_1968_a_HPC2_and_s_in_0__1_, cell_1968_a_HPC2_and_s_in_1__0_,
         cell_1968_a_HPC2_and_z_0__0_, cell_1968_a_HPC2_and_z_1__1_,
         cell_1969_a_HPC2_and_n9, cell_1969_a_HPC2_and_n8,
         cell_1969_a_HPC2_and_n7, cell_1969_a_HPC2_and_p_0_out_0__1_,
         cell_1969_a_HPC2_and_p_0_out_1__0_,
         cell_1969_a_HPC2_and_p_1_out_0__1_,
         cell_1969_a_HPC2_and_p_1_out_1__0_,
         cell_1969_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1969_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1969_a_HPC2_and_p_1_in_0__1_, cell_1969_a_HPC2_and_p_1_in_1__0_,
         cell_1969_a_HPC2_and_s_out_0__1_, cell_1969_a_HPC2_and_s_out_1__0_,
         cell_1969_a_HPC2_and_p_0_in_0__1_, cell_1969_a_HPC2_and_p_0_in_1__0_,
         cell_1969_a_HPC2_and_s_in_0__1_, cell_1969_a_HPC2_and_s_in_1__0_,
         cell_1969_a_HPC2_and_z_0__0_, cell_1969_a_HPC2_and_z_1__1_,
         cell_1970_a_HPC2_and_n9, cell_1970_a_HPC2_and_n8,
         cell_1970_a_HPC2_and_n7, cell_1970_a_HPC2_and_p_0_out_0__1_,
         cell_1970_a_HPC2_and_p_0_out_1__0_,
         cell_1970_a_HPC2_and_p_1_out_0__1_,
         cell_1970_a_HPC2_and_p_1_out_1__0_,
         cell_1970_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1970_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1970_a_HPC2_and_p_1_in_0__1_, cell_1970_a_HPC2_and_p_1_in_1__0_,
         cell_1970_a_HPC2_and_s_out_0__1_, cell_1970_a_HPC2_and_s_out_1__0_,
         cell_1970_a_HPC2_and_p_0_in_0__1_, cell_1970_a_HPC2_and_p_0_in_1__0_,
         cell_1970_a_HPC2_and_s_in_0__1_, cell_1970_a_HPC2_and_s_in_1__0_,
         cell_1970_a_HPC2_and_z_0__0_, cell_1970_a_HPC2_and_z_1__1_,
         cell_1971_a_HPC2_and_n9, cell_1971_a_HPC2_and_n8,
         cell_1971_a_HPC2_and_n7, cell_1971_a_HPC2_and_p_0_out_0__1_,
         cell_1971_a_HPC2_and_p_0_out_1__0_,
         cell_1971_a_HPC2_and_p_1_out_0__1_,
         cell_1971_a_HPC2_and_p_1_out_1__0_,
         cell_1971_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1971_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1971_a_HPC2_and_p_1_in_0__1_, cell_1971_a_HPC2_and_p_1_in_1__0_,
         cell_1971_a_HPC2_and_s_out_0__1_, cell_1971_a_HPC2_and_s_out_1__0_,
         cell_1971_a_HPC2_and_p_0_in_0__1_, cell_1971_a_HPC2_and_p_0_in_1__0_,
         cell_1971_a_HPC2_and_s_in_0__1_, cell_1971_a_HPC2_and_s_in_1__0_,
         cell_1971_a_HPC2_and_z_0__0_, cell_1971_a_HPC2_and_z_1__1_,
         cell_1972_a_HPC2_and_n9, cell_1972_a_HPC2_and_n8,
         cell_1972_a_HPC2_and_n7, cell_1972_a_HPC2_and_p_0_out_0__1_,
         cell_1972_a_HPC2_and_p_0_out_1__0_,
         cell_1972_a_HPC2_and_p_1_out_0__1_,
         cell_1972_a_HPC2_and_p_1_out_1__0_,
         cell_1972_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1972_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1972_a_HPC2_and_p_1_in_0__1_, cell_1972_a_HPC2_and_p_1_in_1__0_,
         cell_1972_a_HPC2_and_s_out_0__1_, cell_1972_a_HPC2_and_s_out_1__0_,
         cell_1972_a_HPC2_and_p_0_in_0__1_, cell_1972_a_HPC2_and_p_0_in_1__0_,
         cell_1972_a_HPC2_and_s_in_0__1_, cell_1972_a_HPC2_and_s_in_1__0_,
         cell_1972_a_HPC2_and_z_0__0_, cell_1972_a_HPC2_and_z_1__1_,
         cell_1973_a_HPC2_and_n9, cell_1973_a_HPC2_and_n8,
         cell_1973_a_HPC2_and_n7, cell_1973_a_HPC2_and_p_0_out_0__1_,
         cell_1973_a_HPC2_and_p_0_out_1__0_,
         cell_1973_a_HPC2_and_p_1_out_0__1_,
         cell_1973_a_HPC2_and_p_1_out_1__0_,
         cell_1973_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1973_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1973_a_HPC2_and_p_1_in_0__1_, cell_1973_a_HPC2_and_p_1_in_1__0_,
         cell_1973_a_HPC2_and_s_out_0__1_, cell_1973_a_HPC2_and_s_out_1__0_,
         cell_1973_a_HPC2_and_p_0_in_0__1_, cell_1973_a_HPC2_and_p_0_in_1__0_,
         cell_1973_a_HPC2_and_s_in_0__1_, cell_1973_a_HPC2_and_s_in_1__0_,
         cell_1973_a_HPC2_and_z_0__0_, cell_1973_a_HPC2_and_z_1__1_,
         cell_1974_a_HPC2_and_n9, cell_1974_a_HPC2_and_n8,
         cell_1974_a_HPC2_and_n7, cell_1974_a_HPC2_and_p_0_out_0__1_,
         cell_1974_a_HPC2_and_p_0_out_1__0_,
         cell_1974_a_HPC2_and_p_1_out_0__1_,
         cell_1974_a_HPC2_and_p_1_out_1__0_,
         cell_1974_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1974_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1974_a_HPC2_and_p_1_in_0__1_, cell_1974_a_HPC2_and_p_1_in_1__0_,
         cell_1974_a_HPC2_and_s_out_0__1_, cell_1974_a_HPC2_and_s_out_1__0_,
         cell_1974_a_HPC2_and_p_0_in_0__1_, cell_1974_a_HPC2_and_p_0_in_1__0_,
         cell_1974_a_HPC2_and_s_in_0__1_, cell_1974_a_HPC2_and_s_in_1__0_,
         cell_1974_a_HPC2_and_z_0__0_, cell_1974_a_HPC2_and_z_1__1_,
         cell_1975_a_HPC2_and_n9, cell_1975_a_HPC2_and_n8,
         cell_1975_a_HPC2_and_n7, cell_1975_a_HPC2_and_p_0_out_0__1_,
         cell_1975_a_HPC2_and_p_0_out_1__0_,
         cell_1975_a_HPC2_and_p_1_out_0__1_,
         cell_1975_a_HPC2_and_p_1_out_1__0_,
         cell_1975_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1975_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1975_a_HPC2_and_p_1_in_0__1_, cell_1975_a_HPC2_and_p_1_in_1__0_,
         cell_1975_a_HPC2_and_s_out_0__1_, cell_1975_a_HPC2_and_s_out_1__0_,
         cell_1975_a_HPC2_and_p_0_in_0__1_, cell_1975_a_HPC2_and_p_0_in_1__0_,
         cell_1975_a_HPC2_and_s_in_0__1_, cell_1975_a_HPC2_and_s_in_1__0_,
         cell_1975_a_HPC2_and_z_0__0_, cell_1975_a_HPC2_and_z_1__1_,
         cell_1976_a_HPC2_and_n9, cell_1976_a_HPC2_and_n8,
         cell_1976_a_HPC2_and_n7, cell_1976_a_HPC2_and_p_0_out_0__1_,
         cell_1976_a_HPC2_and_p_0_out_1__0_,
         cell_1976_a_HPC2_and_p_1_out_0__1_,
         cell_1976_a_HPC2_and_p_1_out_1__0_,
         cell_1976_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1976_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1976_a_HPC2_and_p_1_in_0__1_, cell_1976_a_HPC2_and_p_1_in_1__0_,
         cell_1976_a_HPC2_and_s_out_0__1_, cell_1976_a_HPC2_and_s_out_1__0_,
         cell_1976_a_HPC2_and_p_0_in_0__1_, cell_1976_a_HPC2_and_p_0_in_1__0_,
         cell_1976_a_HPC2_and_s_in_0__1_, cell_1976_a_HPC2_and_s_in_1__0_,
         cell_1976_a_HPC2_and_z_0__0_, cell_1976_a_HPC2_and_z_1__1_,
         cell_1977_a_HPC2_and_n9, cell_1977_a_HPC2_and_n8,
         cell_1977_a_HPC2_and_n7, cell_1977_a_HPC2_and_p_0_out_0__1_,
         cell_1977_a_HPC2_and_p_0_out_1__0_,
         cell_1977_a_HPC2_and_p_1_out_0__1_,
         cell_1977_a_HPC2_and_p_1_out_1__0_,
         cell_1977_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1977_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1977_a_HPC2_and_p_1_in_0__1_, cell_1977_a_HPC2_and_p_1_in_1__0_,
         cell_1977_a_HPC2_and_s_out_0__1_, cell_1977_a_HPC2_and_s_out_1__0_,
         cell_1977_a_HPC2_and_p_0_in_0__1_, cell_1977_a_HPC2_and_p_0_in_1__0_,
         cell_1977_a_HPC2_and_s_in_0__1_, cell_1977_a_HPC2_and_s_in_1__0_,
         cell_1977_a_HPC2_and_z_0__0_, cell_1977_a_HPC2_and_z_1__1_,
         cell_1978_a_HPC2_and_n9, cell_1978_a_HPC2_and_n8,
         cell_1978_a_HPC2_and_n7, cell_1978_a_HPC2_and_p_0_out_0__1_,
         cell_1978_a_HPC2_and_p_0_out_1__0_,
         cell_1978_a_HPC2_and_p_1_out_0__1_,
         cell_1978_a_HPC2_and_p_1_out_1__0_,
         cell_1978_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1978_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1978_a_HPC2_and_p_1_in_0__1_, cell_1978_a_HPC2_and_p_1_in_1__0_,
         cell_1978_a_HPC2_and_s_out_0__1_, cell_1978_a_HPC2_and_s_out_1__0_,
         cell_1978_a_HPC2_and_p_0_in_0__1_, cell_1978_a_HPC2_and_p_0_in_1__0_,
         cell_1978_a_HPC2_and_s_in_0__1_, cell_1978_a_HPC2_and_s_in_1__0_,
         cell_1978_a_HPC2_and_z_0__0_, cell_1978_a_HPC2_and_z_1__1_,
         cell_1979_a_HPC2_and_n9, cell_1979_a_HPC2_and_n8,
         cell_1979_a_HPC2_and_n7, cell_1979_a_HPC2_and_p_0_out_0__1_,
         cell_1979_a_HPC2_and_p_0_out_1__0_,
         cell_1979_a_HPC2_and_p_1_out_0__1_,
         cell_1979_a_HPC2_and_p_1_out_1__0_,
         cell_1979_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1979_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1979_a_HPC2_and_p_1_in_0__1_, cell_1979_a_HPC2_and_p_1_in_1__0_,
         cell_1979_a_HPC2_and_s_out_0__1_, cell_1979_a_HPC2_and_s_out_1__0_,
         cell_1979_a_HPC2_and_p_0_in_0__1_, cell_1979_a_HPC2_and_p_0_in_1__0_,
         cell_1979_a_HPC2_and_s_in_0__1_, cell_1979_a_HPC2_and_s_in_1__0_,
         cell_1979_a_HPC2_and_z_0__0_, cell_1979_a_HPC2_and_z_1__1_,
         cell_1980_a_HPC2_and_n9, cell_1980_a_HPC2_and_n8,
         cell_1980_a_HPC2_and_n7, cell_1980_a_HPC2_and_p_0_out_0__1_,
         cell_1980_a_HPC2_and_p_0_out_1__0_,
         cell_1980_a_HPC2_and_p_1_out_0__1_,
         cell_1980_a_HPC2_and_p_1_out_1__0_,
         cell_1980_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1980_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1980_a_HPC2_and_p_1_in_0__1_, cell_1980_a_HPC2_and_p_1_in_1__0_,
         cell_1980_a_HPC2_and_s_out_0__1_, cell_1980_a_HPC2_and_s_out_1__0_,
         cell_1980_a_HPC2_and_p_0_in_0__1_, cell_1980_a_HPC2_and_p_0_in_1__0_,
         cell_1980_a_HPC2_and_s_in_0__1_, cell_1980_a_HPC2_and_s_in_1__0_,
         cell_1980_a_HPC2_and_z_0__0_, cell_1980_a_HPC2_and_z_1__1_,
         cell_1981_a_HPC2_and_n9, cell_1981_a_HPC2_and_n8,
         cell_1981_a_HPC2_and_n7, cell_1981_a_HPC2_and_p_0_out_0__1_,
         cell_1981_a_HPC2_and_p_0_out_1__0_,
         cell_1981_a_HPC2_and_p_1_out_0__1_,
         cell_1981_a_HPC2_and_p_1_out_1__0_,
         cell_1981_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1981_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1981_a_HPC2_and_p_1_in_0__1_, cell_1981_a_HPC2_and_p_1_in_1__0_,
         cell_1981_a_HPC2_and_s_out_0__1_, cell_1981_a_HPC2_and_s_out_1__0_,
         cell_1981_a_HPC2_and_p_0_in_0__1_, cell_1981_a_HPC2_and_p_0_in_1__0_,
         cell_1981_a_HPC2_and_s_in_0__1_, cell_1981_a_HPC2_and_s_in_1__0_,
         cell_1981_a_HPC2_and_z_0__0_, cell_1981_a_HPC2_and_z_1__1_,
         cell_1982_a_HPC2_and_n9, cell_1982_a_HPC2_and_n8,
         cell_1982_a_HPC2_and_n7, cell_1982_a_HPC2_and_p_0_out_0__1_,
         cell_1982_a_HPC2_and_p_0_out_1__0_,
         cell_1982_a_HPC2_and_p_1_out_0__1_,
         cell_1982_a_HPC2_and_p_1_out_1__0_,
         cell_1982_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1982_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1982_a_HPC2_and_p_1_in_0__1_, cell_1982_a_HPC2_and_p_1_in_1__0_,
         cell_1982_a_HPC2_and_s_out_0__1_, cell_1982_a_HPC2_and_s_out_1__0_,
         cell_1982_a_HPC2_and_p_0_in_0__1_, cell_1982_a_HPC2_and_p_0_in_1__0_,
         cell_1982_a_HPC2_and_s_in_0__1_, cell_1982_a_HPC2_and_s_in_1__0_,
         cell_1982_a_HPC2_and_z_0__0_, cell_1982_a_HPC2_and_z_1__1_,
         cell_1983_a_HPC2_and_n9, cell_1983_a_HPC2_and_n8,
         cell_1983_a_HPC2_and_n7, cell_1983_a_HPC2_and_p_0_out_0__1_,
         cell_1983_a_HPC2_and_p_0_out_1__0_,
         cell_1983_a_HPC2_and_p_1_out_0__1_,
         cell_1983_a_HPC2_and_p_1_out_1__0_,
         cell_1983_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1983_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1983_a_HPC2_and_p_1_in_0__1_, cell_1983_a_HPC2_and_p_1_in_1__0_,
         cell_1983_a_HPC2_and_s_out_0__1_, cell_1983_a_HPC2_and_s_out_1__0_,
         cell_1983_a_HPC2_and_p_0_in_0__1_, cell_1983_a_HPC2_and_p_0_in_1__0_,
         cell_1983_a_HPC2_and_s_in_0__1_, cell_1983_a_HPC2_and_s_in_1__0_,
         cell_1983_a_HPC2_and_z_0__0_, cell_1983_a_HPC2_and_z_1__1_,
         cell_1984_a_HPC2_and_n9, cell_1984_a_HPC2_and_n8,
         cell_1984_a_HPC2_and_n7, cell_1984_a_HPC2_and_p_0_out_0__1_,
         cell_1984_a_HPC2_and_p_0_out_1__0_,
         cell_1984_a_HPC2_and_p_1_out_0__1_,
         cell_1984_a_HPC2_and_p_1_out_1__0_,
         cell_1984_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1984_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1984_a_HPC2_and_p_1_in_0__1_, cell_1984_a_HPC2_and_p_1_in_1__0_,
         cell_1984_a_HPC2_and_s_out_0__1_, cell_1984_a_HPC2_and_s_out_1__0_,
         cell_1984_a_HPC2_and_p_0_in_0__1_, cell_1984_a_HPC2_and_p_0_in_1__0_,
         cell_1984_a_HPC2_and_s_in_0__1_, cell_1984_a_HPC2_and_s_in_1__0_,
         cell_1984_a_HPC2_and_z_0__0_, cell_1984_a_HPC2_and_z_1__1_,
         cell_1985_a_HPC2_and_n9, cell_1985_a_HPC2_and_n8,
         cell_1985_a_HPC2_and_n7, cell_1985_a_HPC2_and_p_0_out_0__1_,
         cell_1985_a_HPC2_and_p_0_out_1__0_,
         cell_1985_a_HPC2_and_p_1_out_0__1_,
         cell_1985_a_HPC2_and_p_1_out_1__0_,
         cell_1985_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1985_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1985_a_HPC2_and_p_1_in_0__1_, cell_1985_a_HPC2_and_p_1_in_1__0_,
         cell_1985_a_HPC2_and_s_out_0__1_, cell_1985_a_HPC2_and_s_out_1__0_,
         cell_1985_a_HPC2_and_p_0_in_0__1_, cell_1985_a_HPC2_and_p_0_in_1__0_,
         cell_1985_a_HPC2_and_s_in_0__1_, cell_1985_a_HPC2_and_s_in_1__0_,
         cell_1985_a_HPC2_and_z_0__0_, cell_1985_a_HPC2_and_z_1__1_,
         cell_1986_a_HPC2_and_n9, cell_1986_a_HPC2_and_n8,
         cell_1986_a_HPC2_and_n7, cell_1986_a_HPC2_and_p_0_out_0__1_,
         cell_1986_a_HPC2_and_p_0_out_1__0_,
         cell_1986_a_HPC2_and_p_1_out_0__1_,
         cell_1986_a_HPC2_and_p_1_out_1__0_,
         cell_1986_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1986_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1986_a_HPC2_and_p_1_in_0__1_, cell_1986_a_HPC2_and_p_1_in_1__0_,
         cell_1986_a_HPC2_and_s_out_0__1_, cell_1986_a_HPC2_and_s_out_1__0_,
         cell_1986_a_HPC2_and_p_0_in_0__1_, cell_1986_a_HPC2_and_p_0_in_1__0_,
         cell_1986_a_HPC2_and_s_in_0__1_, cell_1986_a_HPC2_and_s_in_1__0_,
         cell_1986_a_HPC2_and_z_0__0_, cell_1986_a_HPC2_and_z_1__1_,
         cell_1987_a_HPC2_and_n9, cell_1987_a_HPC2_and_n8,
         cell_1987_a_HPC2_and_n7, cell_1987_a_HPC2_and_p_0_out_0__1_,
         cell_1987_a_HPC2_and_p_0_out_1__0_,
         cell_1987_a_HPC2_and_p_1_out_0__1_,
         cell_1987_a_HPC2_and_p_1_out_1__0_,
         cell_1987_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1987_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1987_a_HPC2_and_p_1_in_0__1_, cell_1987_a_HPC2_and_p_1_in_1__0_,
         cell_1987_a_HPC2_and_s_out_0__1_, cell_1987_a_HPC2_and_s_out_1__0_,
         cell_1987_a_HPC2_and_p_0_in_0__1_, cell_1987_a_HPC2_and_p_0_in_1__0_,
         cell_1987_a_HPC2_and_s_in_0__1_, cell_1987_a_HPC2_and_s_in_1__0_,
         cell_1987_a_HPC2_and_z_0__0_, cell_1987_a_HPC2_and_z_1__1_,
         cell_1988_a_HPC2_and_n9, cell_1988_a_HPC2_and_n8,
         cell_1988_a_HPC2_and_n7, cell_1988_a_HPC2_and_p_0_out_0__1_,
         cell_1988_a_HPC2_and_p_0_out_1__0_,
         cell_1988_a_HPC2_and_p_1_out_0__1_,
         cell_1988_a_HPC2_and_p_1_out_1__0_,
         cell_1988_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1988_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1988_a_HPC2_and_p_1_in_0__1_, cell_1988_a_HPC2_and_p_1_in_1__0_,
         cell_1988_a_HPC2_and_s_out_0__1_, cell_1988_a_HPC2_and_s_out_1__0_,
         cell_1988_a_HPC2_and_p_0_in_0__1_, cell_1988_a_HPC2_and_p_0_in_1__0_,
         cell_1988_a_HPC2_and_s_in_0__1_, cell_1988_a_HPC2_and_s_in_1__0_,
         cell_1988_a_HPC2_and_z_0__0_, cell_1988_a_HPC2_and_z_1__1_,
         cell_1989_a_HPC2_and_n9, cell_1989_a_HPC2_and_n8,
         cell_1989_a_HPC2_and_n7, cell_1989_a_HPC2_and_p_0_out_0__1_,
         cell_1989_a_HPC2_and_p_0_out_1__0_,
         cell_1989_a_HPC2_and_p_1_out_0__1_,
         cell_1989_a_HPC2_and_p_1_out_1__0_,
         cell_1989_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1989_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1989_a_HPC2_and_p_1_in_0__1_, cell_1989_a_HPC2_and_p_1_in_1__0_,
         cell_1989_a_HPC2_and_s_out_0__1_, cell_1989_a_HPC2_and_s_out_1__0_,
         cell_1989_a_HPC2_and_p_0_in_0__1_, cell_1989_a_HPC2_and_p_0_in_1__0_,
         cell_1989_a_HPC2_and_s_in_0__1_, cell_1989_a_HPC2_and_s_in_1__0_,
         cell_1989_a_HPC2_and_z_0__0_, cell_1989_a_HPC2_and_z_1__1_,
         cell_1990_a_HPC2_and_n9, cell_1990_a_HPC2_and_n8,
         cell_1990_a_HPC2_and_n7, cell_1990_a_HPC2_and_p_0_out_0__1_,
         cell_1990_a_HPC2_and_p_0_out_1__0_,
         cell_1990_a_HPC2_and_p_1_out_0__1_,
         cell_1990_a_HPC2_and_p_1_out_1__0_,
         cell_1990_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1990_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1990_a_HPC2_and_p_1_in_0__1_, cell_1990_a_HPC2_and_p_1_in_1__0_,
         cell_1990_a_HPC2_and_s_out_0__1_, cell_1990_a_HPC2_and_s_out_1__0_,
         cell_1990_a_HPC2_and_p_0_in_0__1_, cell_1990_a_HPC2_and_p_0_in_1__0_,
         cell_1990_a_HPC2_and_s_in_0__1_, cell_1990_a_HPC2_and_s_in_1__0_,
         cell_1990_a_HPC2_and_z_0__0_, cell_1990_a_HPC2_and_z_1__1_,
         cell_1991_a_HPC2_and_n9, cell_1991_a_HPC2_and_n8,
         cell_1991_a_HPC2_and_n7, cell_1991_a_HPC2_and_p_0_out_0__1_,
         cell_1991_a_HPC2_and_p_0_out_1__0_,
         cell_1991_a_HPC2_and_p_1_out_0__1_,
         cell_1991_a_HPC2_and_p_1_out_1__0_,
         cell_1991_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1991_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1991_a_HPC2_and_p_1_in_0__1_, cell_1991_a_HPC2_and_p_1_in_1__0_,
         cell_1991_a_HPC2_and_s_out_0__1_, cell_1991_a_HPC2_and_s_out_1__0_,
         cell_1991_a_HPC2_and_p_0_in_0__1_, cell_1991_a_HPC2_and_p_0_in_1__0_,
         cell_1991_a_HPC2_and_s_in_0__1_, cell_1991_a_HPC2_and_s_in_1__0_,
         cell_1991_a_HPC2_and_z_0__0_, cell_1991_a_HPC2_and_z_1__1_,
         cell_1992_a_HPC2_and_n9, cell_1992_a_HPC2_and_n8,
         cell_1992_a_HPC2_and_n7, cell_1992_a_HPC2_and_p_0_out_0__1_,
         cell_1992_a_HPC2_and_p_0_out_1__0_,
         cell_1992_a_HPC2_and_p_1_out_0__1_,
         cell_1992_a_HPC2_and_p_1_out_1__0_,
         cell_1992_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1992_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1992_a_HPC2_and_p_1_in_0__1_, cell_1992_a_HPC2_and_p_1_in_1__0_,
         cell_1992_a_HPC2_and_s_out_0__1_, cell_1992_a_HPC2_and_s_out_1__0_,
         cell_1992_a_HPC2_and_p_0_in_0__1_, cell_1992_a_HPC2_and_p_0_in_1__0_,
         cell_1992_a_HPC2_and_s_in_0__1_, cell_1992_a_HPC2_and_s_in_1__0_,
         cell_1992_a_HPC2_and_z_0__0_, cell_1992_a_HPC2_and_z_1__1_,
         cell_1993_a_HPC2_and_n9, cell_1993_a_HPC2_and_n8,
         cell_1993_a_HPC2_and_n7, cell_1993_a_HPC2_and_p_0_out_0__1_,
         cell_1993_a_HPC2_and_p_0_out_1__0_,
         cell_1993_a_HPC2_and_p_1_out_0__1_,
         cell_1993_a_HPC2_and_p_1_out_1__0_,
         cell_1993_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1993_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1993_a_HPC2_and_p_1_in_0__1_, cell_1993_a_HPC2_and_p_1_in_1__0_,
         cell_1993_a_HPC2_and_s_out_0__1_, cell_1993_a_HPC2_and_s_out_1__0_,
         cell_1993_a_HPC2_and_p_0_in_0__1_, cell_1993_a_HPC2_and_p_0_in_1__0_,
         cell_1993_a_HPC2_and_s_in_0__1_, cell_1993_a_HPC2_and_s_in_1__0_,
         cell_1993_a_HPC2_and_z_0__0_, cell_1993_a_HPC2_and_z_1__1_,
         cell_1994_a_HPC2_and_n9, cell_1994_a_HPC2_and_n8,
         cell_1994_a_HPC2_and_n7, cell_1994_a_HPC2_and_p_0_out_0__1_,
         cell_1994_a_HPC2_and_p_0_out_1__0_,
         cell_1994_a_HPC2_and_p_1_out_0__1_,
         cell_1994_a_HPC2_and_p_1_out_1__0_,
         cell_1994_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1994_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1994_a_HPC2_and_p_1_in_0__1_, cell_1994_a_HPC2_and_p_1_in_1__0_,
         cell_1994_a_HPC2_and_s_out_0__1_, cell_1994_a_HPC2_and_s_out_1__0_,
         cell_1994_a_HPC2_and_p_0_in_0__1_, cell_1994_a_HPC2_and_p_0_in_1__0_,
         cell_1994_a_HPC2_and_s_in_0__1_, cell_1994_a_HPC2_and_s_in_1__0_,
         cell_1994_a_HPC2_and_z_0__0_, cell_1994_a_HPC2_and_z_1__1_,
         cell_1995_a_HPC2_and_n9, cell_1995_a_HPC2_and_n8,
         cell_1995_a_HPC2_and_n7, cell_1995_a_HPC2_and_p_0_out_0__1_,
         cell_1995_a_HPC2_and_p_0_out_1__0_,
         cell_1995_a_HPC2_and_p_1_out_0__1_,
         cell_1995_a_HPC2_and_p_1_out_1__0_,
         cell_1995_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1995_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1995_a_HPC2_and_p_1_in_0__1_, cell_1995_a_HPC2_and_p_1_in_1__0_,
         cell_1995_a_HPC2_and_s_out_0__1_, cell_1995_a_HPC2_and_s_out_1__0_,
         cell_1995_a_HPC2_and_p_0_in_0__1_, cell_1995_a_HPC2_and_p_0_in_1__0_,
         cell_1995_a_HPC2_and_s_in_0__1_, cell_1995_a_HPC2_and_s_in_1__0_,
         cell_1995_a_HPC2_and_z_0__0_, cell_1995_a_HPC2_and_z_1__1_,
         cell_1996_a_HPC2_and_n9, cell_1996_a_HPC2_and_n8,
         cell_1996_a_HPC2_and_n7, cell_1996_a_HPC2_and_p_0_out_0__1_,
         cell_1996_a_HPC2_and_p_0_out_1__0_,
         cell_1996_a_HPC2_and_p_1_out_0__1_,
         cell_1996_a_HPC2_and_p_1_out_1__0_,
         cell_1996_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1996_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1996_a_HPC2_and_p_1_in_0__1_, cell_1996_a_HPC2_and_p_1_in_1__0_,
         cell_1996_a_HPC2_and_s_out_0__1_, cell_1996_a_HPC2_and_s_out_1__0_,
         cell_1996_a_HPC2_and_p_0_in_0__1_, cell_1996_a_HPC2_and_p_0_in_1__0_,
         cell_1996_a_HPC2_and_s_in_0__1_, cell_1996_a_HPC2_and_s_in_1__0_,
         cell_1996_a_HPC2_and_z_0__0_, cell_1996_a_HPC2_and_z_1__1_,
         cell_1997_a_HPC2_and_n9, cell_1997_a_HPC2_and_n8,
         cell_1997_a_HPC2_and_n7, cell_1997_a_HPC2_and_p_0_out_0__1_,
         cell_1997_a_HPC2_and_p_0_out_1__0_,
         cell_1997_a_HPC2_and_p_1_out_0__1_,
         cell_1997_a_HPC2_and_p_1_out_1__0_,
         cell_1997_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1997_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1997_a_HPC2_and_p_1_in_0__1_, cell_1997_a_HPC2_and_p_1_in_1__0_,
         cell_1997_a_HPC2_and_s_out_0__1_, cell_1997_a_HPC2_and_s_out_1__0_,
         cell_1997_a_HPC2_and_p_0_in_0__1_, cell_1997_a_HPC2_and_p_0_in_1__0_,
         cell_1997_a_HPC2_and_s_in_0__1_, cell_1997_a_HPC2_and_s_in_1__0_,
         cell_1997_a_HPC2_and_z_0__0_, cell_1997_a_HPC2_and_z_1__1_,
         cell_1998_a_HPC2_and_n9, cell_1998_a_HPC2_and_n8,
         cell_1998_a_HPC2_and_n7, cell_1998_a_HPC2_and_p_0_out_0__1_,
         cell_1998_a_HPC2_and_p_0_out_1__0_,
         cell_1998_a_HPC2_and_p_1_out_0__1_,
         cell_1998_a_HPC2_and_p_1_out_1__0_,
         cell_1998_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1998_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1998_a_HPC2_and_p_1_in_0__1_, cell_1998_a_HPC2_and_p_1_in_1__0_,
         cell_1998_a_HPC2_and_s_out_0__1_, cell_1998_a_HPC2_and_s_out_1__0_,
         cell_1998_a_HPC2_and_p_0_in_0__1_, cell_1998_a_HPC2_and_p_0_in_1__0_,
         cell_1998_a_HPC2_and_s_in_0__1_, cell_1998_a_HPC2_and_s_in_1__0_,
         cell_1998_a_HPC2_and_z_0__0_, cell_1998_a_HPC2_and_z_1__1_,
         cell_1999_a_HPC2_and_n9, cell_1999_a_HPC2_and_n8,
         cell_1999_a_HPC2_and_n7, cell_1999_a_HPC2_and_p_0_out_0__1_,
         cell_1999_a_HPC2_and_p_0_out_1__0_,
         cell_1999_a_HPC2_and_p_1_out_0__1_,
         cell_1999_a_HPC2_and_p_1_out_1__0_,
         cell_1999_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_1999_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_1999_a_HPC2_and_p_1_in_0__1_, cell_1999_a_HPC2_and_p_1_in_1__0_,
         cell_1999_a_HPC2_and_s_out_0__1_, cell_1999_a_HPC2_and_s_out_1__0_,
         cell_1999_a_HPC2_and_p_0_in_0__1_, cell_1999_a_HPC2_and_p_0_in_1__0_,
         cell_1999_a_HPC2_and_s_in_0__1_, cell_1999_a_HPC2_and_s_in_1__0_,
         cell_1999_a_HPC2_and_z_0__0_, cell_1999_a_HPC2_and_z_1__1_,
         cell_2000_a_HPC2_and_n9, cell_2000_a_HPC2_and_n8,
         cell_2000_a_HPC2_and_n7, cell_2000_a_HPC2_and_p_0_out_0__1_,
         cell_2000_a_HPC2_and_p_0_out_1__0_,
         cell_2000_a_HPC2_and_p_1_out_0__1_,
         cell_2000_a_HPC2_and_p_1_out_1__0_,
         cell_2000_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2000_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2000_a_HPC2_and_p_1_in_0__1_, cell_2000_a_HPC2_and_p_1_in_1__0_,
         cell_2000_a_HPC2_and_s_out_0__1_, cell_2000_a_HPC2_and_s_out_1__0_,
         cell_2000_a_HPC2_and_p_0_in_0__1_, cell_2000_a_HPC2_and_p_0_in_1__0_,
         cell_2000_a_HPC2_and_s_in_0__1_, cell_2000_a_HPC2_and_s_in_1__0_,
         cell_2000_a_HPC2_and_z_0__0_, cell_2000_a_HPC2_and_z_1__1_,
         cell_2001_a_HPC2_and_n9, cell_2001_a_HPC2_and_n8,
         cell_2001_a_HPC2_and_n7, cell_2001_a_HPC2_and_p_0_out_0__1_,
         cell_2001_a_HPC2_and_p_0_out_1__0_,
         cell_2001_a_HPC2_and_p_1_out_0__1_,
         cell_2001_a_HPC2_and_p_1_out_1__0_,
         cell_2001_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2001_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2001_a_HPC2_and_p_1_in_0__1_, cell_2001_a_HPC2_and_p_1_in_1__0_,
         cell_2001_a_HPC2_and_s_out_0__1_, cell_2001_a_HPC2_and_s_out_1__0_,
         cell_2001_a_HPC2_and_p_0_in_0__1_, cell_2001_a_HPC2_and_p_0_in_1__0_,
         cell_2001_a_HPC2_and_s_in_0__1_, cell_2001_a_HPC2_and_s_in_1__0_,
         cell_2001_a_HPC2_and_z_0__0_, cell_2001_a_HPC2_and_z_1__1_,
         cell_2002_a_HPC2_and_n9, cell_2002_a_HPC2_and_n8,
         cell_2002_a_HPC2_and_n7, cell_2002_a_HPC2_and_p_0_out_0__1_,
         cell_2002_a_HPC2_and_p_0_out_1__0_,
         cell_2002_a_HPC2_and_p_1_out_0__1_,
         cell_2002_a_HPC2_and_p_1_out_1__0_,
         cell_2002_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2002_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2002_a_HPC2_and_p_1_in_0__1_, cell_2002_a_HPC2_and_p_1_in_1__0_,
         cell_2002_a_HPC2_and_s_out_0__1_, cell_2002_a_HPC2_and_s_out_1__0_,
         cell_2002_a_HPC2_and_p_0_in_0__1_, cell_2002_a_HPC2_and_p_0_in_1__0_,
         cell_2002_a_HPC2_and_s_in_0__1_, cell_2002_a_HPC2_and_s_in_1__0_,
         cell_2002_a_HPC2_and_z_0__0_, cell_2002_a_HPC2_and_z_1__1_,
         cell_2003_a_HPC2_and_n9, cell_2003_a_HPC2_and_n8,
         cell_2003_a_HPC2_and_n7, cell_2003_a_HPC2_and_p_0_out_0__1_,
         cell_2003_a_HPC2_and_p_0_out_1__0_,
         cell_2003_a_HPC2_and_p_1_out_0__1_,
         cell_2003_a_HPC2_and_p_1_out_1__0_,
         cell_2003_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2003_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2003_a_HPC2_and_p_1_in_0__1_, cell_2003_a_HPC2_and_p_1_in_1__0_,
         cell_2003_a_HPC2_and_s_out_0__1_, cell_2003_a_HPC2_and_s_out_1__0_,
         cell_2003_a_HPC2_and_p_0_in_0__1_, cell_2003_a_HPC2_and_p_0_in_1__0_,
         cell_2003_a_HPC2_and_s_in_0__1_, cell_2003_a_HPC2_and_s_in_1__0_,
         cell_2003_a_HPC2_and_z_0__0_, cell_2003_a_HPC2_and_z_1__1_,
         cell_2004_a_HPC2_and_n9, cell_2004_a_HPC2_and_n8,
         cell_2004_a_HPC2_and_n7, cell_2004_a_HPC2_and_p_0_out_0__1_,
         cell_2004_a_HPC2_and_p_0_out_1__0_,
         cell_2004_a_HPC2_and_p_1_out_0__1_,
         cell_2004_a_HPC2_and_p_1_out_1__0_,
         cell_2004_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2004_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2004_a_HPC2_and_p_1_in_0__1_, cell_2004_a_HPC2_and_p_1_in_1__0_,
         cell_2004_a_HPC2_and_s_out_0__1_, cell_2004_a_HPC2_and_s_out_1__0_,
         cell_2004_a_HPC2_and_p_0_in_0__1_, cell_2004_a_HPC2_and_p_0_in_1__0_,
         cell_2004_a_HPC2_and_s_in_0__1_, cell_2004_a_HPC2_and_s_in_1__0_,
         cell_2004_a_HPC2_and_z_0__0_, cell_2004_a_HPC2_and_z_1__1_,
         cell_2005_a_HPC2_and_n9, cell_2005_a_HPC2_and_n8,
         cell_2005_a_HPC2_and_n7, cell_2005_a_HPC2_and_p_0_out_0__1_,
         cell_2005_a_HPC2_and_p_0_out_1__0_,
         cell_2005_a_HPC2_and_p_1_out_0__1_,
         cell_2005_a_HPC2_and_p_1_out_1__0_,
         cell_2005_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2005_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2005_a_HPC2_and_p_1_in_0__1_, cell_2005_a_HPC2_and_p_1_in_1__0_,
         cell_2005_a_HPC2_and_s_out_0__1_, cell_2005_a_HPC2_and_s_out_1__0_,
         cell_2005_a_HPC2_and_p_0_in_0__1_, cell_2005_a_HPC2_and_p_0_in_1__0_,
         cell_2005_a_HPC2_and_s_in_0__1_, cell_2005_a_HPC2_and_s_in_1__0_,
         cell_2005_a_HPC2_and_z_0__0_, cell_2005_a_HPC2_and_z_1__1_,
         cell_2006_a_HPC2_and_n9, cell_2006_a_HPC2_and_n8,
         cell_2006_a_HPC2_and_n7, cell_2006_a_HPC2_and_p_0_out_0__1_,
         cell_2006_a_HPC2_and_p_0_out_1__0_,
         cell_2006_a_HPC2_and_p_1_out_0__1_,
         cell_2006_a_HPC2_and_p_1_out_1__0_,
         cell_2006_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2006_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2006_a_HPC2_and_p_1_in_0__1_, cell_2006_a_HPC2_and_p_1_in_1__0_,
         cell_2006_a_HPC2_and_s_out_0__1_, cell_2006_a_HPC2_and_s_out_1__0_,
         cell_2006_a_HPC2_and_p_0_in_0__1_, cell_2006_a_HPC2_and_p_0_in_1__0_,
         cell_2006_a_HPC2_and_s_in_0__1_, cell_2006_a_HPC2_and_s_in_1__0_,
         cell_2006_a_HPC2_and_z_0__0_, cell_2006_a_HPC2_and_z_1__1_,
         cell_2007_a_HPC2_and_n9, cell_2007_a_HPC2_and_n8,
         cell_2007_a_HPC2_and_n7, cell_2007_a_HPC2_and_p_0_out_0__1_,
         cell_2007_a_HPC2_and_p_0_out_1__0_,
         cell_2007_a_HPC2_and_p_1_out_0__1_,
         cell_2007_a_HPC2_and_p_1_out_1__0_,
         cell_2007_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2007_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2007_a_HPC2_and_p_1_in_0__1_, cell_2007_a_HPC2_and_p_1_in_1__0_,
         cell_2007_a_HPC2_and_s_out_0__1_, cell_2007_a_HPC2_and_s_out_1__0_,
         cell_2007_a_HPC2_and_p_0_in_0__1_, cell_2007_a_HPC2_and_p_0_in_1__0_,
         cell_2007_a_HPC2_and_s_in_0__1_, cell_2007_a_HPC2_and_s_in_1__0_,
         cell_2007_a_HPC2_and_z_0__0_, cell_2007_a_HPC2_and_z_1__1_,
         cell_2008_a_HPC2_and_n9, cell_2008_a_HPC2_and_n8,
         cell_2008_a_HPC2_and_n7, cell_2008_a_HPC2_and_p_0_out_0__1_,
         cell_2008_a_HPC2_and_p_0_out_1__0_,
         cell_2008_a_HPC2_and_p_1_out_0__1_,
         cell_2008_a_HPC2_and_p_1_out_1__0_,
         cell_2008_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2008_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2008_a_HPC2_and_p_1_in_0__1_, cell_2008_a_HPC2_and_p_1_in_1__0_,
         cell_2008_a_HPC2_and_s_out_0__1_, cell_2008_a_HPC2_and_s_out_1__0_,
         cell_2008_a_HPC2_and_p_0_in_0__1_, cell_2008_a_HPC2_and_p_0_in_1__0_,
         cell_2008_a_HPC2_and_s_in_0__1_, cell_2008_a_HPC2_and_s_in_1__0_,
         cell_2008_a_HPC2_and_z_0__0_, cell_2008_a_HPC2_and_z_1__1_,
         cell_2009_a_HPC2_and_n9, cell_2009_a_HPC2_and_n8,
         cell_2009_a_HPC2_and_n7, cell_2009_a_HPC2_and_p_0_out_0__1_,
         cell_2009_a_HPC2_and_p_0_out_1__0_,
         cell_2009_a_HPC2_and_p_1_out_0__1_,
         cell_2009_a_HPC2_and_p_1_out_1__0_,
         cell_2009_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2009_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2009_a_HPC2_and_p_1_in_0__1_, cell_2009_a_HPC2_and_p_1_in_1__0_,
         cell_2009_a_HPC2_and_s_out_0__1_, cell_2009_a_HPC2_and_s_out_1__0_,
         cell_2009_a_HPC2_and_p_0_in_0__1_, cell_2009_a_HPC2_and_p_0_in_1__0_,
         cell_2009_a_HPC2_and_s_in_0__1_, cell_2009_a_HPC2_and_s_in_1__0_,
         cell_2009_a_HPC2_and_z_0__0_, cell_2009_a_HPC2_and_z_1__1_,
         cell_2010_a_HPC2_and_n9, cell_2010_a_HPC2_and_n8,
         cell_2010_a_HPC2_and_n7, cell_2010_a_HPC2_and_p_0_out_0__1_,
         cell_2010_a_HPC2_and_p_0_out_1__0_,
         cell_2010_a_HPC2_and_p_1_out_0__1_,
         cell_2010_a_HPC2_and_p_1_out_1__0_,
         cell_2010_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2010_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2010_a_HPC2_and_p_1_in_0__1_, cell_2010_a_HPC2_and_p_1_in_1__0_,
         cell_2010_a_HPC2_and_s_out_0__1_, cell_2010_a_HPC2_and_s_out_1__0_,
         cell_2010_a_HPC2_and_p_0_in_0__1_, cell_2010_a_HPC2_and_p_0_in_1__0_,
         cell_2010_a_HPC2_and_s_in_0__1_, cell_2010_a_HPC2_and_s_in_1__0_,
         cell_2010_a_HPC2_and_z_0__0_, cell_2010_a_HPC2_and_z_1__1_,
         cell_2011_a_HPC2_and_n9, cell_2011_a_HPC2_and_n8,
         cell_2011_a_HPC2_and_n7, cell_2011_a_HPC2_and_p_0_out_0__1_,
         cell_2011_a_HPC2_and_p_0_out_1__0_,
         cell_2011_a_HPC2_and_p_1_out_0__1_,
         cell_2011_a_HPC2_and_p_1_out_1__0_,
         cell_2011_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2011_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2011_a_HPC2_and_p_1_in_0__1_, cell_2011_a_HPC2_and_p_1_in_1__0_,
         cell_2011_a_HPC2_and_s_out_0__1_, cell_2011_a_HPC2_and_s_out_1__0_,
         cell_2011_a_HPC2_and_p_0_in_0__1_, cell_2011_a_HPC2_and_p_0_in_1__0_,
         cell_2011_a_HPC2_and_s_in_0__1_, cell_2011_a_HPC2_and_s_in_1__0_,
         cell_2011_a_HPC2_and_z_0__0_, cell_2011_a_HPC2_and_z_1__1_,
         cell_2012_a_HPC2_and_n9, cell_2012_a_HPC2_and_n8,
         cell_2012_a_HPC2_and_n7, cell_2012_a_HPC2_and_p_0_out_0__1_,
         cell_2012_a_HPC2_and_p_0_out_1__0_,
         cell_2012_a_HPC2_and_p_1_out_0__1_,
         cell_2012_a_HPC2_and_p_1_out_1__0_,
         cell_2012_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2012_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2012_a_HPC2_and_p_1_in_0__1_, cell_2012_a_HPC2_and_p_1_in_1__0_,
         cell_2012_a_HPC2_and_s_out_0__1_, cell_2012_a_HPC2_and_s_out_1__0_,
         cell_2012_a_HPC2_and_p_0_in_0__1_, cell_2012_a_HPC2_and_p_0_in_1__0_,
         cell_2012_a_HPC2_and_s_in_0__1_, cell_2012_a_HPC2_and_s_in_1__0_,
         cell_2012_a_HPC2_and_z_0__0_, cell_2012_a_HPC2_and_z_1__1_,
         cell_2013_a_HPC2_and_n9, cell_2013_a_HPC2_and_n8,
         cell_2013_a_HPC2_and_n7, cell_2013_a_HPC2_and_p_0_out_0__1_,
         cell_2013_a_HPC2_and_p_0_out_1__0_,
         cell_2013_a_HPC2_and_p_1_out_0__1_,
         cell_2013_a_HPC2_and_p_1_out_1__0_,
         cell_2013_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2013_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2013_a_HPC2_and_p_1_in_0__1_, cell_2013_a_HPC2_and_p_1_in_1__0_,
         cell_2013_a_HPC2_and_s_out_0__1_, cell_2013_a_HPC2_and_s_out_1__0_,
         cell_2013_a_HPC2_and_p_0_in_0__1_, cell_2013_a_HPC2_and_p_0_in_1__0_,
         cell_2013_a_HPC2_and_s_in_0__1_, cell_2013_a_HPC2_and_s_in_1__0_,
         cell_2013_a_HPC2_and_z_0__0_, cell_2013_a_HPC2_and_z_1__1_,
         cell_2014_a_HPC2_and_n9, cell_2014_a_HPC2_and_n8,
         cell_2014_a_HPC2_and_n7, cell_2014_a_HPC2_and_p_0_out_0__1_,
         cell_2014_a_HPC2_and_p_0_out_1__0_,
         cell_2014_a_HPC2_and_p_1_out_0__1_,
         cell_2014_a_HPC2_and_p_1_out_1__0_,
         cell_2014_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2014_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2014_a_HPC2_and_p_1_in_0__1_, cell_2014_a_HPC2_and_p_1_in_1__0_,
         cell_2014_a_HPC2_and_s_out_0__1_, cell_2014_a_HPC2_and_s_out_1__0_,
         cell_2014_a_HPC2_and_p_0_in_0__1_, cell_2014_a_HPC2_and_p_0_in_1__0_,
         cell_2014_a_HPC2_and_s_in_0__1_, cell_2014_a_HPC2_and_s_in_1__0_,
         cell_2014_a_HPC2_and_z_0__0_, cell_2014_a_HPC2_and_z_1__1_,
         cell_2015_a_HPC2_and_n9, cell_2015_a_HPC2_and_n8,
         cell_2015_a_HPC2_and_n7, cell_2015_a_HPC2_and_p_0_out_0__1_,
         cell_2015_a_HPC2_and_p_0_out_1__0_,
         cell_2015_a_HPC2_and_p_1_out_0__1_,
         cell_2015_a_HPC2_and_p_1_out_1__0_,
         cell_2015_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2015_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2015_a_HPC2_and_p_1_in_0__1_, cell_2015_a_HPC2_and_p_1_in_1__0_,
         cell_2015_a_HPC2_and_s_out_0__1_, cell_2015_a_HPC2_and_s_out_1__0_,
         cell_2015_a_HPC2_and_p_0_in_0__1_, cell_2015_a_HPC2_and_p_0_in_1__0_,
         cell_2015_a_HPC2_and_s_in_0__1_, cell_2015_a_HPC2_and_s_in_1__0_,
         cell_2015_a_HPC2_and_z_0__0_, cell_2015_a_HPC2_and_z_1__1_,
         cell_2016_a_HPC2_and_n9, cell_2016_a_HPC2_and_n8,
         cell_2016_a_HPC2_and_n7, cell_2016_a_HPC2_and_p_0_out_0__1_,
         cell_2016_a_HPC2_and_p_0_out_1__0_,
         cell_2016_a_HPC2_and_p_1_out_0__1_,
         cell_2016_a_HPC2_and_p_1_out_1__0_,
         cell_2016_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2016_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2016_a_HPC2_and_p_1_in_0__1_, cell_2016_a_HPC2_and_p_1_in_1__0_,
         cell_2016_a_HPC2_and_s_out_0__1_, cell_2016_a_HPC2_and_s_out_1__0_,
         cell_2016_a_HPC2_and_p_0_in_0__1_, cell_2016_a_HPC2_and_p_0_in_1__0_,
         cell_2016_a_HPC2_and_s_in_0__1_, cell_2016_a_HPC2_and_s_in_1__0_,
         cell_2016_a_HPC2_and_z_0__0_, cell_2016_a_HPC2_and_z_1__1_,
         cell_2017_a_HPC2_and_n9, cell_2017_a_HPC2_and_n8,
         cell_2017_a_HPC2_and_n7, cell_2017_a_HPC2_and_p_0_out_0__1_,
         cell_2017_a_HPC2_and_p_0_out_1__0_,
         cell_2017_a_HPC2_and_p_1_out_0__1_,
         cell_2017_a_HPC2_and_p_1_out_1__0_,
         cell_2017_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2017_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2017_a_HPC2_and_p_1_in_0__1_, cell_2017_a_HPC2_and_p_1_in_1__0_,
         cell_2017_a_HPC2_and_s_out_0__1_, cell_2017_a_HPC2_and_s_out_1__0_,
         cell_2017_a_HPC2_and_p_0_in_0__1_, cell_2017_a_HPC2_and_p_0_in_1__0_,
         cell_2017_a_HPC2_and_s_in_0__1_, cell_2017_a_HPC2_and_s_in_1__0_,
         cell_2017_a_HPC2_and_z_0__0_, cell_2017_a_HPC2_and_z_1__1_,
         cell_2018_a_HPC2_and_n9, cell_2018_a_HPC2_and_n8,
         cell_2018_a_HPC2_and_n7, cell_2018_a_HPC2_and_p_0_out_0__1_,
         cell_2018_a_HPC2_and_p_0_out_1__0_,
         cell_2018_a_HPC2_and_p_1_out_0__1_,
         cell_2018_a_HPC2_and_p_1_out_1__0_,
         cell_2018_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2018_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2018_a_HPC2_and_p_1_in_0__1_, cell_2018_a_HPC2_and_p_1_in_1__0_,
         cell_2018_a_HPC2_and_s_out_0__1_, cell_2018_a_HPC2_and_s_out_1__0_,
         cell_2018_a_HPC2_and_p_0_in_0__1_, cell_2018_a_HPC2_and_p_0_in_1__0_,
         cell_2018_a_HPC2_and_s_in_0__1_, cell_2018_a_HPC2_and_s_in_1__0_,
         cell_2018_a_HPC2_and_z_0__0_, cell_2018_a_HPC2_and_z_1__1_,
         cell_2019_a_HPC2_and_n9, cell_2019_a_HPC2_and_n8,
         cell_2019_a_HPC2_and_n7, cell_2019_a_HPC2_and_p_0_out_0__1_,
         cell_2019_a_HPC2_and_p_0_out_1__0_,
         cell_2019_a_HPC2_and_p_1_out_0__1_,
         cell_2019_a_HPC2_and_p_1_out_1__0_,
         cell_2019_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2019_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2019_a_HPC2_and_p_1_in_0__1_, cell_2019_a_HPC2_and_p_1_in_1__0_,
         cell_2019_a_HPC2_and_s_out_0__1_, cell_2019_a_HPC2_and_s_out_1__0_,
         cell_2019_a_HPC2_and_p_0_in_0__1_, cell_2019_a_HPC2_and_p_0_in_1__0_,
         cell_2019_a_HPC2_and_s_in_0__1_, cell_2019_a_HPC2_and_s_in_1__0_,
         cell_2019_a_HPC2_and_z_0__0_, cell_2019_a_HPC2_and_z_1__1_,
         cell_2020_a_HPC2_and_n9, cell_2020_a_HPC2_and_n8,
         cell_2020_a_HPC2_and_n7, cell_2020_a_HPC2_and_p_0_out_0__1_,
         cell_2020_a_HPC2_and_p_0_out_1__0_,
         cell_2020_a_HPC2_and_p_1_out_0__1_,
         cell_2020_a_HPC2_and_p_1_out_1__0_,
         cell_2020_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2020_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2020_a_HPC2_and_p_1_in_0__1_, cell_2020_a_HPC2_and_p_1_in_1__0_,
         cell_2020_a_HPC2_and_s_out_0__1_, cell_2020_a_HPC2_and_s_out_1__0_,
         cell_2020_a_HPC2_and_p_0_in_0__1_, cell_2020_a_HPC2_and_p_0_in_1__0_,
         cell_2020_a_HPC2_and_s_in_0__1_, cell_2020_a_HPC2_and_s_in_1__0_,
         cell_2020_a_HPC2_and_z_0__0_, cell_2020_a_HPC2_and_z_1__1_,
         cell_2021_a_HPC2_and_n9, cell_2021_a_HPC2_and_n8,
         cell_2021_a_HPC2_and_n7, cell_2021_a_HPC2_and_p_0_out_0__1_,
         cell_2021_a_HPC2_and_p_0_out_1__0_,
         cell_2021_a_HPC2_and_p_1_out_0__1_,
         cell_2021_a_HPC2_and_p_1_out_1__0_,
         cell_2021_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2021_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2021_a_HPC2_and_p_1_in_0__1_, cell_2021_a_HPC2_and_p_1_in_1__0_,
         cell_2021_a_HPC2_and_s_out_0__1_, cell_2021_a_HPC2_and_s_out_1__0_,
         cell_2021_a_HPC2_and_p_0_in_0__1_, cell_2021_a_HPC2_and_p_0_in_1__0_,
         cell_2021_a_HPC2_and_s_in_0__1_, cell_2021_a_HPC2_and_s_in_1__0_,
         cell_2021_a_HPC2_and_z_0__0_, cell_2021_a_HPC2_and_z_1__1_,
         cell_2022_a_HPC2_and_n9, cell_2022_a_HPC2_and_n8,
         cell_2022_a_HPC2_and_n7, cell_2022_a_HPC2_and_p_0_out_0__1_,
         cell_2022_a_HPC2_and_p_0_out_1__0_,
         cell_2022_a_HPC2_and_p_1_out_0__1_,
         cell_2022_a_HPC2_and_p_1_out_1__0_,
         cell_2022_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2022_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2022_a_HPC2_and_p_1_in_0__1_, cell_2022_a_HPC2_and_p_1_in_1__0_,
         cell_2022_a_HPC2_and_s_out_0__1_, cell_2022_a_HPC2_and_s_out_1__0_,
         cell_2022_a_HPC2_and_p_0_in_0__1_, cell_2022_a_HPC2_and_p_0_in_1__0_,
         cell_2022_a_HPC2_and_s_in_0__1_, cell_2022_a_HPC2_and_s_in_1__0_,
         cell_2022_a_HPC2_and_z_0__0_, cell_2022_a_HPC2_and_z_1__1_,
         cell_2023_a_HPC2_and_n9, cell_2023_a_HPC2_and_n8,
         cell_2023_a_HPC2_and_n7, cell_2023_a_HPC2_and_p_0_out_0__1_,
         cell_2023_a_HPC2_and_p_0_out_1__0_,
         cell_2023_a_HPC2_and_p_1_out_0__1_,
         cell_2023_a_HPC2_and_p_1_out_1__0_,
         cell_2023_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2023_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2023_a_HPC2_and_p_1_in_0__1_, cell_2023_a_HPC2_and_p_1_in_1__0_,
         cell_2023_a_HPC2_and_s_out_0__1_, cell_2023_a_HPC2_and_s_out_1__0_,
         cell_2023_a_HPC2_and_p_0_in_0__1_, cell_2023_a_HPC2_and_p_0_in_1__0_,
         cell_2023_a_HPC2_and_s_in_0__1_, cell_2023_a_HPC2_and_s_in_1__0_,
         cell_2023_a_HPC2_and_z_0__0_, cell_2023_a_HPC2_and_z_1__1_,
         cell_2024_a_HPC2_and_n9, cell_2024_a_HPC2_and_n8,
         cell_2024_a_HPC2_and_n7, cell_2024_a_HPC2_and_p_0_out_0__1_,
         cell_2024_a_HPC2_and_p_0_out_1__0_,
         cell_2024_a_HPC2_and_p_1_out_0__1_,
         cell_2024_a_HPC2_and_p_1_out_1__0_,
         cell_2024_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2024_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2024_a_HPC2_and_p_1_in_0__1_, cell_2024_a_HPC2_and_p_1_in_1__0_,
         cell_2024_a_HPC2_and_s_out_0__1_, cell_2024_a_HPC2_and_s_out_1__0_,
         cell_2024_a_HPC2_and_p_0_in_0__1_, cell_2024_a_HPC2_and_p_0_in_1__0_,
         cell_2024_a_HPC2_and_s_in_0__1_, cell_2024_a_HPC2_and_s_in_1__0_,
         cell_2024_a_HPC2_and_z_0__0_, cell_2024_a_HPC2_and_z_1__1_,
         cell_2025_a_HPC2_and_n9, cell_2025_a_HPC2_and_n8,
         cell_2025_a_HPC2_and_n7, cell_2025_a_HPC2_and_p_0_out_0__1_,
         cell_2025_a_HPC2_and_p_0_out_1__0_,
         cell_2025_a_HPC2_and_p_1_out_0__1_,
         cell_2025_a_HPC2_and_p_1_out_1__0_,
         cell_2025_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2025_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2025_a_HPC2_and_p_1_in_0__1_, cell_2025_a_HPC2_and_p_1_in_1__0_,
         cell_2025_a_HPC2_and_s_out_0__1_, cell_2025_a_HPC2_and_s_out_1__0_,
         cell_2025_a_HPC2_and_p_0_in_0__1_, cell_2025_a_HPC2_and_p_0_in_1__0_,
         cell_2025_a_HPC2_and_s_in_0__1_, cell_2025_a_HPC2_and_s_in_1__0_,
         cell_2025_a_HPC2_and_z_0__0_, cell_2025_a_HPC2_and_z_1__1_,
         cell_2026_a_HPC2_and_n9, cell_2026_a_HPC2_and_n8,
         cell_2026_a_HPC2_and_n7, cell_2026_a_HPC2_and_p_0_out_0__1_,
         cell_2026_a_HPC2_and_p_0_out_1__0_,
         cell_2026_a_HPC2_and_p_1_out_0__1_,
         cell_2026_a_HPC2_and_p_1_out_1__0_,
         cell_2026_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2026_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2026_a_HPC2_and_p_1_in_0__1_, cell_2026_a_HPC2_and_p_1_in_1__0_,
         cell_2026_a_HPC2_and_s_out_0__1_, cell_2026_a_HPC2_and_s_out_1__0_,
         cell_2026_a_HPC2_and_p_0_in_0__1_, cell_2026_a_HPC2_and_p_0_in_1__0_,
         cell_2026_a_HPC2_and_s_in_0__1_, cell_2026_a_HPC2_and_s_in_1__0_,
         cell_2026_a_HPC2_and_z_0__0_, cell_2026_a_HPC2_and_z_1__1_,
         cell_2027_a_HPC2_and_n9, cell_2027_a_HPC2_and_n8,
         cell_2027_a_HPC2_and_n7, cell_2027_a_HPC2_and_p_0_out_0__1_,
         cell_2027_a_HPC2_and_p_0_out_1__0_,
         cell_2027_a_HPC2_and_p_1_out_0__1_,
         cell_2027_a_HPC2_and_p_1_out_1__0_,
         cell_2027_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2027_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2027_a_HPC2_and_p_1_in_0__1_, cell_2027_a_HPC2_and_p_1_in_1__0_,
         cell_2027_a_HPC2_and_s_out_0__1_, cell_2027_a_HPC2_and_s_out_1__0_,
         cell_2027_a_HPC2_and_p_0_in_0__1_, cell_2027_a_HPC2_and_p_0_in_1__0_,
         cell_2027_a_HPC2_and_s_in_0__1_, cell_2027_a_HPC2_and_s_in_1__0_,
         cell_2027_a_HPC2_and_z_0__0_, cell_2027_a_HPC2_and_z_1__1_,
         cell_2028_a_HPC2_and_n9, cell_2028_a_HPC2_and_n8,
         cell_2028_a_HPC2_and_n7, cell_2028_a_HPC2_and_p_0_out_0__1_,
         cell_2028_a_HPC2_and_p_0_out_1__0_,
         cell_2028_a_HPC2_and_p_1_out_0__1_,
         cell_2028_a_HPC2_and_p_1_out_1__0_,
         cell_2028_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2028_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2028_a_HPC2_and_p_1_in_0__1_, cell_2028_a_HPC2_and_p_1_in_1__0_,
         cell_2028_a_HPC2_and_s_out_0__1_, cell_2028_a_HPC2_and_s_out_1__0_,
         cell_2028_a_HPC2_and_p_0_in_0__1_, cell_2028_a_HPC2_and_p_0_in_1__0_,
         cell_2028_a_HPC2_and_s_in_0__1_, cell_2028_a_HPC2_and_s_in_1__0_,
         cell_2028_a_HPC2_and_z_0__0_, cell_2028_a_HPC2_and_z_1__1_,
         cell_2029_a_HPC2_and_n9, cell_2029_a_HPC2_and_n8,
         cell_2029_a_HPC2_and_n7, cell_2029_a_HPC2_and_p_0_out_0__1_,
         cell_2029_a_HPC2_and_p_0_out_1__0_,
         cell_2029_a_HPC2_and_p_1_out_0__1_,
         cell_2029_a_HPC2_and_p_1_out_1__0_,
         cell_2029_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2029_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2029_a_HPC2_and_p_1_in_0__1_, cell_2029_a_HPC2_and_p_1_in_1__0_,
         cell_2029_a_HPC2_and_s_out_0__1_, cell_2029_a_HPC2_and_s_out_1__0_,
         cell_2029_a_HPC2_and_p_0_in_0__1_, cell_2029_a_HPC2_and_p_0_in_1__0_,
         cell_2029_a_HPC2_and_s_in_0__1_, cell_2029_a_HPC2_and_s_in_1__0_,
         cell_2029_a_HPC2_and_z_0__0_, cell_2029_a_HPC2_and_z_1__1_,
         cell_2030_a_HPC2_and_n9, cell_2030_a_HPC2_and_n8,
         cell_2030_a_HPC2_and_n7, cell_2030_a_HPC2_and_p_0_out_0__1_,
         cell_2030_a_HPC2_and_p_0_out_1__0_,
         cell_2030_a_HPC2_and_p_1_out_0__1_,
         cell_2030_a_HPC2_and_p_1_out_1__0_,
         cell_2030_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2030_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2030_a_HPC2_and_p_1_in_0__1_, cell_2030_a_HPC2_and_p_1_in_1__0_,
         cell_2030_a_HPC2_and_s_out_0__1_, cell_2030_a_HPC2_and_s_out_1__0_,
         cell_2030_a_HPC2_and_p_0_in_0__1_, cell_2030_a_HPC2_and_p_0_in_1__0_,
         cell_2030_a_HPC2_and_s_in_0__1_, cell_2030_a_HPC2_and_s_in_1__0_,
         cell_2030_a_HPC2_and_z_0__0_, cell_2030_a_HPC2_and_z_1__1_,
         cell_2031_a_HPC2_and_n9, cell_2031_a_HPC2_and_n8,
         cell_2031_a_HPC2_and_n7, cell_2031_a_HPC2_and_p_0_out_0__1_,
         cell_2031_a_HPC2_and_p_0_out_1__0_,
         cell_2031_a_HPC2_and_p_1_out_0__1_,
         cell_2031_a_HPC2_and_p_1_out_1__0_,
         cell_2031_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2031_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2031_a_HPC2_and_p_1_in_0__1_, cell_2031_a_HPC2_and_p_1_in_1__0_,
         cell_2031_a_HPC2_and_s_out_0__1_, cell_2031_a_HPC2_and_s_out_1__0_,
         cell_2031_a_HPC2_and_p_0_in_0__1_, cell_2031_a_HPC2_and_p_0_in_1__0_,
         cell_2031_a_HPC2_and_s_in_0__1_, cell_2031_a_HPC2_and_s_in_1__0_,
         cell_2031_a_HPC2_and_z_0__0_, cell_2031_a_HPC2_and_z_1__1_,
         cell_2032_a_HPC2_and_n9, cell_2032_a_HPC2_and_n8,
         cell_2032_a_HPC2_and_n7, cell_2032_a_HPC2_and_p_0_out_0__1_,
         cell_2032_a_HPC2_and_p_0_out_1__0_,
         cell_2032_a_HPC2_and_p_1_out_0__1_,
         cell_2032_a_HPC2_and_p_1_out_1__0_,
         cell_2032_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2032_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2032_a_HPC2_and_p_1_in_0__1_, cell_2032_a_HPC2_and_p_1_in_1__0_,
         cell_2032_a_HPC2_and_s_out_0__1_, cell_2032_a_HPC2_and_s_out_1__0_,
         cell_2032_a_HPC2_and_p_0_in_0__1_, cell_2032_a_HPC2_and_p_0_in_1__0_,
         cell_2032_a_HPC2_and_s_in_0__1_, cell_2032_a_HPC2_and_s_in_1__0_,
         cell_2032_a_HPC2_and_z_0__0_, cell_2032_a_HPC2_and_z_1__1_,
         cell_2033_a_HPC2_and_n9, cell_2033_a_HPC2_and_n8,
         cell_2033_a_HPC2_and_n7, cell_2033_a_HPC2_and_p_0_out_0__1_,
         cell_2033_a_HPC2_and_p_0_out_1__0_,
         cell_2033_a_HPC2_and_p_1_out_0__1_,
         cell_2033_a_HPC2_and_p_1_out_1__0_,
         cell_2033_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2033_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2033_a_HPC2_and_p_1_in_0__1_, cell_2033_a_HPC2_and_p_1_in_1__0_,
         cell_2033_a_HPC2_and_s_out_0__1_, cell_2033_a_HPC2_and_s_out_1__0_,
         cell_2033_a_HPC2_and_p_0_in_0__1_, cell_2033_a_HPC2_and_p_0_in_1__0_,
         cell_2033_a_HPC2_and_s_in_0__1_, cell_2033_a_HPC2_and_s_in_1__0_,
         cell_2033_a_HPC2_and_z_0__0_, cell_2033_a_HPC2_and_z_1__1_,
         cell_2034_a_HPC2_and_n9, cell_2034_a_HPC2_and_n8,
         cell_2034_a_HPC2_and_n7, cell_2034_a_HPC2_and_p_0_out_0__1_,
         cell_2034_a_HPC2_and_p_0_out_1__0_,
         cell_2034_a_HPC2_and_p_1_out_0__1_,
         cell_2034_a_HPC2_and_p_1_out_1__0_,
         cell_2034_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2034_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2034_a_HPC2_and_p_1_in_0__1_, cell_2034_a_HPC2_and_p_1_in_1__0_,
         cell_2034_a_HPC2_and_s_out_0__1_, cell_2034_a_HPC2_and_s_out_1__0_,
         cell_2034_a_HPC2_and_p_0_in_0__1_, cell_2034_a_HPC2_and_p_0_in_1__0_,
         cell_2034_a_HPC2_and_s_in_0__1_, cell_2034_a_HPC2_and_s_in_1__0_,
         cell_2034_a_HPC2_and_z_0__0_, cell_2034_a_HPC2_and_z_1__1_,
         cell_2035_a_HPC2_and_n9, cell_2035_a_HPC2_and_n8,
         cell_2035_a_HPC2_and_n7, cell_2035_a_HPC2_and_p_0_out_0__1_,
         cell_2035_a_HPC2_and_p_0_out_1__0_,
         cell_2035_a_HPC2_and_p_1_out_0__1_,
         cell_2035_a_HPC2_and_p_1_out_1__0_,
         cell_2035_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2035_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2035_a_HPC2_and_p_1_in_0__1_, cell_2035_a_HPC2_and_p_1_in_1__0_,
         cell_2035_a_HPC2_and_s_out_0__1_, cell_2035_a_HPC2_and_s_out_1__0_,
         cell_2035_a_HPC2_and_p_0_in_0__1_, cell_2035_a_HPC2_and_p_0_in_1__0_,
         cell_2035_a_HPC2_and_s_in_0__1_, cell_2035_a_HPC2_and_s_in_1__0_,
         cell_2035_a_HPC2_and_z_0__0_, cell_2035_a_HPC2_and_z_1__1_,
         cell_2036_a_HPC2_and_n9, cell_2036_a_HPC2_and_n8,
         cell_2036_a_HPC2_and_n7, cell_2036_a_HPC2_and_p_0_out_0__1_,
         cell_2036_a_HPC2_and_p_0_out_1__0_,
         cell_2036_a_HPC2_and_p_1_out_0__1_,
         cell_2036_a_HPC2_and_p_1_out_1__0_,
         cell_2036_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2036_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2036_a_HPC2_and_p_1_in_0__1_, cell_2036_a_HPC2_and_p_1_in_1__0_,
         cell_2036_a_HPC2_and_s_out_0__1_, cell_2036_a_HPC2_and_s_out_1__0_,
         cell_2036_a_HPC2_and_p_0_in_0__1_, cell_2036_a_HPC2_and_p_0_in_1__0_,
         cell_2036_a_HPC2_and_s_in_0__1_, cell_2036_a_HPC2_and_s_in_1__0_,
         cell_2036_a_HPC2_and_z_0__0_, cell_2036_a_HPC2_and_z_1__1_,
         cell_2037_a_HPC2_and_n9, cell_2037_a_HPC2_and_n8,
         cell_2037_a_HPC2_and_n7, cell_2037_a_HPC2_and_p_0_out_0__1_,
         cell_2037_a_HPC2_and_p_0_out_1__0_,
         cell_2037_a_HPC2_and_p_1_out_0__1_,
         cell_2037_a_HPC2_and_p_1_out_1__0_,
         cell_2037_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2037_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2037_a_HPC2_and_p_1_in_0__1_, cell_2037_a_HPC2_and_p_1_in_1__0_,
         cell_2037_a_HPC2_and_s_out_0__1_, cell_2037_a_HPC2_and_s_out_1__0_,
         cell_2037_a_HPC2_and_p_0_in_0__1_, cell_2037_a_HPC2_and_p_0_in_1__0_,
         cell_2037_a_HPC2_and_s_in_0__1_, cell_2037_a_HPC2_and_s_in_1__0_,
         cell_2037_a_HPC2_and_z_0__0_, cell_2037_a_HPC2_and_z_1__1_,
         cell_2038_a_HPC2_and_n9, cell_2038_a_HPC2_and_n8,
         cell_2038_a_HPC2_and_n7, cell_2038_a_HPC2_and_p_0_out_0__1_,
         cell_2038_a_HPC2_and_p_0_out_1__0_,
         cell_2038_a_HPC2_and_p_1_out_0__1_,
         cell_2038_a_HPC2_and_p_1_out_1__0_,
         cell_2038_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2038_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2038_a_HPC2_and_p_1_in_0__1_, cell_2038_a_HPC2_and_p_1_in_1__0_,
         cell_2038_a_HPC2_and_s_out_0__1_, cell_2038_a_HPC2_and_s_out_1__0_,
         cell_2038_a_HPC2_and_p_0_in_0__1_, cell_2038_a_HPC2_and_p_0_in_1__0_,
         cell_2038_a_HPC2_and_s_in_0__1_, cell_2038_a_HPC2_and_s_in_1__0_,
         cell_2038_a_HPC2_and_z_0__0_, cell_2038_a_HPC2_and_z_1__1_,
         cell_2039_a_HPC2_and_n9, cell_2039_a_HPC2_and_n8,
         cell_2039_a_HPC2_and_n7, cell_2039_a_HPC2_and_p_0_out_0__1_,
         cell_2039_a_HPC2_and_p_0_out_1__0_,
         cell_2039_a_HPC2_and_p_1_out_0__1_,
         cell_2039_a_HPC2_and_p_1_out_1__0_,
         cell_2039_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2039_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2039_a_HPC2_and_p_1_in_0__1_, cell_2039_a_HPC2_and_p_1_in_1__0_,
         cell_2039_a_HPC2_and_s_out_0__1_, cell_2039_a_HPC2_and_s_out_1__0_,
         cell_2039_a_HPC2_and_p_0_in_0__1_, cell_2039_a_HPC2_and_p_0_in_1__0_,
         cell_2039_a_HPC2_and_s_in_0__1_, cell_2039_a_HPC2_and_s_in_1__0_,
         cell_2039_a_HPC2_and_z_0__0_, cell_2039_a_HPC2_and_z_1__1_,
         cell_2040_a_HPC2_and_n9, cell_2040_a_HPC2_and_n8,
         cell_2040_a_HPC2_and_n7, cell_2040_a_HPC2_and_p_0_out_0__1_,
         cell_2040_a_HPC2_and_p_0_out_1__0_,
         cell_2040_a_HPC2_and_p_1_out_0__1_,
         cell_2040_a_HPC2_and_p_1_out_1__0_,
         cell_2040_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2040_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2040_a_HPC2_and_p_1_in_0__1_, cell_2040_a_HPC2_and_p_1_in_1__0_,
         cell_2040_a_HPC2_and_s_out_0__1_, cell_2040_a_HPC2_and_s_out_1__0_,
         cell_2040_a_HPC2_and_p_0_in_0__1_, cell_2040_a_HPC2_and_p_0_in_1__0_,
         cell_2040_a_HPC2_and_s_in_0__1_, cell_2040_a_HPC2_and_s_in_1__0_,
         cell_2040_a_HPC2_and_z_0__0_, cell_2040_a_HPC2_and_z_1__1_,
         cell_2041_a_HPC2_and_n9, cell_2041_a_HPC2_and_n8,
         cell_2041_a_HPC2_and_n7, cell_2041_a_HPC2_and_p_0_out_0__1_,
         cell_2041_a_HPC2_and_p_0_out_1__0_,
         cell_2041_a_HPC2_and_p_1_out_0__1_,
         cell_2041_a_HPC2_and_p_1_out_1__0_,
         cell_2041_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2041_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2041_a_HPC2_and_p_1_in_0__1_, cell_2041_a_HPC2_and_p_1_in_1__0_,
         cell_2041_a_HPC2_and_s_out_0__1_, cell_2041_a_HPC2_and_s_out_1__0_,
         cell_2041_a_HPC2_and_p_0_in_0__1_, cell_2041_a_HPC2_and_p_0_in_1__0_,
         cell_2041_a_HPC2_and_s_in_0__1_, cell_2041_a_HPC2_and_s_in_1__0_,
         cell_2041_a_HPC2_and_z_0__0_, cell_2041_a_HPC2_and_z_1__1_,
         cell_2042_a_HPC2_and_n9, cell_2042_a_HPC2_and_n8,
         cell_2042_a_HPC2_and_n7, cell_2042_a_HPC2_and_p_0_out_0__1_,
         cell_2042_a_HPC2_and_p_0_out_1__0_,
         cell_2042_a_HPC2_and_p_1_out_0__1_,
         cell_2042_a_HPC2_and_p_1_out_1__0_,
         cell_2042_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2042_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2042_a_HPC2_and_p_1_in_0__1_, cell_2042_a_HPC2_and_p_1_in_1__0_,
         cell_2042_a_HPC2_and_s_out_0__1_, cell_2042_a_HPC2_and_s_out_1__0_,
         cell_2042_a_HPC2_and_p_0_in_0__1_, cell_2042_a_HPC2_and_p_0_in_1__0_,
         cell_2042_a_HPC2_and_s_in_0__1_, cell_2042_a_HPC2_and_s_in_1__0_,
         cell_2042_a_HPC2_and_z_0__0_, cell_2042_a_HPC2_and_z_1__1_,
         cell_2043_a_HPC2_and_n9, cell_2043_a_HPC2_and_n8,
         cell_2043_a_HPC2_and_n7, cell_2043_a_HPC2_and_p_0_out_0__1_,
         cell_2043_a_HPC2_and_p_0_out_1__0_,
         cell_2043_a_HPC2_and_p_1_out_0__1_,
         cell_2043_a_HPC2_and_p_1_out_1__0_,
         cell_2043_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2043_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2043_a_HPC2_and_p_1_in_0__1_, cell_2043_a_HPC2_and_p_1_in_1__0_,
         cell_2043_a_HPC2_and_s_out_0__1_, cell_2043_a_HPC2_and_s_out_1__0_,
         cell_2043_a_HPC2_and_p_0_in_0__1_, cell_2043_a_HPC2_and_p_0_in_1__0_,
         cell_2043_a_HPC2_and_s_in_0__1_, cell_2043_a_HPC2_and_s_in_1__0_,
         cell_2043_a_HPC2_and_z_0__0_, cell_2043_a_HPC2_and_z_1__1_,
         cell_2044_a_HPC2_and_n9, cell_2044_a_HPC2_and_n8,
         cell_2044_a_HPC2_and_n7, cell_2044_a_HPC2_and_p_0_out_0__1_,
         cell_2044_a_HPC2_and_p_0_out_1__0_,
         cell_2044_a_HPC2_and_p_1_out_0__1_,
         cell_2044_a_HPC2_and_p_1_out_1__0_,
         cell_2044_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2044_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2044_a_HPC2_and_p_1_in_0__1_, cell_2044_a_HPC2_and_p_1_in_1__0_,
         cell_2044_a_HPC2_and_s_out_0__1_, cell_2044_a_HPC2_and_s_out_1__0_,
         cell_2044_a_HPC2_and_p_0_in_0__1_, cell_2044_a_HPC2_and_p_0_in_1__0_,
         cell_2044_a_HPC2_and_s_in_0__1_, cell_2044_a_HPC2_and_s_in_1__0_,
         cell_2044_a_HPC2_and_z_0__0_, cell_2044_a_HPC2_and_z_1__1_,
         cell_2045_a_HPC2_and_n9, cell_2045_a_HPC2_and_n8,
         cell_2045_a_HPC2_and_n7, cell_2045_a_HPC2_and_p_0_out_0__1_,
         cell_2045_a_HPC2_and_p_0_out_1__0_,
         cell_2045_a_HPC2_and_p_1_out_0__1_,
         cell_2045_a_HPC2_and_p_1_out_1__0_,
         cell_2045_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2045_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2045_a_HPC2_and_p_1_in_0__1_, cell_2045_a_HPC2_and_p_1_in_1__0_,
         cell_2045_a_HPC2_and_s_out_0__1_, cell_2045_a_HPC2_and_s_out_1__0_,
         cell_2045_a_HPC2_and_p_0_in_0__1_, cell_2045_a_HPC2_and_p_0_in_1__0_,
         cell_2045_a_HPC2_and_s_in_0__1_, cell_2045_a_HPC2_and_s_in_1__0_,
         cell_2045_a_HPC2_and_z_0__0_, cell_2045_a_HPC2_and_z_1__1_,
         cell_2046_a_HPC2_and_n9, cell_2046_a_HPC2_and_n8,
         cell_2046_a_HPC2_and_n7, cell_2046_a_HPC2_and_p_0_out_0__1_,
         cell_2046_a_HPC2_and_p_0_out_1__0_,
         cell_2046_a_HPC2_and_p_1_out_0__1_,
         cell_2046_a_HPC2_and_p_1_out_1__0_,
         cell_2046_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2046_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2046_a_HPC2_and_p_1_in_0__1_, cell_2046_a_HPC2_and_p_1_in_1__0_,
         cell_2046_a_HPC2_and_s_out_0__1_, cell_2046_a_HPC2_and_s_out_1__0_,
         cell_2046_a_HPC2_and_p_0_in_0__1_, cell_2046_a_HPC2_and_p_0_in_1__0_,
         cell_2046_a_HPC2_and_s_in_0__1_, cell_2046_a_HPC2_and_s_in_1__0_,
         cell_2046_a_HPC2_and_z_0__0_, cell_2046_a_HPC2_and_z_1__1_,
         cell_2047_a_HPC2_and_n9, cell_2047_a_HPC2_and_n8,
         cell_2047_a_HPC2_and_n7, cell_2047_a_HPC2_and_p_0_out_0__1_,
         cell_2047_a_HPC2_and_p_0_out_1__0_,
         cell_2047_a_HPC2_and_p_1_out_0__1_,
         cell_2047_a_HPC2_and_p_1_out_1__0_,
         cell_2047_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2047_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2047_a_HPC2_and_p_1_in_0__1_, cell_2047_a_HPC2_and_p_1_in_1__0_,
         cell_2047_a_HPC2_and_s_out_0__1_, cell_2047_a_HPC2_and_s_out_1__0_,
         cell_2047_a_HPC2_and_p_0_in_0__1_, cell_2047_a_HPC2_and_p_0_in_1__0_,
         cell_2047_a_HPC2_and_s_in_0__1_, cell_2047_a_HPC2_and_s_in_1__0_,
         cell_2047_a_HPC2_and_z_0__0_, cell_2047_a_HPC2_and_z_1__1_,
         cell_2048_a_HPC2_and_n9, cell_2048_a_HPC2_and_n8,
         cell_2048_a_HPC2_and_n7, cell_2048_a_HPC2_and_p_0_out_0__1_,
         cell_2048_a_HPC2_and_p_0_out_1__0_,
         cell_2048_a_HPC2_and_p_1_out_0__1_,
         cell_2048_a_HPC2_and_p_1_out_1__0_,
         cell_2048_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2048_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2048_a_HPC2_and_p_1_in_0__1_, cell_2048_a_HPC2_and_p_1_in_1__0_,
         cell_2048_a_HPC2_and_s_out_0__1_, cell_2048_a_HPC2_and_s_out_1__0_,
         cell_2048_a_HPC2_and_p_0_in_0__1_, cell_2048_a_HPC2_and_p_0_in_1__0_,
         cell_2048_a_HPC2_and_s_in_0__1_, cell_2048_a_HPC2_and_s_in_1__0_,
         cell_2048_a_HPC2_and_z_0__0_, cell_2048_a_HPC2_and_z_1__1_,
         cell_2049_a_HPC2_and_n9, cell_2049_a_HPC2_and_n8,
         cell_2049_a_HPC2_and_n7, cell_2049_a_HPC2_and_p_0_out_0__1_,
         cell_2049_a_HPC2_and_p_0_out_1__0_,
         cell_2049_a_HPC2_and_p_1_out_0__1_,
         cell_2049_a_HPC2_and_p_1_out_1__0_,
         cell_2049_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2049_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2049_a_HPC2_and_p_1_in_0__1_, cell_2049_a_HPC2_and_p_1_in_1__0_,
         cell_2049_a_HPC2_and_s_out_0__1_, cell_2049_a_HPC2_and_s_out_1__0_,
         cell_2049_a_HPC2_and_p_0_in_0__1_, cell_2049_a_HPC2_and_p_0_in_1__0_,
         cell_2049_a_HPC2_and_s_in_0__1_, cell_2049_a_HPC2_and_s_in_1__0_,
         cell_2049_a_HPC2_and_z_0__0_, cell_2049_a_HPC2_and_z_1__1_,
         cell_2050_a_HPC2_and_n9, cell_2050_a_HPC2_and_n8,
         cell_2050_a_HPC2_and_n7, cell_2050_a_HPC2_and_p_0_out_0__1_,
         cell_2050_a_HPC2_and_p_0_out_1__0_,
         cell_2050_a_HPC2_and_p_1_out_0__1_,
         cell_2050_a_HPC2_and_p_1_out_1__0_,
         cell_2050_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2050_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2050_a_HPC2_and_p_1_in_0__1_, cell_2050_a_HPC2_and_p_1_in_1__0_,
         cell_2050_a_HPC2_and_s_out_0__1_, cell_2050_a_HPC2_and_s_out_1__0_,
         cell_2050_a_HPC2_and_p_0_in_0__1_, cell_2050_a_HPC2_and_p_0_in_1__0_,
         cell_2050_a_HPC2_and_s_in_0__1_, cell_2050_a_HPC2_and_s_in_1__0_,
         cell_2050_a_HPC2_and_z_0__0_, cell_2050_a_HPC2_and_z_1__1_,
         cell_2051_a_HPC2_and_n9, cell_2051_a_HPC2_and_n8,
         cell_2051_a_HPC2_and_n7, cell_2051_a_HPC2_and_p_0_out_0__1_,
         cell_2051_a_HPC2_and_p_0_out_1__0_,
         cell_2051_a_HPC2_and_p_1_out_0__1_,
         cell_2051_a_HPC2_and_p_1_out_1__0_,
         cell_2051_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2051_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2051_a_HPC2_and_p_1_in_0__1_, cell_2051_a_HPC2_and_p_1_in_1__0_,
         cell_2051_a_HPC2_and_s_out_0__1_, cell_2051_a_HPC2_and_s_out_1__0_,
         cell_2051_a_HPC2_and_p_0_in_0__1_, cell_2051_a_HPC2_and_p_0_in_1__0_,
         cell_2051_a_HPC2_and_s_in_0__1_, cell_2051_a_HPC2_and_s_in_1__0_,
         cell_2051_a_HPC2_and_z_0__0_, cell_2051_a_HPC2_and_z_1__1_,
         cell_2052_a_HPC2_and_n9, cell_2052_a_HPC2_and_n8,
         cell_2052_a_HPC2_and_n7, cell_2052_a_HPC2_and_p_0_out_0__1_,
         cell_2052_a_HPC2_and_p_0_out_1__0_,
         cell_2052_a_HPC2_and_p_1_out_0__1_,
         cell_2052_a_HPC2_and_p_1_out_1__0_,
         cell_2052_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2052_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2052_a_HPC2_and_p_1_in_0__1_, cell_2052_a_HPC2_and_p_1_in_1__0_,
         cell_2052_a_HPC2_and_s_out_0__1_, cell_2052_a_HPC2_and_s_out_1__0_,
         cell_2052_a_HPC2_and_p_0_in_0__1_, cell_2052_a_HPC2_and_p_0_in_1__0_,
         cell_2052_a_HPC2_and_s_in_0__1_, cell_2052_a_HPC2_and_s_in_1__0_,
         cell_2052_a_HPC2_and_z_0__0_, cell_2052_a_HPC2_and_z_1__1_,
         cell_2053_a_HPC2_and_n9, cell_2053_a_HPC2_and_n8,
         cell_2053_a_HPC2_and_n7, cell_2053_a_HPC2_and_p_0_out_0__1_,
         cell_2053_a_HPC2_and_p_0_out_1__0_,
         cell_2053_a_HPC2_and_p_1_out_0__1_,
         cell_2053_a_HPC2_and_p_1_out_1__0_,
         cell_2053_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2053_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2053_a_HPC2_and_p_1_in_0__1_, cell_2053_a_HPC2_and_p_1_in_1__0_,
         cell_2053_a_HPC2_and_s_out_0__1_, cell_2053_a_HPC2_and_s_out_1__0_,
         cell_2053_a_HPC2_and_p_0_in_0__1_, cell_2053_a_HPC2_and_p_0_in_1__0_,
         cell_2053_a_HPC2_and_s_in_0__1_, cell_2053_a_HPC2_and_s_in_1__0_,
         cell_2053_a_HPC2_and_z_0__0_, cell_2053_a_HPC2_and_z_1__1_,
         cell_2054_a_HPC2_and_n9, cell_2054_a_HPC2_and_n8,
         cell_2054_a_HPC2_and_n7, cell_2054_a_HPC2_and_p_0_out_0__1_,
         cell_2054_a_HPC2_and_p_0_out_1__0_,
         cell_2054_a_HPC2_and_p_1_out_0__1_,
         cell_2054_a_HPC2_and_p_1_out_1__0_,
         cell_2054_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2054_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2054_a_HPC2_and_p_1_in_0__1_, cell_2054_a_HPC2_and_p_1_in_1__0_,
         cell_2054_a_HPC2_and_s_out_0__1_, cell_2054_a_HPC2_and_s_out_1__0_,
         cell_2054_a_HPC2_and_p_0_in_0__1_, cell_2054_a_HPC2_and_p_0_in_1__0_,
         cell_2054_a_HPC2_and_s_in_0__1_, cell_2054_a_HPC2_and_s_in_1__0_,
         cell_2054_a_HPC2_and_z_0__0_, cell_2054_a_HPC2_and_z_1__1_,
         cell_2055_a_HPC2_and_n9, cell_2055_a_HPC2_and_n8,
         cell_2055_a_HPC2_and_n7, cell_2055_a_HPC2_and_p_0_out_0__1_,
         cell_2055_a_HPC2_and_p_0_out_1__0_,
         cell_2055_a_HPC2_and_p_1_out_0__1_,
         cell_2055_a_HPC2_and_p_1_out_1__0_,
         cell_2055_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2055_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2055_a_HPC2_and_p_1_in_0__1_, cell_2055_a_HPC2_and_p_1_in_1__0_,
         cell_2055_a_HPC2_and_s_out_0__1_, cell_2055_a_HPC2_and_s_out_1__0_,
         cell_2055_a_HPC2_and_p_0_in_0__1_, cell_2055_a_HPC2_and_p_0_in_1__0_,
         cell_2055_a_HPC2_and_s_in_0__1_, cell_2055_a_HPC2_and_s_in_1__0_,
         cell_2055_a_HPC2_and_z_0__0_, cell_2055_a_HPC2_and_z_1__1_,
         cell_2056_a_HPC2_and_n9, cell_2056_a_HPC2_and_n8,
         cell_2056_a_HPC2_and_n7, cell_2056_a_HPC2_and_p_0_out_0__1_,
         cell_2056_a_HPC2_and_p_0_out_1__0_,
         cell_2056_a_HPC2_and_p_1_out_0__1_,
         cell_2056_a_HPC2_and_p_1_out_1__0_,
         cell_2056_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2056_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2056_a_HPC2_and_p_1_in_0__1_, cell_2056_a_HPC2_and_p_1_in_1__0_,
         cell_2056_a_HPC2_and_s_out_0__1_, cell_2056_a_HPC2_and_s_out_1__0_,
         cell_2056_a_HPC2_and_p_0_in_0__1_, cell_2056_a_HPC2_and_p_0_in_1__0_,
         cell_2056_a_HPC2_and_s_in_0__1_, cell_2056_a_HPC2_and_s_in_1__0_,
         cell_2056_a_HPC2_and_z_0__0_, cell_2056_a_HPC2_and_z_1__1_,
         cell_2057_a_HPC2_and_n9, cell_2057_a_HPC2_and_n8,
         cell_2057_a_HPC2_and_n7, cell_2057_a_HPC2_and_p_0_out_0__1_,
         cell_2057_a_HPC2_and_p_0_out_1__0_,
         cell_2057_a_HPC2_and_p_1_out_0__1_,
         cell_2057_a_HPC2_and_p_1_out_1__0_,
         cell_2057_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2057_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2057_a_HPC2_and_p_1_in_0__1_, cell_2057_a_HPC2_and_p_1_in_1__0_,
         cell_2057_a_HPC2_and_s_out_0__1_, cell_2057_a_HPC2_and_s_out_1__0_,
         cell_2057_a_HPC2_and_p_0_in_0__1_, cell_2057_a_HPC2_and_p_0_in_1__0_,
         cell_2057_a_HPC2_and_s_in_0__1_, cell_2057_a_HPC2_and_s_in_1__0_,
         cell_2057_a_HPC2_and_z_0__0_, cell_2057_a_HPC2_and_z_1__1_,
         cell_2058_a_HPC2_and_n9, cell_2058_a_HPC2_and_n8,
         cell_2058_a_HPC2_and_n7, cell_2058_a_HPC2_and_p_0_out_0__1_,
         cell_2058_a_HPC2_and_p_0_out_1__0_,
         cell_2058_a_HPC2_and_p_1_out_0__1_,
         cell_2058_a_HPC2_and_p_1_out_1__0_,
         cell_2058_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2058_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2058_a_HPC2_and_p_1_in_0__1_, cell_2058_a_HPC2_and_p_1_in_1__0_,
         cell_2058_a_HPC2_and_s_out_0__1_, cell_2058_a_HPC2_and_s_out_1__0_,
         cell_2058_a_HPC2_and_p_0_in_0__1_, cell_2058_a_HPC2_and_p_0_in_1__0_,
         cell_2058_a_HPC2_and_s_in_0__1_, cell_2058_a_HPC2_and_s_in_1__0_,
         cell_2058_a_HPC2_and_z_0__0_, cell_2058_a_HPC2_and_z_1__1_,
         cell_2059_a_HPC2_and_n9, cell_2059_a_HPC2_and_n8,
         cell_2059_a_HPC2_and_n7, cell_2059_a_HPC2_and_p_0_out_0__1_,
         cell_2059_a_HPC2_and_p_0_out_1__0_,
         cell_2059_a_HPC2_and_p_1_out_0__1_,
         cell_2059_a_HPC2_and_p_1_out_1__0_,
         cell_2059_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2059_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2059_a_HPC2_and_p_1_in_0__1_, cell_2059_a_HPC2_and_p_1_in_1__0_,
         cell_2059_a_HPC2_and_s_out_0__1_, cell_2059_a_HPC2_and_s_out_1__0_,
         cell_2059_a_HPC2_and_p_0_in_0__1_, cell_2059_a_HPC2_and_p_0_in_1__0_,
         cell_2059_a_HPC2_and_s_in_0__1_, cell_2059_a_HPC2_and_s_in_1__0_,
         cell_2059_a_HPC2_and_z_0__0_, cell_2059_a_HPC2_and_z_1__1_,
         cell_2060_a_HPC2_and_n9, cell_2060_a_HPC2_and_n8,
         cell_2060_a_HPC2_and_n7, cell_2060_a_HPC2_and_p_0_out_0__1_,
         cell_2060_a_HPC2_and_p_0_out_1__0_,
         cell_2060_a_HPC2_and_p_1_out_0__1_,
         cell_2060_a_HPC2_and_p_1_out_1__0_,
         cell_2060_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2060_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2060_a_HPC2_and_p_1_in_0__1_, cell_2060_a_HPC2_and_p_1_in_1__0_,
         cell_2060_a_HPC2_and_s_out_0__1_, cell_2060_a_HPC2_and_s_out_1__0_,
         cell_2060_a_HPC2_and_p_0_in_0__1_, cell_2060_a_HPC2_and_p_0_in_1__0_,
         cell_2060_a_HPC2_and_s_in_0__1_, cell_2060_a_HPC2_and_s_in_1__0_,
         cell_2060_a_HPC2_and_z_0__0_, cell_2060_a_HPC2_and_z_1__1_,
         cell_2061_a_HPC2_and_n9, cell_2061_a_HPC2_and_n8,
         cell_2061_a_HPC2_and_n7, cell_2061_a_HPC2_and_p_0_out_0__1_,
         cell_2061_a_HPC2_and_p_0_out_1__0_,
         cell_2061_a_HPC2_and_p_1_out_0__1_,
         cell_2061_a_HPC2_and_p_1_out_1__0_,
         cell_2061_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2061_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2061_a_HPC2_and_p_1_in_0__1_, cell_2061_a_HPC2_and_p_1_in_1__0_,
         cell_2061_a_HPC2_and_s_out_0__1_, cell_2061_a_HPC2_and_s_out_1__0_,
         cell_2061_a_HPC2_and_p_0_in_0__1_, cell_2061_a_HPC2_and_p_0_in_1__0_,
         cell_2061_a_HPC2_and_s_in_0__1_, cell_2061_a_HPC2_and_s_in_1__0_,
         cell_2061_a_HPC2_and_z_0__0_, cell_2061_a_HPC2_and_z_1__1_,
         cell_2062_a_HPC2_and_n9, cell_2062_a_HPC2_and_n8,
         cell_2062_a_HPC2_and_n7, cell_2062_a_HPC2_and_p_0_out_0__1_,
         cell_2062_a_HPC2_and_p_0_out_1__0_,
         cell_2062_a_HPC2_and_p_1_out_0__1_,
         cell_2062_a_HPC2_and_p_1_out_1__0_,
         cell_2062_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2062_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2062_a_HPC2_and_p_1_in_0__1_, cell_2062_a_HPC2_and_p_1_in_1__0_,
         cell_2062_a_HPC2_and_s_out_0__1_, cell_2062_a_HPC2_and_s_out_1__0_,
         cell_2062_a_HPC2_and_p_0_in_0__1_, cell_2062_a_HPC2_and_p_0_in_1__0_,
         cell_2062_a_HPC2_and_s_in_0__1_, cell_2062_a_HPC2_and_s_in_1__0_,
         cell_2062_a_HPC2_and_z_0__0_, cell_2062_a_HPC2_and_z_1__1_,
         cell_2063_a_HPC2_and_n9, cell_2063_a_HPC2_and_n8,
         cell_2063_a_HPC2_and_n7, cell_2063_a_HPC2_and_p_0_out_0__1_,
         cell_2063_a_HPC2_and_p_0_out_1__0_,
         cell_2063_a_HPC2_and_p_1_out_0__1_,
         cell_2063_a_HPC2_and_p_1_out_1__0_,
         cell_2063_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2063_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2063_a_HPC2_and_p_1_in_0__1_, cell_2063_a_HPC2_and_p_1_in_1__0_,
         cell_2063_a_HPC2_and_s_out_0__1_, cell_2063_a_HPC2_and_s_out_1__0_,
         cell_2063_a_HPC2_and_p_0_in_0__1_, cell_2063_a_HPC2_and_p_0_in_1__0_,
         cell_2063_a_HPC2_and_s_in_0__1_, cell_2063_a_HPC2_and_s_in_1__0_,
         cell_2063_a_HPC2_and_z_0__0_, cell_2063_a_HPC2_and_z_1__1_,
         cell_2064_a_HPC2_and_n9, cell_2064_a_HPC2_and_n8,
         cell_2064_a_HPC2_and_n7, cell_2064_a_HPC2_and_p_0_out_0__1_,
         cell_2064_a_HPC2_and_p_0_out_1__0_,
         cell_2064_a_HPC2_and_p_1_out_0__1_,
         cell_2064_a_HPC2_and_p_1_out_1__0_,
         cell_2064_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2064_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2064_a_HPC2_and_p_1_in_0__1_, cell_2064_a_HPC2_and_p_1_in_1__0_,
         cell_2064_a_HPC2_and_s_out_0__1_, cell_2064_a_HPC2_and_s_out_1__0_,
         cell_2064_a_HPC2_and_p_0_in_0__1_, cell_2064_a_HPC2_and_p_0_in_1__0_,
         cell_2064_a_HPC2_and_s_in_0__1_, cell_2064_a_HPC2_and_s_in_1__0_,
         cell_2064_a_HPC2_and_z_0__0_, cell_2064_a_HPC2_and_z_1__1_,
         cell_2065_a_HPC2_and_n9, cell_2065_a_HPC2_and_n8,
         cell_2065_a_HPC2_and_n7, cell_2065_a_HPC2_and_p_0_out_0__1_,
         cell_2065_a_HPC2_and_p_0_out_1__0_,
         cell_2065_a_HPC2_and_p_1_out_0__1_,
         cell_2065_a_HPC2_and_p_1_out_1__0_,
         cell_2065_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2065_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2065_a_HPC2_and_p_1_in_0__1_, cell_2065_a_HPC2_and_p_1_in_1__0_,
         cell_2065_a_HPC2_and_s_out_0__1_, cell_2065_a_HPC2_and_s_out_1__0_,
         cell_2065_a_HPC2_and_p_0_in_0__1_, cell_2065_a_HPC2_and_p_0_in_1__0_,
         cell_2065_a_HPC2_and_s_in_0__1_, cell_2065_a_HPC2_and_s_in_1__0_,
         cell_2065_a_HPC2_and_z_0__0_, cell_2065_a_HPC2_and_z_1__1_,
         cell_2066_a_HPC2_and_n9, cell_2066_a_HPC2_and_n8,
         cell_2066_a_HPC2_and_n7, cell_2066_a_HPC2_and_p_0_out_0__1_,
         cell_2066_a_HPC2_and_p_0_out_1__0_,
         cell_2066_a_HPC2_and_p_1_out_0__1_,
         cell_2066_a_HPC2_and_p_1_out_1__0_,
         cell_2066_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2066_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2066_a_HPC2_and_p_1_in_0__1_, cell_2066_a_HPC2_and_p_1_in_1__0_,
         cell_2066_a_HPC2_and_s_out_0__1_, cell_2066_a_HPC2_and_s_out_1__0_,
         cell_2066_a_HPC2_and_p_0_in_0__1_, cell_2066_a_HPC2_and_p_0_in_1__0_,
         cell_2066_a_HPC2_and_s_in_0__1_, cell_2066_a_HPC2_and_s_in_1__0_,
         cell_2066_a_HPC2_and_z_0__0_, cell_2066_a_HPC2_and_z_1__1_,
         cell_2067_a_HPC2_and_n9, cell_2067_a_HPC2_and_n8,
         cell_2067_a_HPC2_and_n7, cell_2067_a_HPC2_and_p_0_out_0__1_,
         cell_2067_a_HPC2_and_p_0_out_1__0_,
         cell_2067_a_HPC2_and_p_1_out_0__1_,
         cell_2067_a_HPC2_and_p_1_out_1__0_,
         cell_2067_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2067_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2067_a_HPC2_and_p_1_in_0__1_, cell_2067_a_HPC2_and_p_1_in_1__0_,
         cell_2067_a_HPC2_and_s_out_0__1_, cell_2067_a_HPC2_and_s_out_1__0_,
         cell_2067_a_HPC2_and_p_0_in_0__1_, cell_2067_a_HPC2_and_p_0_in_1__0_,
         cell_2067_a_HPC2_and_s_in_0__1_, cell_2067_a_HPC2_and_s_in_1__0_,
         cell_2067_a_HPC2_and_z_0__0_, cell_2067_a_HPC2_and_z_1__1_,
         cell_2068_a_HPC2_and_n9, cell_2068_a_HPC2_and_n8,
         cell_2068_a_HPC2_and_n7, cell_2068_a_HPC2_and_p_0_out_0__1_,
         cell_2068_a_HPC2_and_p_0_out_1__0_,
         cell_2068_a_HPC2_and_p_1_out_0__1_,
         cell_2068_a_HPC2_and_p_1_out_1__0_,
         cell_2068_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2068_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2068_a_HPC2_and_p_1_in_0__1_, cell_2068_a_HPC2_and_p_1_in_1__0_,
         cell_2068_a_HPC2_and_s_out_0__1_, cell_2068_a_HPC2_and_s_out_1__0_,
         cell_2068_a_HPC2_and_p_0_in_0__1_, cell_2068_a_HPC2_and_p_0_in_1__0_,
         cell_2068_a_HPC2_and_s_in_0__1_, cell_2068_a_HPC2_and_s_in_1__0_,
         cell_2068_a_HPC2_and_z_0__0_, cell_2068_a_HPC2_and_z_1__1_,
         cell_2069_a_HPC2_and_n9, cell_2069_a_HPC2_and_n8,
         cell_2069_a_HPC2_and_n7, cell_2069_a_HPC2_and_p_0_out_0__1_,
         cell_2069_a_HPC2_and_p_0_out_1__0_,
         cell_2069_a_HPC2_and_p_1_out_0__1_,
         cell_2069_a_HPC2_and_p_1_out_1__0_,
         cell_2069_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2069_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2069_a_HPC2_and_p_1_in_0__1_, cell_2069_a_HPC2_and_p_1_in_1__0_,
         cell_2069_a_HPC2_and_s_out_0__1_, cell_2069_a_HPC2_and_s_out_1__0_,
         cell_2069_a_HPC2_and_p_0_in_0__1_, cell_2069_a_HPC2_and_p_0_in_1__0_,
         cell_2069_a_HPC2_and_s_in_0__1_, cell_2069_a_HPC2_and_s_in_1__0_,
         cell_2069_a_HPC2_and_z_0__0_, cell_2069_a_HPC2_and_z_1__1_,
         cell_2070_a_HPC2_and_n9, cell_2070_a_HPC2_and_n8,
         cell_2070_a_HPC2_and_n7, cell_2070_a_HPC2_and_p_0_out_0__1_,
         cell_2070_a_HPC2_and_p_0_out_1__0_,
         cell_2070_a_HPC2_and_p_1_out_0__1_,
         cell_2070_a_HPC2_and_p_1_out_1__0_,
         cell_2070_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2070_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2070_a_HPC2_and_p_1_in_0__1_, cell_2070_a_HPC2_and_p_1_in_1__0_,
         cell_2070_a_HPC2_and_s_out_0__1_, cell_2070_a_HPC2_and_s_out_1__0_,
         cell_2070_a_HPC2_and_p_0_in_0__1_, cell_2070_a_HPC2_and_p_0_in_1__0_,
         cell_2070_a_HPC2_and_s_in_0__1_, cell_2070_a_HPC2_and_s_in_1__0_,
         cell_2070_a_HPC2_and_z_0__0_, cell_2070_a_HPC2_and_z_1__1_,
         cell_2071_a_HPC2_and_n9, cell_2071_a_HPC2_and_n8,
         cell_2071_a_HPC2_and_n7, cell_2071_a_HPC2_and_p_0_out_0__1_,
         cell_2071_a_HPC2_and_p_0_out_1__0_,
         cell_2071_a_HPC2_and_p_1_out_0__1_,
         cell_2071_a_HPC2_and_p_1_out_1__0_,
         cell_2071_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2071_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2071_a_HPC2_and_p_1_in_0__1_, cell_2071_a_HPC2_and_p_1_in_1__0_,
         cell_2071_a_HPC2_and_s_out_0__1_, cell_2071_a_HPC2_and_s_out_1__0_,
         cell_2071_a_HPC2_and_p_0_in_0__1_, cell_2071_a_HPC2_and_p_0_in_1__0_,
         cell_2071_a_HPC2_and_s_in_0__1_, cell_2071_a_HPC2_and_s_in_1__0_,
         cell_2071_a_HPC2_and_z_0__0_, cell_2071_a_HPC2_and_z_1__1_,
         cell_2072_a_HPC2_and_n9, cell_2072_a_HPC2_and_n8,
         cell_2072_a_HPC2_and_n7, cell_2072_a_HPC2_and_p_0_out_0__1_,
         cell_2072_a_HPC2_and_p_0_out_1__0_,
         cell_2072_a_HPC2_and_p_1_out_0__1_,
         cell_2072_a_HPC2_and_p_1_out_1__0_,
         cell_2072_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2072_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2072_a_HPC2_and_p_1_in_0__1_, cell_2072_a_HPC2_and_p_1_in_1__0_,
         cell_2072_a_HPC2_and_s_out_0__1_, cell_2072_a_HPC2_and_s_out_1__0_,
         cell_2072_a_HPC2_and_p_0_in_0__1_, cell_2072_a_HPC2_and_p_0_in_1__0_,
         cell_2072_a_HPC2_and_s_in_0__1_, cell_2072_a_HPC2_and_s_in_1__0_,
         cell_2072_a_HPC2_and_z_0__0_, cell_2072_a_HPC2_and_z_1__1_,
         cell_2073_a_HPC2_and_n9, cell_2073_a_HPC2_and_n8,
         cell_2073_a_HPC2_and_n7, cell_2073_a_HPC2_and_p_0_out_0__1_,
         cell_2073_a_HPC2_and_p_0_out_1__0_,
         cell_2073_a_HPC2_and_p_1_out_0__1_,
         cell_2073_a_HPC2_and_p_1_out_1__0_,
         cell_2073_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2073_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2073_a_HPC2_and_p_1_in_0__1_, cell_2073_a_HPC2_and_p_1_in_1__0_,
         cell_2073_a_HPC2_and_s_out_0__1_, cell_2073_a_HPC2_and_s_out_1__0_,
         cell_2073_a_HPC2_and_p_0_in_0__1_, cell_2073_a_HPC2_and_p_0_in_1__0_,
         cell_2073_a_HPC2_and_s_in_0__1_, cell_2073_a_HPC2_and_s_in_1__0_,
         cell_2073_a_HPC2_and_z_0__0_, cell_2073_a_HPC2_and_z_1__1_,
         cell_2074_a_HPC2_and_n9, cell_2074_a_HPC2_and_n8,
         cell_2074_a_HPC2_and_n7, cell_2074_a_HPC2_and_p_0_out_0__1_,
         cell_2074_a_HPC2_and_p_0_out_1__0_,
         cell_2074_a_HPC2_and_p_1_out_0__1_,
         cell_2074_a_HPC2_and_p_1_out_1__0_,
         cell_2074_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2074_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2074_a_HPC2_and_p_1_in_0__1_, cell_2074_a_HPC2_and_p_1_in_1__0_,
         cell_2074_a_HPC2_and_s_out_0__1_, cell_2074_a_HPC2_and_s_out_1__0_,
         cell_2074_a_HPC2_and_p_0_in_0__1_, cell_2074_a_HPC2_and_p_0_in_1__0_,
         cell_2074_a_HPC2_and_s_in_0__1_, cell_2074_a_HPC2_and_s_in_1__0_,
         cell_2074_a_HPC2_and_z_0__0_, cell_2074_a_HPC2_and_z_1__1_,
         cell_2075_a_HPC2_and_n9, cell_2075_a_HPC2_and_n8,
         cell_2075_a_HPC2_and_n7, cell_2075_a_HPC2_and_p_0_out_0__1_,
         cell_2075_a_HPC2_and_p_0_out_1__0_,
         cell_2075_a_HPC2_and_p_1_out_0__1_,
         cell_2075_a_HPC2_and_p_1_out_1__0_,
         cell_2075_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2075_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2075_a_HPC2_and_p_1_in_0__1_, cell_2075_a_HPC2_and_p_1_in_1__0_,
         cell_2075_a_HPC2_and_s_out_0__1_, cell_2075_a_HPC2_and_s_out_1__0_,
         cell_2075_a_HPC2_and_p_0_in_0__1_, cell_2075_a_HPC2_and_p_0_in_1__0_,
         cell_2075_a_HPC2_and_s_in_0__1_, cell_2075_a_HPC2_and_s_in_1__0_,
         cell_2075_a_HPC2_and_z_0__0_, cell_2075_a_HPC2_and_z_1__1_,
         cell_2076_a_HPC2_and_n9, cell_2076_a_HPC2_and_n8,
         cell_2076_a_HPC2_and_n7, cell_2076_a_HPC2_and_p_0_out_0__1_,
         cell_2076_a_HPC2_and_p_0_out_1__0_,
         cell_2076_a_HPC2_and_p_1_out_0__1_,
         cell_2076_a_HPC2_and_p_1_out_1__0_,
         cell_2076_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2076_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2076_a_HPC2_and_p_1_in_0__1_, cell_2076_a_HPC2_and_p_1_in_1__0_,
         cell_2076_a_HPC2_and_s_out_0__1_, cell_2076_a_HPC2_and_s_out_1__0_,
         cell_2076_a_HPC2_and_p_0_in_0__1_, cell_2076_a_HPC2_and_p_0_in_1__0_,
         cell_2076_a_HPC2_and_s_in_0__1_, cell_2076_a_HPC2_and_s_in_1__0_,
         cell_2076_a_HPC2_and_z_0__0_, cell_2076_a_HPC2_and_z_1__1_,
         cell_2077_a_HPC2_and_n9, cell_2077_a_HPC2_and_n8,
         cell_2077_a_HPC2_and_n7, cell_2077_a_HPC2_and_p_0_out_0__1_,
         cell_2077_a_HPC2_and_p_0_out_1__0_,
         cell_2077_a_HPC2_and_p_1_out_0__1_,
         cell_2077_a_HPC2_and_p_1_out_1__0_,
         cell_2077_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2077_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2077_a_HPC2_and_p_1_in_0__1_, cell_2077_a_HPC2_and_p_1_in_1__0_,
         cell_2077_a_HPC2_and_s_out_0__1_, cell_2077_a_HPC2_and_s_out_1__0_,
         cell_2077_a_HPC2_and_p_0_in_0__1_, cell_2077_a_HPC2_and_p_0_in_1__0_,
         cell_2077_a_HPC2_and_s_in_0__1_, cell_2077_a_HPC2_and_s_in_1__0_,
         cell_2077_a_HPC2_and_z_0__0_, cell_2077_a_HPC2_and_z_1__1_,
         cell_2078_a_HPC2_and_n9, cell_2078_a_HPC2_and_n8,
         cell_2078_a_HPC2_and_n7, cell_2078_a_HPC2_and_p_0_out_0__1_,
         cell_2078_a_HPC2_and_p_0_out_1__0_,
         cell_2078_a_HPC2_and_p_1_out_0__1_,
         cell_2078_a_HPC2_and_p_1_out_1__0_,
         cell_2078_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2078_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2078_a_HPC2_and_p_1_in_0__1_, cell_2078_a_HPC2_and_p_1_in_1__0_,
         cell_2078_a_HPC2_and_s_out_0__1_, cell_2078_a_HPC2_and_s_out_1__0_,
         cell_2078_a_HPC2_and_p_0_in_0__1_, cell_2078_a_HPC2_and_p_0_in_1__0_,
         cell_2078_a_HPC2_and_s_in_0__1_, cell_2078_a_HPC2_and_s_in_1__0_,
         cell_2078_a_HPC2_and_z_0__0_, cell_2078_a_HPC2_and_z_1__1_,
         cell_2079_a_HPC2_and_n9, cell_2079_a_HPC2_and_n8,
         cell_2079_a_HPC2_and_n7, cell_2079_a_HPC2_and_p_0_out_0__1_,
         cell_2079_a_HPC2_and_p_0_out_1__0_,
         cell_2079_a_HPC2_and_p_1_out_0__1_,
         cell_2079_a_HPC2_and_p_1_out_1__0_,
         cell_2079_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2079_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2079_a_HPC2_and_p_1_in_0__1_, cell_2079_a_HPC2_and_p_1_in_1__0_,
         cell_2079_a_HPC2_and_s_out_0__1_, cell_2079_a_HPC2_and_s_out_1__0_,
         cell_2079_a_HPC2_and_p_0_in_0__1_, cell_2079_a_HPC2_and_p_0_in_1__0_,
         cell_2079_a_HPC2_and_s_in_0__1_, cell_2079_a_HPC2_and_s_in_1__0_,
         cell_2079_a_HPC2_and_z_0__0_, cell_2079_a_HPC2_and_z_1__1_,
         cell_2080_a_HPC2_and_n9, cell_2080_a_HPC2_and_n8,
         cell_2080_a_HPC2_and_n7, cell_2080_a_HPC2_and_p_0_out_0__1_,
         cell_2080_a_HPC2_and_p_0_out_1__0_,
         cell_2080_a_HPC2_and_p_1_out_0__1_,
         cell_2080_a_HPC2_and_p_1_out_1__0_,
         cell_2080_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2080_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2080_a_HPC2_and_p_1_in_0__1_, cell_2080_a_HPC2_and_p_1_in_1__0_,
         cell_2080_a_HPC2_and_s_out_0__1_, cell_2080_a_HPC2_and_s_out_1__0_,
         cell_2080_a_HPC2_and_p_0_in_0__1_, cell_2080_a_HPC2_and_p_0_in_1__0_,
         cell_2080_a_HPC2_and_s_in_0__1_, cell_2080_a_HPC2_and_s_in_1__0_,
         cell_2080_a_HPC2_and_z_0__0_, cell_2080_a_HPC2_and_z_1__1_,
         cell_2081_a_HPC2_and_n9, cell_2081_a_HPC2_and_n8,
         cell_2081_a_HPC2_and_n7, cell_2081_a_HPC2_and_p_0_out_0__1_,
         cell_2081_a_HPC2_and_p_0_out_1__0_,
         cell_2081_a_HPC2_and_p_1_out_0__1_,
         cell_2081_a_HPC2_and_p_1_out_1__0_,
         cell_2081_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2081_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2081_a_HPC2_and_p_1_in_0__1_, cell_2081_a_HPC2_and_p_1_in_1__0_,
         cell_2081_a_HPC2_and_s_out_0__1_, cell_2081_a_HPC2_and_s_out_1__0_,
         cell_2081_a_HPC2_and_p_0_in_0__1_, cell_2081_a_HPC2_and_p_0_in_1__0_,
         cell_2081_a_HPC2_and_s_in_0__1_, cell_2081_a_HPC2_and_s_in_1__0_,
         cell_2081_a_HPC2_and_z_0__0_, cell_2081_a_HPC2_and_z_1__1_,
         cell_2082_a_HPC2_and_n9, cell_2082_a_HPC2_and_n8,
         cell_2082_a_HPC2_and_n7, cell_2082_a_HPC2_and_p_0_out_0__1_,
         cell_2082_a_HPC2_and_p_0_out_1__0_,
         cell_2082_a_HPC2_and_p_1_out_0__1_,
         cell_2082_a_HPC2_and_p_1_out_1__0_,
         cell_2082_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2082_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2082_a_HPC2_and_p_1_in_0__1_, cell_2082_a_HPC2_and_p_1_in_1__0_,
         cell_2082_a_HPC2_and_s_out_0__1_, cell_2082_a_HPC2_and_s_out_1__0_,
         cell_2082_a_HPC2_and_p_0_in_0__1_, cell_2082_a_HPC2_and_p_0_in_1__0_,
         cell_2082_a_HPC2_and_s_in_0__1_, cell_2082_a_HPC2_and_s_in_1__0_,
         cell_2082_a_HPC2_and_z_0__0_, cell_2082_a_HPC2_and_z_1__1_,
         cell_2083_a_HPC2_and_n9, cell_2083_a_HPC2_and_n8,
         cell_2083_a_HPC2_and_n7, cell_2083_a_HPC2_and_p_0_out_0__1_,
         cell_2083_a_HPC2_and_p_0_out_1__0_,
         cell_2083_a_HPC2_and_p_1_out_0__1_,
         cell_2083_a_HPC2_and_p_1_out_1__0_,
         cell_2083_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2083_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2083_a_HPC2_and_p_1_in_0__1_, cell_2083_a_HPC2_and_p_1_in_1__0_,
         cell_2083_a_HPC2_and_s_out_0__1_, cell_2083_a_HPC2_and_s_out_1__0_,
         cell_2083_a_HPC2_and_p_0_in_0__1_, cell_2083_a_HPC2_and_p_0_in_1__0_,
         cell_2083_a_HPC2_and_s_in_0__1_, cell_2083_a_HPC2_and_s_in_1__0_,
         cell_2083_a_HPC2_and_z_0__0_, cell_2083_a_HPC2_and_z_1__1_,
         cell_2084_a_HPC2_and_n9, cell_2084_a_HPC2_and_n8,
         cell_2084_a_HPC2_and_n7, cell_2084_a_HPC2_and_p_0_out_0__1_,
         cell_2084_a_HPC2_and_p_0_out_1__0_,
         cell_2084_a_HPC2_and_p_1_out_0__1_,
         cell_2084_a_HPC2_and_p_1_out_1__0_,
         cell_2084_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2084_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2084_a_HPC2_and_p_1_in_0__1_, cell_2084_a_HPC2_and_p_1_in_1__0_,
         cell_2084_a_HPC2_and_s_out_0__1_, cell_2084_a_HPC2_and_s_out_1__0_,
         cell_2084_a_HPC2_and_p_0_in_0__1_, cell_2084_a_HPC2_and_p_0_in_1__0_,
         cell_2084_a_HPC2_and_s_in_0__1_, cell_2084_a_HPC2_and_s_in_1__0_,
         cell_2084_a_HPC2_and_z_0__0_, cell_2084_a_HPC2_and_z_1__1_,
         cell_2085_a_HPC2_and_n9, cell_2085_a_HPC2_and_n8,
         cell_2085_a_HPC2_and_n7, cell_2085_a_HPC2_and_p_0_out_0__1_,
         cell_2085_a_HPC2_and_p_0_out_1__0_,
         cell_2085_a_HPC2_and_p_1_out_0__1_,
         cell_2085_a_HPC2_and_p_1_out_1__0_,
         cell_2085_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2085_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2085_a_HPC2_and_p_1_in_0__1_, cell_2085_a_HPC2_and_p_1_in_1__0_,
         cell_2085_a_HPC2_and_s_out_0__1_, cell_2085_a_HPC2_and_s_out_1__0_,
         cell_2085_a_HPC2_and_p_0_in_0__1_, cell_2085_a_HPC2_and_p_0_in_1__0_,
         cell_2085_a_HPC2_and_s_in_0__1_, cell_2085_a_HPC2_and_s_in_1__0_,
         cell_2085_a_HPC2_and_z_0__0_, cell_2085_a_HPC2_and_z_1__1_,
         cell_2086_a_HPC2_and_n9, cell_2086_a_HPC2_and_n8,
         cell_2086_a_HPC2_and_n7, cell_2086_a_HPC2_and_p_0_out_0__1_,
         cell_2086_a_HPC2_and_p_0_out_1__0_,
         cell_2086_a_HPC2_and_p_1_out_0__1_,
         cell_2086_a_HPC2_and_p_1_out_1__0_,
         cell_2086_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2086_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2086_a_HPC2_and_p_1_in_0__1_, cell_2086_a_HPC2_and_p_1_in_1__0_,
         cell_2086_a_HPC2_and_s_out_0__1_, cell_2086_a_HPC2_and_s_out_1__0_,
         cell_2086_a_HPC2_and_p_0_in_0__1_, cell_2086_a_HPC2_and_p_0_in_1__0_,
         cell_2086_a_HPC2_and_s_in_0__1_, cell_2086_a_HPC2_and_s_in_1__0_,
         cell_2086_a_HPC2_and_z_0__0_, cell_2086_a_HPC2_and_z_1__1_,
         cell_2087_a_HPC2_and_n9, cell_2087_a_HPC2_and_n8,
         cell_2087_a_HPC2_and_n7, cell_2087_a_HPC2_and_p_0_out_0__1_,
         cell_2087_a_HPC2_and_p_0_out_1__0_,
         cell_2087_a_HPC2_and_p_1_out_0__1_,
         cell_2087_a_HPC2_and_p_1_out_1__0_,
         cell_2087_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2087_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2087_a_HPC2_and_p_1_in_0__1_, cell_2087_a_HPC2_and_p_1_in_1__0_,
         cell_2087_a_HPC2_and_s_out_0__1_, cell_2087_a_HPC2_and_s_out_1__0_,
         cell_2087_a_HPC2_and_p_0_in_0__1_, cell_2087_a_HPC2_and_p_0_in_1__0_,
         cell_2087_a_HPC2_and_s_in_0__1_, cell_2087_a_HPC2_and_s_in_1__0_,
         cell_2087_a_HPC2_and_z_0__0_, cell_2087_a_HPC2_and_z_1__1_,
         cell_2088_a_HPC2_and_n9, cell_2088_a_HPC2_and_n8,
         cell_2088_a_HPC2_and_n7, cell_2088_a_HPC2_and_p_0_out_0__1_,
         cell_2088_a_HPC2_and_p_0_out_1__0_,
         cell_2088_a_HPC2_and_p_1_out_0__1_,
         cell_2088_a_HPC2_and_p_1_out_1__0_,
         cell_2088_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2088_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2088_a_HPC2_and_p_1_in_0__1_, cell_2088_a_HPC2_and_p_1_in_1__0_,
         cell_2088_a_HPC2_and_s_out_0__1_, cell_2088_a_HPC2_and_s_out_1__0_,
         cell_2088_a_HPC2_and_p_0_in_0__1_, cell_2088_a_HPC2_and_p_0_in_1__0_,
         cell_2088_a_HPC2_and_s_in_0__1_, cell_2088_a_HPC2_and_s_in_1__0_,
         cell_2088_a_HPC2_and_z_0__0_, cell_2088_a_HPC2_and_z_1__1_,
         cell_2089_a_HPC2_and_n9, cell_2089_a_HPC2_and_n8,
         cell_2089_a_HPC2_and_n7, cell_2089_a_HPC2_and_p_0_out_0__1_,
         cell_2089_a_HPC2_and_p_0_out_1__0_,
         cell_2089_a_HPC2_and_p_1_out_0__1_,
         cell_2089_a_HPC2_and_p_1_out_1__0_,
         cell_2089_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2089_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2089_a_HPC2_and_p_1_in_0__1_, cell_2089_a_HPC2_and_p_1_in_1__0_,
         cell_2089_a_HPC2_and_s_out_0__1_, cell_2089_a_HPC2_and_s_out_1__0_,
         cell_2089_a_HPC2_and_p_0_in_0__1_, cell_2089_a_HPC2_and_p_0_in_1__0_,
         cell_2089_a_HPC2_and_s_in_0__1_, cell_2089_a_HPC2_and_s_in_1__0_,
         cell_2089_a_HPC2_and_z_0__0_, cell_2089_a_HPC2_and_z_1__1_,
         cell_2090_a_HPC2_and_n9, cell_2090_a_HPC2_and_n8,
         cell_2090_a_HPC2_and_n7, cell_2090_a_HPC2_and_p_0_out_0__1_,
         cell_2090_a_HPC2_and_p_0_out_1__0_,
         cell_2090_a_HPC2_and_p_1_out_0__1_,
         cell_2090_a_HPC2_and_p_1_out_1__0_,
         cell_2090_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2090_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2090_a_HPC2_and_p_1_in_0__1_, cell_2090_a_HPC2_and_p_1_in_1__0_,
         cell_2090_a_HPC2_and_s_out_0__1_, cell_2090_a_HPC2_and_s_out_1__0_,
         cell_2090_a_HPC2_and_p_0_in_0__1_, cell_2090_a_HPC2_and_p_0_in_1__0_,
         cell_2090_a_HPC2_and_s_in_0__1_, cell_2090_a_HPC2_and_s_in_1__0_,
         cell_2090_a_HPC2_and_z_0__0_, cell_2090_a_HPC2_and_z_1__1_,
         cell_2091_a_HPC2_and_n9, cell_2091_a_HPC2_and_n8,
         cell_2091_a_HPC2_and_n7, cell_2091_a_HPC2_and_p_0_out_0__1_,
         cell_2091_a_HPC2_and_p_0_out_1__0_,
         cell_2091_a_HPC2_and_p_1_out_0__1_,
         cell_2091_a_HPC2_and_p_1_out_1__0_,
         cell_2091_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2091_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2091_a_HPC2_and_p_1_in_0__1_, cell_2091_a_HPC2_and_p_1_in_1__0_,
         cell_2091_a_HPC2_and_s_out_0__1_, cell_2091_a_HPC2_and_s_out_1__0_,
         cell_2091_a_HPC2_and_p_0_in_0__1_, cell_2091_a_HPC2_and_p_0_in_1__0_,
         cell_2091_a_HPC2_and_s_in_0__1_, cell_2091_a_HPC2_and_s_in_1__0_,
         cell_2091_a_HPC2_and_z_0__0_, cell_2091_a_HPC2_and_z_1__1_,
         cell_2092_a_HPC2_and_n9, cell_2092_a_HPC2_and_n8,
         cell_2092_a_HPC2_and_n7, cell_2092_a_HPC2_and_p_0_out_0__1_,
         cell_2092_a_HPC2_and_p_0_out_1__0_,
         cell_2092_a_HPC2_and_p_1_out_0__1_,
         cell_2092_a_HPC2_and_p_1_out_1__0_,
         cell_2092_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2092_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2092_a_HPC2_and_p_1_in_0__1_, cell_2092_a_HPC2_and_p_1_in_1__0_,
         cell_2092_a_HPC2_and_s_out_0__1_, cell_2092_a_HPC2_and_s_out_1__0_,
         cell_2092_a_HPC2_and_p_0_in_0__1_, cell_2092_a_HPC2_and_p_0_in_1__0_,
         cell_2092_a_HPC2_and_s_in_0__1_, cell_2092_a_HPC2_and_s_in_1__0_,
         cell_2092_a_HPC2_and_z_0__0_, cell_2092_a_HPC2_and_z_1__1_,
         cell_2093_a_HPC2_and_n9, cell_2093_a_HPC2_and_n8,
         cell_2093_a_HPC2_and_n7, cell_2093_a_HPC2_and_p_0_out_0__1_,
         cell_2093_a_HPC2_and_p_0_out_1__0_,
         cell_2093_a_HPC2_and_p_1_out_0__1_,
         cell_2093_a_HPC2_and_p_1_out_1__0_,
         cell_2093_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2093_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2093_a_HPC2_and_p_1_in_0__1_, cell_2093_a_HPC2_and_p_1_in_1__0_,
         cell_2093_a_HPC2_and_s_out_0__1_, cell_2093_a_HPC2_and_s_out_1__0_,
         cell_2093_a_HPC2_and_p_0_in_0__1_, cell_2093_a_HPC2_and_p_0_in_1__0_,
         cell_2093_a_HPC2_and_s_in_0__1_, cell_2093_a_HPC2_and_s_in_1__0_,
         cell_2093_a_HPC2_and_z_0__0_, cell_2093_a_HPC2_and_z_1__1_,
         cell_2094_a_HPC2_and_n9, cell_2094_a_HPC2_and_n8,
         cell_2094_a_HPC2_and_n7, cell_2094_a_HPC2_and_p_0_out_0__1_,
         cell_2094_a_HPC2_and_p_0_out_1__0_,
         cell_2094_a_HPC2_and_p_1_out_0__1_,
         cell_2094_a_HPC2_and_p_1_out_1__0_,
         cell_2094_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2094_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2094_a_HPC2_and_p_1_in_0__1_, cell_2094_a_HPC2_and_p_1_in_1__0_,
         cell_2094_a_HPC2_and_s_out_0__1_, cell_2094_a_HPC2_and_s_out_1__0_,
         cell_2094_a_HPC2_and_p_0_in_0__1_, cell_2094_a_HPC2_and_p_0_in_1__0_,
         cell_2094_a_HPC2_and_s_in_0__1_, cell_2094_a_HPC2_and_s_in_1__0_,
         cell_2094_a_HPC2_and_z_0__0_, cell_2094_a_HPC2_and_z_1__1_,
         cell_2095_a_HPC2_and_n9, cell_2095_a_HPC2_and_n8,
         cell_2095_a_HPC2_and_n7, cell_2095_a_HPC2_and_p_0_out_0__1_,
         cell_2095_a_HPC2_and_p_0_out_1__0_,
         cell_2095_a_HPC2_and_p_1_out_0__1_,
         cell_2095_a_HPC2_and_p_1_out_1__0_,
         cell_2095_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2095_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2095_a_HPC2_and_p_1_in_0__1_, cell_2095_a_HPC2_and_p_1_in_1__0_,
         cell_2095_a_HPC2_and_s_out_0__1_, cell_2095_a_HPC2_and_s_out_1__0_,
         cell_2095_a_HPC2_and_p_0_in_0__1_, cell_2095_a_HPC2_and_p_0_in_1__0_,
         cell_2095_a_HPC2_and_s_in_0__1_, cell_2095_a_HPC2_and_s_in_1__0_,
         cell_2095_a_HPC2_and_z_0__0_, cell_2095_a_HPC2_and_z_1__1_,
         cell_2096_a_HPC2_and_n9, cell_2096_a_HPC2_and_n8,
         cell_2096_a_HPC2_and_n7, cell_2096_a_HPC2_and_p_0_out_0__1_,
         cell_2096_a_HPC2_and_p_0_out_1__0_,
         cell_2096_a_HPC2_and_p_1_out_0__1_,
         cell_2096_a_HPC2_and_p_1_out_1__0_,
         cell_2096_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2096_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2096_a_HPC2_and_p_1_in_0__1_, cell_2096_a_HPC2_and_p_1_in_1__0_,
         cell_2096_a_HPC2_and_s_out_0__1_, cell_2096_a_HPC2_and_s_out_1__0_,
         cell_2096_a_HPC2_and_p_0_in_0__1_, cell_2096_a_HPC2_and_p_0_in_1__0_,
         cell_2096_a_HPC2_and_s_in_0__1_, cell_2096_a_HPC2_and_s_in_1__0_,
         cell_2096_a_HPC2_and_z_0__0_, cell_2096_a_HPC2_and_z_1__1_,
         cell_2097_a_HPC2_and_n9, cell_2097_a_HPC2_and_n8,
         cell_2097_a_HPC2_and_n7, cell_2097_a_HPC2_and_p_0_out_0__1_,
         cell_2097_a_HPC2_and_p_0_out_1__0_,
         cell_2097_a_HPC2_and_p_1_out_0__1_,
         cell_2097_a_HPC2_and_p_1_out_1__0_,
         cell_2097_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2097_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2097_a_HPC2_and_p_1_in_0__1_, cell_2097_a_HPC2_and_p_1_in_1__0_,
         cell_2097_a_HPC2_and_s_out_0__1_, cell_2097_a_HPC2_and_s_out_1__0_,
         cell_2097_a_HPC2_and_p_0_in_0__1_, cell_2097_a_HPC2_and_p_0_in_1__0_,
         cell_2097_a_HPC2_and_s_in_0__1_, cell_2097_a_HPC2_and_s_in_1__0_,
         cell_2097_a_HPC2_and_z_0__0_, cell_2097_a_HPC2_and_z_1__1_,
         cell_2098_a_HPC2_and_n9, cell_2098_a_HPC2_and_n8,
         cell_2098_a_HPC2_and_n7, cell_2098_a_HPC2_and_p_0_out_0__1_,
         cell_2098_a_HPC2_and_p_0_out_1__0_,
         cell_2098_a_HPC2_and_p_1_out_0__1_,
         cell_2098_a_HPC2_and_p_1_out_1__0_,
         cell_2098_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2098_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2098_a_HPC2_and_p_1_in_0__1_, cell_2098_a_HPC2_and_p_1_in_1__0_,
         cell_2098_a_HPC2_and_s_out_0__1_, cell_2098_a_HPC2_and_s_out_1__0_,
         cell_2098_a_HPC2_and_p_0_in_0__1_, cell_2098_a_HPC2_and_p_0_in_1__0_,
         cell_2098_a_HPC2_and_s_in_0__1_, cell_2098_a_HPC2_and_s_in_1__0_,
         cell_2098_a_HPC2_and_z_0__0_, cell_2098_a_HPC2_and_z_1__1_,
         cell_2099_a_HPC2_and_n9, cell_2099_a_HPC2_and_n8,
         cell_2099_a_HPC2_and_n7, cell_2099_a_HPC2_and_p_0_out_0__1_,
         cell_2099_a_HPC2_and_p_0_out_1__0_,
         cell_2099_a_HPC2_and_p_1_out_0__1_,
         cell_2099_a_HPC2_and_p_1_out_1__0_,
         cell_2099_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2099_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2099_a_HPC2_and_p_1_in_0__1_, cell_2099_a_HPC2_and_p_1_in_1__0_,
         cell_2099_a_HPC2_and_s_out_0__1_, cell_2099_a_HPC2_and_s_out_1__0_,
         cell_2099_a_HPC2_and_p_0_in_0__1_, cell_2099_a_HPC2_and_p_0_in_1__0_,
         cell_2099_a_HPC2_and_s_in_0__1_, cell_2099_a_HPC2_and_s_in_1__0_,
         cell_2099_a_HPC2_and_z_0__0_, cell_2099_a_HPC2_and_z_1__1_,
         cell_2100_a_HPC2_and_n9, cell_2100_a_HPC2_and_n8,
         cell_2100_a_HPC2_and_n7, cell_2100_a_HPC2_and_p_0_out_0__1_,
         cell_2100_a_HPC2_and_p_0_out_1__0_,
         cell_2100_a_HPC2_and_p_1_out_0__1_,
         cell_2100_a_HPC2_and_p_1_out_1__0_,
         cell_2100_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2100_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2100_a_HPC2_and_p_1_in_0__1_, cell_2100_a_HPC2_and_p_1_in_1__0_,
         cell_2100_a_HPC2_and_s_out_0__1_, cell_2100_a_HPC2_and_s_out_1__0_,
         cell_2100_a_HPC2_and_p_0_in_0__1_, cell_2100_a_HPC2_and_p_0_in_1__0_,
         cell_2100_a_HPC2_and_s_in_0__1_, cell_2100_a_HPC2_and_s_in_1__0_,
         cell_2100_a_HPC2_and_z_0__0_, cell_2100_a_HPC2_and_z_1__1_,
         cell_2101_a_HPC2_and_n9, cell_2101_a_HPC2_and_n8,
         cell_2101_a_HPC2_and_n7, cell_2101_a_HPC2_and_p_0_out_0__1_,
         cell_2101_a_HPC2_and_p_0_out_1__0_,
         cell_2101_a_HPC2_and_p_1_out_0__1_,
         cell_2101_a_HPC2_and_p_1_out_1__0_,
         cell_2101_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2101_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2101_a_HPC2_and_p_1_in_0__1_, cell_2101_a_HPC2_and_p_1_in_1__0_,
         cell_2101_a_HPC2_and_s_out_0__1_, cell_2101_a_HPC2_and_s_out_1__0_,
         cell_2101_a_HPC2_and_p_0_in_0__1_, cell_2101_a_HPC2_and_p_0_in_1__0_,
         cell_2101_a_HPC2_and_s_in_0__1_, cell_2101_a_HPC2_and_s_in_1__0_,
         cell_2101_a_HPC2_and_z_0__0_, cell_2101_a_HPC2_and_z_1__1_,
         cell_2102_a_HPC2_and_n9, cell_2102_a_HPC2_and_n8,
         cell_2102_a_HPC2_and_n7, cell_2102_a_HPC2_and_p_0_out_0__1_,
         cell_2102_a_HPC2_and_p_0_out_1__0_,
         cell_2102_a_HPC2_and_p_1_out_0__1_,
         cell_2102_a_HPC2_and_p_1_out_1__0_,
         cell_2102_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2102_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2102_a_HPC2_and_p_1_in_0__1_, cell_2102_a_HPC2_and_p_1_in_1__0_,
         cell_2102_a_HPC2_and_s_out_0__1_, cell_2102_a_HPC2_and_s_out_1__0_,
         cell_2102_a_HPC2_and_p_0_in_0__1_, cell_2102_a_HPC2_and_p_0_in_1__0_,
         cell_2102_a_HPC2_and_s_in_0__1_, cell_2102_a_HPC2_and_s_in_1__0_,
         cell_2102_a_HPC2_and_z_0__0_, cell_2102_a_HPC2_and_z_1__1_,
         cell_2103_a_HPC2_and_n9, cell_2103_a_HPC2_and_n8,
         cell_2103_a_HPC2_and_n7, cell_2103_a_HPC2_and_p_0_out_0__1_,
         cell_2103_a_HPC2_and_p_0_out_1__0_,
         cell_2103_a_HPC2_and_p_1_out_0__1_,
         cell_2103_a_HPC2_and_p_1_out_1__0_,
         cell_2103_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2103_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2103_a_HPC2_and_p_1_in_0__1_, cell_2103_a_HPC2_and_p_1_in_1__0_,
         cell_2103_a_HPC2_and_s_out_0__1_, cell_2103_a_HPC2_and_s_out_1__0_,
         cell_2103_a_HPC2_and_p_0_in_0__1_, cell_2103_a_HPC2_and_p_0_in_1__0_,
         cell_2103_a_HPC2_and_s_in_0__1_, cell_2103_a_HPC2_and_s_in_1__0_,
         cell_2103_a_HPC2_and_z_0__0_, cell_2103_a_HPC2_and_z_1__1_,
         cell_2104_a_HPC2_and_n9, cell_2104_a_HPC2_and_n8,
         cell_2104_a_HPC2_and_n7, cell_2104_a_HPC2_and_p_0_out_0__1_,
         cell_2104_a_HPC2_and_p_0_out_1__0_,
         cell_2104_a_HPC2_and_p_1_out_0__1_,
         cell_2104_a_HPC2_and_p_1_out_1__0_,
         cell_2104_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2104_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2104_a_HPC2_and_p_1_in_0__1_, cell_2104_a_HPC2_and_p_1_in_1__0_,
         cell_2104_a_HPC2_and_s_out_0__1_, cell_2104_a_HPC2_and_s_out_1__0_,
         cell_2104_a_HPC2_and_p_0_in_0__1_, cell_2104_a_HPC2_and_p_0_in_1__0_,
         cell_2104_a_HPC2_and_s_in_0__1_, cell_2104_a_HPC2_and_s_in_1__0_,
         cell_2104_a_HPC2_and_z_0__0_, cell_2104_a_HPC2_and_z_1__1_,
         cell_2105_a_HPC2_and_n9, cell_2105_a_HPC2_and_n8,
         cell_2105_a_HPC2_and_n7, cell_2105_a_HPC2_and_p_0_out_0__1_,
         cell_2105_a_HPC2_and_p_0_out_1__0_,
         cell_2105_a_HPC2_and_p_1_out_0__1_,
         cell_2105_a_HPC2_and_p_1_out_1__0_,
         cell_2105_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2105_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2105_a_HPC2_and_p_1_in_0__1_, cell_2105_a_HPC2_and_p_1_in_1__0_,
         cell_2105_a_HPC2_and_s_out_0__1_, cell_2105_a_HPC2_and_s_out_1__0_,
         cell_2105_a_HPC2_and_p_0_in_0__1_, cell_2105_a_HPC2_and_p_0_in_1__0_,
         cell_2105_a_HPC2_and_s_in_0__1_, cell_2105_a_HPC2_and_s_in_1__0_,
         cell_2105_a_HPC2_and_z_0__0_, cell_2105_a_HPC2_and_z_1__1_,
         cell_2106_a_HPC2_and_n9, cell_2106_a_HPC2_and_n8,
         cell_2106_a_HPC2_and_n7, cell_2106_a_HPC2_and_p_0_out_0__1_,
         cell_2106_a_HPC2_and_p_0_out_1__0_,
         cell_2106_a_HPC2_and_p_1_out_0__1_,
         cell_2106_a_HPC2_and_p_1_out_1__0_,
         cell_2106_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2106_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2106_a_HPC2_and_p_1_in_0__1_, cell_2106_a_HPC2_and_p_1_in_1__0_,
         cell_2106_a_HPC2_and_s_out_0__1_, cell_2106_a_HPC2_and_s_out_1__0_,
         cell_2106_a_HPC2_and_p_0_in_0__1_, cell_2106_a_HPC2_and_p_0_in_1__0_,
         cell_2106_a_HPC2_and_s_in_0__1_, cell_2106_a_HPC2_and_s_in_1__0_,
         cell_2106_a_HPC2_and_z_0__0_, cell_2106_a_HPC2_and_z_1__1_,
         cell_2107_a_HPC2_and_n9, cell_2107_a_HPC2_and_n8,
         cell_2107_a_HPC2_and_n7, cell_2107_a_HPC2_and_p_0_out_0__1_,
         cell_2107_a_HPC2_and_p_0_out_1__0_,
         cell_2107_a_HPC2_and_p_1_out_0__1_,
         cell_2107_a_HPC2_and_p_1_out_1__0_,
         cell_2107_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2107_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2107_a_HPC2_and_p_1_in_0__1_, cell_2107_a_HPC2_and_p_1_in_1__0_,
         cell_2107_a_HPC2_and_s_out_0__1_, cell_2107_a_HPC2_and_s_out_1__0_,
         cell_2107_a_HPC2_and_p_0_in_0__1_, cell_2107_a_HPC2_and_p_0_in_1__0_,
         cell_2107_a_HPC2_and_s_in_0__1_, cell_2107_a_HPC2_and_s_in_1__0_,
         cell_2107_a_HPC2_and_z_0__0_, cell_2107_a_HPC2_and_z_1__1_,
         cell_2108_a_HPC2_and_n9, cell_2108_a_HPC2_and_n8,
         cell_2108_a_HPC2_and_n7, cell_2108_a_HPC2_and_p_0_out_0__1_,
         cell_2108_a_HPC2_and_p_0_out_1__0_,
         cell_2108_a_HPC2_and_p_1_out_0__1_,
         cell_2108_a_HPC2_and_p_1_out_1__0_,
         cell_2108_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2108_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2108_a_HPC2_and_p_1_in_0__1_, cell_2108_a_HPC2_and_p_1_in_1__0_,
         cell_2108_a_HPC2_and_s_out_0__1_, cell_2108_a_HPC2_and_s_out_1__0_,
         cell_2108_a_HPC2_and_p_0_in_0__1_, cell_2108_a_HPC2_and_p_0_in_1__0_,
         cell_2108_a_HPC2_and_s_in_0__1_, cell_2108_a_HPC2_and_s_in_1__0_,
         cell_2108_a_HPC2_and_z_0__0_, cell_2108_a_HPC2_and_z_1__1_,
         cell_2109_a_HPC2_and_n9, cell_2109_a_HPC2_and_n8,
         cell_2109_a_HPC2_and_n7, cell_2109_a_HPC2_and_p_0_out_0__1_,
         cell_2109_a_HPC2_and_p_0_out_1__0_,
         cell_2109_a_HPC2_and_p_1_out_0__1_,
         cell_2109_a_HPC2_and_p_1_out_1__0_,
         cell_2109_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2109_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2109_a_HPC2_and_p_1_in_0__1_, cell_2109_a_HPC2_and_p_1_in_1__0_,
         cell_2109_a_HPC2_and_s_out_0__1_, cell_2109_a_HPC2_and_s_out_1__0_,
         cell_2109_a_HPC2_and_p_0_in_0__1_, cell_2109_a_HPC2_and_p_0_in_1__0_,
         cell_2109_a_HPC2_and_s_in_0__1_, cell_2109_a_HPC2_and_s_in_1__0_,
         cell_2109_a_HPC2_and_z_0__0_, cell_2109_a_HPC2_and_z_1__1_,
         cell_2110_a_HPC2_and_n9, cell_2110_a_HPC2_and_n8,
         cell_2110_a_HPC2_and_n7, cell_2110_a_HPC2_and_p_0_out_0__1_,
         cell_2110_a_HPC2_and_p_0_out_1__0_,
         cell_2110_a_HPC2_and_p_1_out_0__1_,
         cell_2110_a_HPC2_and_p_1_out_1__0_,
         cell_2110_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2110_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2110_a_HPC2_and_p_1_in_0__1_, cell_2110_a_HPC2_and_p_1_in_1__0_,
         cell_2110_a_HPC2_and_s_out_0__1_, cell_2110_a_HPC2_and_s_out_1__0_,
         cell_2110_a_HPC2_and_p_0_in_0__1_, cell_2110_a_HPC2_and_p_0_in_1__0_,
         cell_2110_a_HPC2_and_s_in_0__1_, cell_2110_a_HPC2_and_s_in_1__0_,
         cell_2110_a_HPC2_and_z_0__0_, cell_2110_a_HPC2_and_z_1__1_,
         cell_2111_a_HPC2_and_n9, cell_2111_a_HPC2_and_n8,
         cell_2111_a_HPC2_and_n7, cell_2111_a_HPC2_and_p_0_out_0__1_,
         cell_2111_a_HPC2_and_p_0_out_1__0_,
         cell_2111_a_HPC2_and_p_1_out_0__1_,
         cell_2111_a_HPC2_and_p_1_out_1__0_,
         cell_2111_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2111_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2111_a_HPC2_and_p_1_in_0__1_, cell_2111_a_HPC2_and_p_1_in_1__0_,
         cell_2111_a_HPC2_and_s_out_0__1_, cell_2111_a_HPC2_and_s_out_1__0_,
         cell_2111_a_HPC2_and_p_0_in_0__1_, cell_2111_a_HPC2_and_p_0_in_1__0_,
         cell_2111_a_HPC2_and_s_in_0__1_, cell_2111_a_HPC2_and_s_in_1__0_,
         cell_2111_a_HPC2_and_z_0__0_, cell_2111_a_HPC2_and_z_1__1_,
         cell_2112_a_HPC2_and_n9, cell_2112_a_HPC2_and_n8,
         cell_2112_a_HPC2_and_n7, cell_2112_a_HPC2_and_p_0_out_0__1_,
         cell_2112_a_HPC2_and_p_0_out_1__0_,
         cell_2112_a_HPC2_and_p_1_out_0__1_,
         cell_2112_a_HPC2_and_p_1_out_1__0_,
         cell_2112_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2112_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2112_a_HPC2_and_p_1_in_0__1_, cell_2112_a_HPC2_and_p_1_in_1__0_,
         cell_2112_a_HPC2_and_s_out_0__1_, cell_2112_a_HPC2_and_s_out_1__0_,
         cell_2112_a_HPC2_and_p_0_in_0__1_, cell_2112_a_HPC2_and_p_0_in_1__0_,
         cell_2112_a_HPC2_and_s_in_0__1_, cell_2112_a_HPC2_and_s_in_1__0_,
         cell_2112_a_HPC2_and_z_0__0_, cell_2112_a_HPC2_and_z_1__1_,
         cell_2113_a_HPC2_and_n9, cell_2113_a_HPC2_and_n8,
         cell_2113_a_HPC2_and_n7, cell_2113_a_HPC2_and_p_0_out_0__1_,
         cell_2113_a_HPC2_and_p_0_out_1__0_,
         cell_2113_a_HPC2_and_p_1_out_0__1_,
         cell_2113_a_HPC2_and_p_1_out_1__0_,
         cell_2113_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2113_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2113_a_HPC2_and_p_1_in_0__1_, cell_2113_a_HPC2_and_p_1_in_1__0_,
         cell_2113_a_HPC2_and_s_out_0__1_, cell_2113_a_HPC2_and_s_out_1__0_,
         cell_2113_a_HPC2_and_p_0_in_0__1_, cell_2113_a_HPC2_and_p_0_in_1__0_,
         cell_2113_a_HPC2_and_s_in_0__1_, cell_2113_a_HPC2_and_s_in_1__0_,
         cell_2113_a_HPC2_and_z_0__0_, cell_2113_a_HPC2_and_z_1__1_,
         cell_2114_a_HPC2_and_n9, cell_2114_a_HPC2_and_n8,
         cell_2114_a_HPC2_and_n7, cell_2114_a_HPC2_and_p_0_out_0__1_,
         cell_2114_a_HPC2_and_p_0_out_1__0_,
         cell_2114_a_HPC2_and_p_1_out_0__1_,
         cell_2114_a_HPC2_and_p_1_out_1__0_,
         cell_2114_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2114_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2114_a_HPC2_and_p_1_in_0__1_, cell_2114_a_HPC2_and_p_1_in_1__0_,
         cell_2114_a_HPC2_and_s_out_0__1_, cell_2114_a_HPC2_and_s_out_1__0_,
         cell_2114_a_HPC2_and_p_0_in_0__1_, cell_2114_a_HPC2_and_p_0_in_1__0_,
         cell_2114_a_HPC2_and_s_in_0__1_, cell_2114_a_HPC2_and_s_in_1__0_,
         cell_2114_a_HPC2_and_z_0__0_, cell_2114_a_HPC2_and_z_1__1_,
         cell_2115_a_HPC2_and_n9, cell_2115_a_HPC2_and_n8,
         cell_2115_a_HPC2_and_n7, cell_2115_a_HPC2_and_p_0_out_0__1_,
         cell_2115_a_HPC2_and_p_0_out_1__0_,
         cell_2115_a_HPC2_and_p_1_out_0__1_,
         cell_2115_a_HPC2_and_p_1_out_1__0_,
         cell_2115_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2115_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2115_a_HPC2_and_p_1_in_0__1_, cell_2115_a_HPC2_and_p_1_in_1__0_,
         cell_2115_a_HPC2_and_s_out_0__1_, cell_2115_a_HPC2_and_s_out_1__0_,
         cell_2115_a_HPC2_and_p_0_in_0__1_, cell_2115_a_HPC2_and_p_0_in_1__0_,
         cell_2115_a_HPC2_and_s_in_0__1_, cell_2115_a_HPC2_and_s_in_1__0_,
         cell_2115_a_HPC2_and_z_0__0_, cell_2115_a_HPC2_and_z_1__1_,
         cell_2116_a_HPC2_and_n9, cell_2116_a_HPC2_and_n8,
         cell_2116_a_HPC2_and_n7, cell_2116_a_HPC2_and_p_0_out_0__1_,
         cell_2116_a_HPC2_and_p_0_out_1__0_,
         cell_2116_a_HPC2_and_p_1_out_0__1_,
         cell_2116_a_HPC2_and_p_1_out_1__0_,
         cell_2116_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2116_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2116_a_HPC2_and_p_1_in_0__1_, cell_2116_a_HPC2_and_p_1_in_1__0_,
         cell_2116_a_HPC2_and_s_out_0__1_, cell_2116_a_HPC2_and_s_out_1__0_,
         cell_2116_a_HPC2_and_p_0_in_0__1_, cell_2116_a_HPC2_and_p_0_in_1__0_,
         cell_2116_a_HPC2_and_s_in_0__1_, cell_2116_a_HPC2_and_s_in_1__0_,
         cell_2116_a_HPC2_and_z_0__0_, cell_2116_a_HPC2_and_z_1__1_,
         cell_2117_a_HPC2_and_n9, cell_2117_a_HPC2_and_n8,
         cell_2117_a_HPC2_and_n7, cell_2117_a_HPC2_and_p_0_out_0__1_,
         cell_2117_a_HPC2_and_p_0_out_1__0_,
         cell_2117_a_HPC2_and_p_1_out_0__1_,
         cell_2117_a_HPC2_and_p_1_out_1__0_,
         cell_2117_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2117_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2117_a_HPC2_and_p_1_in_0__1_, cell_2117_a_HPC2_and_p_1_in_1__0_,
         cell_2117_a_HPC2_and_s_out_0__1_, cell_2117_a_HPC2_and_s_out_1__0_,
         cell_2117_a_HPC2_and_p_0_in_0__1_, cell_2117_a_HPC2_and_p_0_in_1__0_,
         cell_2117_a_HPC2_and_s_in_0__1_, cell_2117_a_HPC2_and_s_in_1__0_,
         cell_2117_a_HPC2_and_z_0__0_, cell_2117_a_HPC2_and_z_1__1_,
         cell_2118_a_HPC2_and_n9, cell_2118_a_HPC2_and_n8,
         cell_2118_a_HPC2_and_n7, cell_2118_a_HPC2_and_p_0_out_0__1_,
         cell_2118_a_HPC2_and_p_0_out_1__0_,
         cell_2118_a_HPC2_and_p_1_out_0__1_,
         cell_2118_a_HPC2_and_p_1_out_1__0_,
         cell_2118_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2118_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2118_a_HPC2_and_p_1_in_0__1_, cell_2118_a_HPC2_and_p_1_in_1__0_,
         cell_2118_a_HPC2_and_s_out_0__1_, cell_2118_a_HPC2_and_s_out_1__0_,
         cell_2118_a_HPC2_and_p_0_in_0__1_, cell_2118_a_HPC2_and_p_0_in_1__0_,
         cell_2118_a_HPC2_and_s_in_0__1_, cell_2118_a_HPC2_and_s_in_1__0_,
         cell_2118_a_HPC2_and_z_0__0_, cell_2118_a_HPC2_and_z_1__1_,
         cell_2119_a_HPC2_and_n9, cell_2119_a_HPC2_and_n8,
         cell_2119_a_HPC2_and_n7, cell_2119_a_HPC2_and_p_0_out_0__1_,
         cell_2119_a_HPC2_and_p_0_out_1__0_,
         cell_2119_a_HPC2_and_p_1_out_0__1_,
         cell_2119_a_HPC2_and_p_1_out_1__0_,
         cell_2119_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2119_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2119_a_HPC2_and_p_1_in_0__1_, cell_2119_a_HPC2_and_p_1_in_1__0_,
         cell_2119_a_HPC2_and_s_out_0__1_, cell_2119_a_HPC2_and_s_out_1__0_,
         cell_2119_a_HPC2_and_p_0_in_0__1_, cell_2119_a_HPC2_and_p_0_in_1__0_,
         cell_2119_a_HPC2_and_s_in_0__1_, cell_2119_a_HPC2_and_s_in_1__0_,
         cell_2119_a_HPC2_and_z_0__0_, cell_2119_a_HPC2_and_z_1__1_,
         cell_2120_a_HPC2_and_n9, cell_2120_a_HPC2_and_n8,
         cell_2120_a_HPC2_and_n7, cell_2120_a_HPC2_and_p_0_out_0__1_,
         cell_2120_a_HPC2_and_p_0_out_1__0_,
         cell_2120_a_HPC2_and_p_1_out_0__1_,
         cell_2120_a_HPC2_and_p_1_out_1__0_,
         cell_2120_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2120_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2120_a_HPC2_and_p_1_in_0__1_, cell_2120_a_HPC2_and_p_1_in_1__0_,
         cell_2120_a_HPC2_and_s_out_0__1_, cell_2120_a_HPC2_and_s_out_1__0_,
         cell_2120_a_HPC2_and_p_0_in_0__1_, cell_2120_a_HPC2_and_p_0_in_1__0_,
         cell_2120_a_HPC2_and_s_in_0__1_, cell_2120_a_HPC2_and_s_in_1__0_,
         cell_2120_a_HPC2_and_z_0__0_, cell_2120_a_HPC2_and_z_1__1_,
         cell_2121_a_HPC2_and_n9, cell_2121_a_HPC2_and_n8,
         cell_2121_a_HPC2_and_n7, cell_2121_a_HPC2_and_p_0_out_0__1_,
         cell_2121_a_HPC2_and_p_0_out_1__0_,
         cell_2121_a_HPC2_and_p_1_out_0__1_,
         cell_2121_a_HPC2_and_p_1_out_1__0_,
         cell_2121_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2121_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2121_a_HPC2_and_p_1_in_0__1_, cell_2121_a_HPC2_and_p_1_in_1__0_,
         cell_2121_a_HPC2_and_s_out_0__1_, cell_2121_a_HPC2_and_s_out_1__0_,
         cell_2121_a_HPC2_and_p_0_in_0__1_, cell_2121_a_HPC2_and_p_0_in_1__0_,
         cell_2121_a_HPC2_and_s_in_0__1_, cell_2121_a_HPC2_and_s_in_1__0_,
         cell_2121_a_HPC2_and_z_0__0_, cell_2121_a_HPC2_and_z_1__1_,
         cell_2122_a_HPC2_and_n9, cell_2122_a_HPC2_and_n8,
         cell_2122_a_HPC2_and_n7, cell_2122_a_HPC2_and_p_0_out_0__1_,
         cell_2122_a_HPC2_and_p_0_out_1__0_,
         cell_2122_a_HPC2_and_p_1_out_0__1_,
         cell_2122_a_HPC2_and_p_1_out_1__0_,
         cell_2122_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2122_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2122_a_HPC2_and_p_1_in_0__1_, cell_2122_a_HPC2_and_p_1_in_1__0_,
         cell_2122_a_HPC2_and_s_out_0__1_, cell_2122_a_HPC2_and_s_out_1__0_,
         cell_2122_a_HPC2_and_p_0_in_0__1_, cell_2122_a_HPC2_and_p_0_in_1__0_,
         cell_2122_a_HPC2_and_s_in_0__1_, cell_2122_a_HPC2_and_s_in_1__0_,
         cell_2122_a_HPC2_and_z_0__0_, cell_2122_a_HPC2_and_z_1__1_,
         cell_2123_a_HPC2_and_n9, cell_2123_a_HPC2_and_n8,
         cell_2123_a_HPC2_and_n7, cell_2123_a_HPC2_and_p_0_out_0__1_,
         cell_2123_a_HPC2_and_p_0_out_1__0_,
         cell_2123_a_HPC2_and_p_1_out_0__1_,
         cell_2123_a_HPC2_and_p_1_out_1__0_,
         cell_2123_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2123_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2123_a_HPC2_and_p_1_in_0__1_, cell_2123_a_HPC2_and_p_1_in_1__0_,
         cell_2123_a_HPC2_and_s_out_0__1_, cell_2123_a_HPC2_and_s_out_1__0_,
         cell_2123_a_HPC2_and_p_0_in_0__1_, cell_2123_a_HPC2_and_p_0_in_1__0_,
         cell_2123_a_HPC2_and_s_in_0__1_, cell_2123_a_HPC2_and_s_in_1__0_,
         cell_2123_a_HPC2_and_z_0__0_, cell_2123_a_HPC2_and_z_1__1_,
         cell_2124_a_HPC2_and_n9, cell_2124_a_HPC2_and_n8,
         cell_2124_a_HPC2_and_n7, cell_2124_a_HPC2_and_p_0_out_0__1_,
         cell_2124_a_HPC2_and_p_0_out_1__0_,
         cell_2124_a_HPC2_and_p_1_out_0__1_,
         cell_2124_a_HPC2_and_p_1_out_1__0_,
         cell_2124_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2124_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2124_a_HPC2_and_p_1_in_0__1_, cell_2124_a_HPC2_and_p_1_in_1__0_,
         cell_2124_a_HPC2_and_s_out_0__1_, cell_2124_a_HPC2_and_s_out_1__0_,
         cell_2124_a_HPC2_and_p_0_in_0__1_, cell_2124_a_HPC2_and_p_0_in_1__0_,
         cell_2124_a_HPC2_and_s_in_0__1_, cell_2124_a_HPC2_and_s_in_1__0_,
         cell_2124_a_HPC2_and_z_0__0_, cell_2124_a_HPC2_and_z_1__1_,
         cell_2125_a_HPC2_and_n9, cell_2125_a_HPC2_and_n8,
         cell_2125_a_HPC2_and_n7, cell_2125_a_HPC2_and_p_0_out_0__1_,
         cell_2125_a_HPC2_and_p_0_out_1__0_,
         cell_2125_a_HPC2_and_p_1_out_0__1_,
         cell_2125_a_HPC2_and_p_1_out_1__0_,
         cell_2125_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2125_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2125_a_HPC2_and_p_1_in_0__1_, cell_2125_a_HPC2_and_p_1_in_1__0_,
         cell_2125_a_HPC2_and_s_out_0__1_, cell_2125_a_HPC2_and_s_out_1__0_,
         cell_2125_a_HPC2_and_p_0_in_0__1_, cell_2125_a_HPC2_and_p_0_in_1__0_,
         cell_2125_a_HPC2_and_s_in_0__1_, cell_2125_a_HPC2_and_s_in_1__0_,
         cell_2125_a_HPC2_and_z_0__0_, cell_2125_a_HPC2_and_z_1__1_,
         cell_2126_a_HPC2_and_n9, cell_2126_a_HPC2_and_n8,
         cell_2126_a_HPC2_and_n7, cell_2126_a_HPC2_and_p_0_out_0__1_,
         cell_2126_a_HPC2_and_p_0_out_1__0_,
         cell_2126_a_HPC2_and_p_1_out_0__1_,
         cell_2126_a_HPC2_and_p_1_out_1__0_,
         cell_2126_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2126_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2126_a_HPC2_and_p_1_in_0__1_, cell_2126_a_HPC2_and_p_1_in_1__0_,
         cell_2126_a_HPC2_and_s_out_0__1_, cell_2126_a_HPC2_and_s_out_1__0_,
         cell_2126_a_HPC2_and_p_0_in_0__1_, cell_2126_a_HPC2_and_p_0_in_1__0_,
         cell_2126_a_HPC2_and_s_in_0__1_, cell_2126_a_HPC2_and_s_in_1__0_,
         cell_2126_a_HPC2_and_z_0__0_, cell_2126_a_HPC2_and_z_1__1_,
         cell_2127_a_HPC2_and_n9, cell_2127_a_HPC2_and_n8,
         cell_2127_a_HPC2_and_n7, cell_2127_a_HPC2_and_p_0_out_0__1_,
         cell_2127_a_HPC2_and_p_0_out_1__0_,
         cell_2127_a_HPC2_and_p_1_out_0__1_,
         cell_2127_a_HPC2_and_p_1_out_1__0_,
         cell_2127_a_HPC2_and_p_0_pipe_out_0__1_,
         cell_2127_a_HPC2_and_p_0_pipe_out_1__0_,
         cell_2127_a_HPC2_and_p_1_in_0__1_, cell_2127_a_HPC2_and_p_1_in_1__0_,
         cell_2127_a_HPC2_and_s_out_0__1_, cell_2127_a_HPC2_and_s_out_1__0_,
         cell_2127_a_HPC2_and_p_0_in_0__1_, cell_2127_a_HPC2_and_p_0_in_1__0_,
         cell_2127_a_HPC2_and_s_in_0__1_, cell_2127_a_HPC2_and_s_in_1__0_,
         cell_2127_a_HPC2_and_z_0__0_, cell_2127_a_HPC2_and_z_1__1_;
  wire   [1:0] cell_1714_and_out;
  wire   [1:0] cell_1714_and_in;
  wire   [1:0] cell_1714_a_HPC2_and_a_reg;
  wire   [1:0] cell_1714_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1714_a_HPC2_and_mul;
  wire   [1:0] cell_1715_and_out;
  wire   [1:0] cell_1715_and_in;
  wire   [1:0] cell_1715_a_HPC2_and_a_reg;
  wire   [1:0] cell_1715_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1715_a_HPC2_and_mul;
  wire   [1:0] cell_1716_and_out;
  wire   [1:0] cell_1716_and_in;
  wire   [1:0] cell_1716_a_HPC2_and_a_reg;
  wire   [1:0] cell_1716_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1716_a_HPC2_and_mul;
  wire   [1:0] cell_1717_and_out;
  wire   [1:0] cell_1717_and_in;
  wire   [1:0] cell_1717_a_HPC2_and_a_reg;
  wire   [1:0] cell_1717_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1717_a_HPC2_and_mul;
  wire   [1:0] cell_1718_and_out;
  wire   [1:0] cell_1718_and_in;
  wire   [1:0] cell_1718_a_HPC2_and_a_reg;
  wire   [1:0] cell_1718_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1718_a_HPC2_and_mul;
  wire   [1:0] cell_1719_and_out;
  wire   [1:0] cell_1719_and_in;
  wire   [1:0] cell_1719_a_HPC2_and_a_reg;
  wire   [1:0] cell_1719_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1719_a_HPC2_and_mul;
  wire   [1:0] cell_1720_and_out;
  wire   [1:0] cell_1720_and_in;
  wire   [1:0] cell_1720_a_HPC2_and_a_reg;
  wire   [1:0] cell_1720_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1720_a_HPC2_and_mul;
  wire   [1:0] cell_1721_and_out;
  wire   [1:0] cell_1721_and_in;
  wire   [1:0] cell_1721_a_HPC2_and_a_reg;
  wire   [1:0] cell_1721_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1721_a_HPC2_and_mul;
  wire   [1:0] cell_1722_and_out;
  wire   [1:0] cell_1722_and_in;
  wire   [1:0] cell_1722_a_HPC2_and_a_reg;
  wire   [1:0] cell_1722_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1722_a_HPC2_and_mul;
  wire   [1:0] cell_1723_and_out;
  wire   [1:0] cell_1723_and_in;
  wire   [1:0] cell_1723_a_HPC2_and_a_reg;
  wire   [1:0] cell_1723_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1723_a_HPC2_and_mul;
  wire   [1:0] cell_1724_and_out;
  wire   [1:0] cell_1724_and_in;
  wire   [1:0] cell_1724_a_HPC2_and_a_reg;
  wire   [1:0] cell_1724_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1724_a_HPC2_and_mul;
  wire   [1:0] cell_1725_and_out;
  wire   [1:0] cell_1725_and_in;
  wire   [1:0] cell_1725_a_HPC2_and_a_reg;
  wire   [1:0] cell_1725_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1725_a_HPC2_and_mul;
  wire   [1:0] cell_1726_and_out;
  wire   [1:0] cell_1726_and_in;
  wire   [1:0] cell_1726_a_HPC2_and_a_reg;
  wire   [1:0] cell_1726_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1726_a_HPC2_and_mul;
  wire   [1:0] cell_1727_and_out;
  wire   [1:0] cell_1727_and_in;
  wire   [1:0] cell_1727_a_HPC2_and_a_reg;
  wire   [1:0] cell_1727_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1727_a_HPC2_and_mul;
  wire   [1:0] cell_1728_and_out;
  wire   [1:0] cell_1728_and_in;
  wire   [1:0] cell_1728_a_HPC2_and_a_reg;
  wire   [1:0] cell_1728_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1728_a_HPC2_and_mul;
  wire   [1:0] cell_1729_and_out;
  wire   [1:0] cell_1729_and_in;
  wire   [1:0] cell_1729_a_HPC2_and_a_reg;
  wire   [1:0] cell_1729_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1729_a_HPC2_and_mul;
  wire   [1:0] cell_1730_and_out;
  wire   [1:0] cell_1730_and_in;
  wire   [1:0] cell_1730_a_HPC2_and_a_reg;
  wire   [1:0] cell_1730_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1730_a_HPC2_and_mul;
  wire   [1:0] cell_1731_and_out;
  wire   [1:0] cell_1731_and_in;
  wire   [1:0] cell_1731_a_HPC2_and_a_reg;
  wire   [1:0] cell_1731_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1731_a_HPC2_and_mul;
  wire   [1:0] cell_1732_and_out;
  wire   [1:0] cell_1732_and_in;
  wire   [1:0] cell_1732_a_HPC2_and_a_reg;
  wire   [1:0] cell_1732_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1732_a_HPC2_and_mul;
  wire   [1:0] cell_1733_and_out;
  wire   [1:0] cell_1733_and_in;
  wire   [1:0] cell_1733_a_HPC2_and_a_reg;
  wire   [1:0] cell_1733_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1733_a_HPC2_and_mul;
  wire   [1:0] cell_1734_and_out;
  wire   [1:0] cell_1734_and_in;
  wire   [1:0] cell_1734_a_HPC2_and_a_reg;
  wire   [1:0] cell_1734_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1734_a_HPC2_and_mul;
  wire   [1:0] cell_1735_and_out;
  wire   [1:0] cell_1735_and_in;
  wire   [1:0] cell_1735_a_HPC2_and_a_reg;
  wire   [1:0] cell_1735_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1735_a_HPC2_and_mul;
  wire   [1:0] cell_1736_and_out;
  wire   [1:0] cell_1736_and_in;
  wire   [1:0] cell_1736_a_HPC2_and_a_reg;
  wire   [1:0] cell_1736_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1736_a_HPC2_and_mul;
  wire   [1:0] cell_1737_and_out;
  wire   [1:0] cell_1737_and_in;
  wire   [1:0] cell_1737_a_HPC2_and_a_reg;
  wire   [1:0] cell_1737_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1737_a_HPC2_and_mul;
  wire   [1:0] cell_1738_and_out;
  wire   [1:0] cell_1738_and_in;
  wire   [1:0] cell_1738_a_HPC2_and_a_reg;
  wire   [1:0] cell_1738_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1738_a_HPC2_and_mul;
  wire   [1:0] cell_1739_and_out;
  wire   [1:0] cell_1739_and_in;
  wire   [1:0] cell_1739_a_HPC2_and_a_reg;
  wire   [1:0] cell_1739_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1739_a_HPC2_and_mul;
  wire   [1:0] cell_1740_and_out;
  wire   [1:0] cell_1740_and_in;
  wire   [1:0] cell_1740_a_HPC2_and_a_reg;
  wire   [1:0] cell_1740_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1740_a_HPC2_and_mul;
  wire   [1:0] cell_1741_and_out;
  wire   [1:0] cell_1741_and_in;
  wire   [1:0] cell_1741_a_HPC2_and_a_reg;
  wire   [1:0] cell_1741_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1741_a_HPC2_and_mul;
  wire   [1:0] cell_1742_and_out;
  wire   [1:0] cell_1742_and_in;
  wire   [1:0] cell_1742_a_HPC2_and_a_reg;
  wire   [1:0] cell_1742_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1742_a_HPC2_and_mul;
  wire   [1:0] cell_1743_and_out;
  wire   [1:0] cell_1743_and_in;
  wire   [1:0] cell_1743_a_HPC2_and_a_reg;
  wire   [1:0] cell_1743_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1743_a_HPC2_and_mul;
  wire   [1:0] cell_1744_and_out;
  wire   [1:0] cell_1744_and_in;
  wire   [1:0] cell_1744_a_HPC2_and_a_reg;
  wire   [1:0] cell_1744_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1744_a_HPC2_and_mul;
  wire   [1:0] cell_1745_and_out;
  wire   [1:0] cell_1745_and_in;
  wire   [1:0] cell_1745_a_HPC2_and_a_reg;
  wire   [1:0] cell_1745_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1745_a_HPC2_and_mul;
  wire   [1:0] cell_1746_and_out;
  wire   [1:0] cell_1746_and_in;
  wire   [1:0] cell_1746_a_HPC2_and_a_reg;
  wire   [1:0] cell_1746_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1746_a_HPC2_and_mul;
  wire   [1:0] cell_1747_and_out;
  wire   [1:0] cell_1747_and_in;
  wire   [1:0] cell_1747_a_HPC2_and_a_reg;
  wire   [1:0] cell_1747_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1747_a_HPC2_and_mul;
  wire   [1:0] cell_1748_and_out;
  wire   [1:0] cell_1748_and_in;
  wire   [1:0] cell_1748_a_HPC2_and_a_reg;
  wire   [1:0] cell_1748_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1748_a_HPC2_and_mul;
  wire   [1:0] cell_1749_and_out;
  wire   [1:0] cell_1749_and_in;
  wire   [1:0] cell_1749_a_HPC2_and_a_reg;
  wire   [1:0] cell_1749_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1749_a_HPC2_and_mul;
  wire   [1:0] cell_1750_and_out;
  wire   [1:0] cell_1750_and_in;
  wire   [1:0] cell_1750_a_HPC2_and_a_reg;
  wire   [1:0] cell_1750_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1750_a_HPC2_and_mul;
  wire   [1:0] cell_1751_and_out;
  wire   [1:0] cell_1751_and_in;
  wire   [1:0] cell_1751_a_HPC2_and_a_reg;
  wire   [1:0] cell_1751_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1751_a_HPC2_and_mul;
  wire   [1:0] cell_1752_and_out;
  wire   [1:0] cell_1752_and_in;
  wire   [1:0] cell_1752_a_HPC2_and_a_reg;
  wire   [1:0] cell_1752_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1752_a_HPC2_and_mul;
  wire   [1:0] cell_1753_and_out;
  wire   [1:0] cell_1753_and_in;
  wire   [1:0] cell_1753_a_HPC2_and_a_reg;
  wire   [1:0] cell_1753_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1753_a_HPC2_and_mul;
  wire   [1:0] cell_1754_and_out;
  wire   [1:0] cell_1754_and_in;
  wire   [1:0] cell_1754_a_HPC2_and_a_reg;
  wire   [1:0] cell_1754_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1754_a_HPC2_and_mul;
  wire   [1:0] cell_1755_and_out;
  wire   [1:0] cell_1755_and_in;
  wire   [1:0] cell_1755_a_HPC2_and_a_reg;
  wire   [1:0] cell_1755_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1755_a_HPC2_and_mul;
  wire   [1:0] cell_1756_and_out;
  wire   [1:0] cell_1756_and_in;
  wire   [1:0] cell_1756_a_HPC2_and_a_reg;
  wire   [1:0] cell_1756_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1756_a_HPC2_and_mul;
  wire   [1:0] cell_1757_and_out;
  wire   [1:0] cell_1757_and_in;
  wire   [1:0] cell_1757_a_HPC2_and_a_reg;
  wire   [1:0] cell_1757_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1757_a_HPC2_and_mul;
  wire   [1:0] cell_1758_and_out;
  wire   [1:0] cell_1758_and_in;
  wire   [1:0] cell_1758_a_HPC2_and_a_reg;
  wire   [1:0] cell_1758_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1758_a_HPC2_and_mul;
  wire   [1:0] cell_1759_and_out;
  wire   [1:0] cell_1759_and_in;
  wire   [1:0] cell_1759_a_HPC2_and_a_reg;
  wire   [1:0] cell_1759_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1759_a_HPC2_and_mul;
  wire   [1:0] cell_1760_and_out;
  wire   [1:0] cell_1760_and_in;
  wire   [1:0] cell_1760_a_HPC2_and_a_reg;
  wire   [1:0] cell_1760_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1760_a_HPC2_and_mul;
  wire   [1:0] cell_1761_and_out;
  wire   [1:0] cell_1761_and_in;
  wire   [1:0] cell_1761_a_HPC2_and_a_reg;
  wire   [1:0] cell_1761_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1761_a_HPC2_and_mul;
  wire   [1:0] cell_1762_and_out;
  wire   [1:0] cell_1762_and_in;
  wire   [1:0] cell_1762_a_HPC2_and_a_reg;
  wire   [1:0] cell_1762_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1762_a_HPC2_and_mul;
  wire   [1:0] cell_1763_and_out;
  wire   [1:0] cell_1763_and_in;
  wire   [1:0] cell_1763_a_HPC2_and_a_reg;
  wire   [1:0] cell_1763_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1763_a_HPC2_and_mul;
  wire   [1:0] cell_1764_and_out;
  wire   [1:0] cell_1764_and_in;
  wire   [1:0] cell_1764_a_HPC2_and_a_reg;
  wire   [1:0] cell_1764_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1764_a_HPC2_and_mul;
  wire   [1:0] cell_1765_and_out;
  wire   [1:0] cell_1765_and_in;
  wire   [1:0] cell_1765_a_HPC2_and_a_reg;
  wire   [1:0] cell_1765_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1765_a_HPC2_and_mul;
  wire   [1:0] cell_1766_and_out;
  wire   [1:0] cell_1766_and_in;
  wire   [1:0] cell_1766_a_HPC2_and_a_reg;
  wire   [1:0] cell_1766_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1766_a_HPC2_and_mul;
  wire   [1:0] cell_1767_and_out;
  wire   [1:0] cell_1767_and_in;
  wire   [1:0] cell_1767_a_HPC2_and_a_reg;
  wire   [1:0] cell_1767_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1767_a_HPC2_and_mul;
  wire   [1:0] cell_1768_and_out;
  wire   [1:0] cell_1768_and_in;
  wire   [1:0] cell_1768_a_HPC2_and_a_reg;
  wire   [1:0] cell_1768_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1768_a_HPC2_and_mul;
  wire   [1:0] cell_1769_and_out;
  wire   [1:0] cell_1769_and_in;
  wire   [1:0] cell_1769_a_HPC2_and_a_reg;
  wire   [1:0] cell_1769_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1769_a_HPC2_and_mul;
  wire   [1:0] cell_1770_and_out;
  wire   [1:0] cell_1770_and_in;
  wire   [1:0] cell_1770_a_HPC2_and_a_reg;
  wire   [1:0] cell_1770_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1770_a_HPC2_and_mul;
  wire   [1:0] cell_1771_and_out;
  wire   [1:0] cell_1771_and_in;
  wire   [1:0] cell_1771_a_HPC2_and_a_reg;
  wire   [1:0] cell_1771_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1771_a_HPC2_and_mul;
  wire   [1:0] cell_1772_and_out;
  wire   [1:0] cell_1772_and_in;
  wire   [1:0] cell_1772_a_HPC2_and_a_reg;
  wire   [1:0] cell_1772_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1772_a_HPC2_and_mul;
  wire   [1:0] cell_1773_and_out;
  wire   [1:0] cell_1773_and_in;
  wire   [1:0] cell_1773_a_HPC2_and_a_reg;
  wire   [1:0] cell_1773_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1773_a_HPC2_and_mul;
  wire   [1:0] cell_1774_and_out;
  wire   [1:0] cell_1774_and_in;
  wire   [1:0] cell_1774_a_HPC2_and_a_reg;
  wire   [1:0] cell_1774_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1774_a_HPC2_and_mul;
  wire   [1:0] cell_1775_and_out;
  wire   [1:0] cell_1775_and_in;
  wire   [1:0] cell_1775_a_HPC2_and_a_reg;
  wire   [1:0] cell_1775_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1775_a_HPC2_and_mul;
  wire   [1:0] cell_1776_and_out;
  wire   [1:0] cell_1776_and_in;
  wire   [1:0] cell_1776_a_HPC2_and_a_reg;
  wire   [1:0] cell_1776_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1776_a_HPC2_and_mul;
  wire   [1:0] cell_1777_and_out;
  wire   [1:0] cell_1777_and_in;
  wire   [1:0] cell_1777_a_HPC2_and_a_reg;
  wire   [1:0] cell_1777_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1777_a_HPC2_and_mul;
  wire   [1:0] cell_1778_and_out;
  wire   [1:0] cell_1778_and_in;
  wire   [1:0] cell_1778_a_HPC2_and_a_reg;
  wire   [1:0] cell_1778_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1778_a_HPC2_and_mul;
  wire   [1:0] cell_1779_and_out;
  wire   [1:0] cell_1779_and_in;
  wire   [1:0] cell_1779_a_HPC2_and_a_reg;
  wire   [1:0] cell_1779_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1779_a_HPC2_and_mul;
  wire   [1:0] cell_1780_and_out;
  wire   [1:0] cell_1780_and_in;
  wire   [1:0] cell_1780_a_HPC2_and_a_reg;
  wire   [1:0] cell_1780_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1780_a_HPC2_and_mul;
  wire   [1:0] cell_1781_and_out;
  wire   [1:0] cell_1781_and_in;
  wire   [1:0] cell_1781_a_HPC2_and_a_reg;
  wire   [1:0] cell_1781_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1781_a_HPC2_and_mul;
  wire   [1:0] cell_1782_and_out;
  wire   [1:0] cell_1782_and_in;
  wire   [1:0] cell_1782_a_HPC2_and_a_reg;
  wire   [1:0] cell_1782_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1782_a_HPC2_and_mul;
  wire   [1:0] cell_1783_and_out;
  wire   [1:0] cell_1783_and_in;
  wire   [1:0] cell_1783_a_HPC2_and_a_reg;
  wire   [1:0] cell_1783_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1783_a_HPC2_and_mul;
  wire   [1:0] cell_1784_and_out;
  wire   [1:0] cell_1784_and_in;
  wire   [1:0] cell_1784_a_HPC2_and_a_reg;
  wire   [1:0] cell_1784_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1784_a_HPC2_and_mul;
  wire   [1:0] cell_1785_and_out;
  wire   [1:0] cell_1785_and_in;
  wire   [1:0] cell_1785_a_HPC2_and_a_reg;
  wire   [1:0] cell_1785_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1785_a_HPC2_and_mul;
  wire   [1:0] cell_1786_and_out;
  wire   [1:0] cell_1786_and_in;
  wire   [1:0] cell_1786_a_HPC2_and_a_reg;
  wire   [1:0] cell_1786_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1786_a_HPC2_and_mul;
  wire   [1:0] cell_1787_and_out;
  wire   [1:0] cell_1787_and_in;
  wire   [1:0] cell_1787_a_HPC2_and_a_reg;
  wire   [1:0] cell_1787_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1787_a_HPC2_and_mul;
  wire   [1:0] cell_1788_and_out;
  wire   [1:0] cell_1788_and_in;
  wire   [1:0] cell_1788_a_HPC2_and_a_reg;
  wire   [1:0] cell_1788_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1788_a_HPC2_and_mul;
  wire   [1:0] cell_1789_and_out;
  wire   [1:0] cell_1789_and_in;
  wire   [1:0] cell_1789_a_HPC2_and_a_reg;
  wire   [1:0] cell_1789_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1789_a_HPC2_and_mul;
  wire   [1:0] cell_1790_and_out;
  wire   [1:0] cell_1790_and_in;
  wire   [1:0] cell_1790_a_HPC2_and_a_reg;
  wire   [1:0] cell_1790_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1790_a_HPC2_and_mul;
  wire   [1:0] cell_1791_and_out;
  wire   [1:0] cell_1791_and_in;
  wire   [1:0] cell_1791_a_HPC2_and_a_reg;
  wire   [1:0] cell_1791_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1791_a_HPC2_and_mul;
  wire   [1:0] cell_1792_and_out;
  wire   [1:0] cell_1792_and_in;
  wire   [1:0] cell_1792_a_HPC2_and_a_reg;
  wire   [1:0] cell_1792_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1792_a_HPC2_and_mul;
  wire   [1:0] cell_1793_and_out;
  wire   [1:0] cell_1793_and_in;
  wire   [1:0] cell_1793_a_HPC2_and_a_reg;
  wire   [1:0] cell_1793_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1793_a_HPC2_and_mul;
  wire   [1:0] cell_1794_and_out;
  wire   [1:0] cell_1794_and_in;
  wire   [1:0] cell_1794_a_HPC2_and_a_reg;
  wire   [1:0] cell_1794_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1794_a_HPC2_and_mul;
  wire   [1:0] cell_1795_and_out;
  wire   [1:0] cell_1795_and_in;
  wire   [1:0] cell_1795_a_HPC2_and_a_reg;
  wire   [1:0] cell_1795_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1795_a_HPC2_and_mul;
  wire   [1:0] cell_1796_and_out;
  wire   [1:0] cell_1796_and_in;
  wire   [1:0] cell_1796_a_HPC2_and_a_reg;
  wire   [1:0] cell_1796_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1796_a_HPC2_and_mul;
  wire   [1:0] cell_1797_and_out;
  wire   [1:0] cell_1797_and_in;
  wire   [1:0] cell_1797_a_HPC2_and_a_reg;
  wire   [1:0] cell_1797_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1797_a_HPC2_and_mul;
  wire   [1:0] cell_1798_and_out;
  wire   [1:0] cell_1798_and_in;
  wire   [1:0] cell_1798_a_HPC2_and_a_reg;
  wire   [1:0] cell_1798_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1798_a_HPC2_and_mul;
  wire   [1:0] cell_1799_and_out;
  wire   [1:0] cell_1799_and_in;
  wire   [1:0] cell_1799_a_HPC2_and_a_reg;
  wire   [1:0] cell_1799_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1799_a_HPC2_and_mul;
  wire   [1:0] cell_1800_and_out;
  wire   [1:0] cell_1800_and_in;
  wire   [1:0] cell_1800_a_HPC2_and_a_reg;
  wire   [1:0] cell_1800_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1800_a_HPC2_and_mul;
  wire   [1:0] cell_1801_and_out;
  wire   [1:0] cell_1801_and_in;
  wire   [1:0] cell_1801_a_HPC2_and_a_reg;
  wire   [1:0] cell_1801_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1801_a_HPC2_and_mul;
  wire   [1:0] cell_1802_and_out;
  wire   [1:0] cell_1802_and_in;
  wire   [1:0] cell_1802_a_HPC2_and_a_reg;
  wire   [1:0] cell_1802_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1802_a_HPC2_and_mul;
  wire   [1:0] cell_1803_and_out;
  wire   [1:0] cell_1803_and_in;
  wire   [1:0] cell_1803_a_HPC2_and_a_reg;
  wire   [1:0] cell_1803_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1803_a_HPC2_and_mul;
  wire   [1:0] cell_1804_and_out;
  wire   [1:0] cell_1804_and_in;
  wire   [1:0] cell_1804_a_HPC2_and_a_reg;
  wire   [1:0] cell_1804_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1804_a_HPC2_and_mul;
  wire   [1:0] cell_1805_and_out;
  wire   [1:0] cell_1805_and_in;
  wire   [1:0] cell_1805_a_HPC2_and_a_reg;
  wire   [1:0] cell_1805_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1805_a_HPC2_and_mul;
  wire   [1:0] cell_1806_and_out;
  wire   [1:0] cell_1806_and_in;
  wire   [1:0] cell_1806_a_HPC2_and_a_reg;
  wire   [1:0] cell_1806_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1806_a_HPC2_and_mul;
  wire   [1:0] cell_1807_and_out;
  wire   [1:0] cell_1807_and_in;
  wire   [1:0] cell_1807_a_HPC2_and_a_reg;
  wire   [1:0] cell_1807_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1807_a_HPC2_and_mul;
  wire   [1:0] cell_1808_and_out;
  wire   [1:0] cell_1808_and_in;
  wire   [1:0] cell_1808_a_HPC2_and_a_reg;
  wire   [1:0] cell_1808_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1808_a_HPC2_and_mul;
  wire   [1:0] cell_1809_and_out;
  wire   [1:0] cell_1809_and_in;
  wire   [1:0] cell_1809_a_HPC2_and_a_reg;
  wire   [1:0] cell_1809_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1809_a_HPC2_and_mul;
  wire   [1:0] cell_1810_and_out;
  wire   [1:0] cell_1810_and_in;
  wire   [1:0] cell_1810_a_HPC2_and_a_reg;
  wire   [1:0] cell_1810_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1810_a_HPC2_and_mul;
  wire   [1:0] cell_1811_and_out;
  wire   [1:0] cell_1811_and_in;
  wire   [1:0] cell_1811_a_HPC2_and_a_reg;
  wire   [1:0] cell_1811_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1811_a_HPC2_and_mul;
  wire   [1:0] cell_1812_and_out;
  wire   [1:0] cell_1812_and_in;
  wire   [1:0] cell_1812_a_HPC2_and_a_reg;
  wire   [1:0] cell_1812_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1812_a_HPC2_and_mul;
  wire   [1:0] cell_1813_and_out;
  wire   [1:0] cell_1813_and_in;
  wire   [1:0] cell_1813_a_HPC2_and_a_reg;
  wire   [1:0] cell_1813_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1813_a_HPC2_and_mul;
  wire   [1:0] cell_1814_and_out;
  wire   [1:0] cell_1814_and_in;
  wire   [1:0] cell_1814_a_HPC2_and_a_reg;
  wire   [1:0] cell_1814_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1814_a_HPC2_and_mul;
  wire   [1:0] cell_1815_and_out;
  wire   [1:0] cell_1815_and_in;
  wire   [1:0] cell_1815_a_HPC2_and_a_reg;
  wire   [1:0] cell_1815_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1815_a_HPC2_and_mul;
  wire   [1:0] cell_1816_and_out;
  wire   [1:0] cell_1816_and_in;
  wire   [1:0] cell_1816_a_HPC2_and_a_reg;
  wire   [1:0] cell_1816_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1816_a_HPC2_and_mul;
  wire   [1:0] cell_1817_and_out;
  wire   [1:0] cell_1817_and_in;
  wire   [1:0] cell_1817_a_HPC2_and_a_reg;
  wire   [1:0] cell_1817_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1817_a_HPC2_and_mul;
  wire   [1:0] cell_1818_and_out;
  wire   [1:0] cell_1818_and_in;
  wire   [1:0] cell_1818_a_HPC2_and_a_reg;
  wire   [1:0] cell_1818_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1818_a_HPC2_and_mul;
  wire   [1:0] cell_1819_and_out;
  wire   [1:0] cell_1819_and_in;
  wire   [1:0] cell_1819_a_HPC2_and_a_reg;
  wire   [1:0] cell_1819_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1819_a_HPC2_and_mul;
  wire   [1:0] cell_1820_and_out;
  wire   [1:0] cell_1820_and_in;
  wire   [1:0] cell_1820_a_HPC2_and_a_reg;
  wire   [1:0] cell_1820_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1820_a_HPC2_and_mul;
  wire   [1:0] cell_1821_and_out;
  wire   [1:0] cell_1821_and_in;
  wire   [1:0] cell_1821_a_HPC2_and_a_reg;
  wire   [1:0] cell_1821_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1821_a_HPC2_and_mul;
  wire   [1:0] cell_1822_and_out;
  wire   [1:0] cell_1822_and_in;
  wire   [1:0] cell_1822_a_HPC2_and_a_reg;
  wire   [1:0] cell_1822_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1822_a_HPC2_and_mul;
  wire   [1:0] cell_1823_and_out;
  wire   [1:0] cell_1823_and_in;
  wire   [1:0] cell_1823_a_HPC2_and_a_reg;
  wire   [1:0] cell_1823_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1823_a_HPC2_and_mul;
  wire   [1:0] cell_1824_and_out;
  wire   [1:0] cell_1824_and_in;
  wire   [1:0] cell_1824_a_HPC2_and_a_reg;
  wire   [1:0] cell_1824_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1824_a_HPC2_and_mul;
  wire   [1:0] cell_1825_and_out;
  wire   [1:0] cell_1825_and_in;
  wire   [1:0] cell_1825_a_HPC2_and_a_reg;
  wire   [1:0] cell_1825_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1825_a_HPC2_and_mul;
  wire   [1:0] cell_1826_and_out;
  wire   [1:0] cell_1826_and_in;
  wire   [1:0] cell_1826_a_HPC2_and_a_reg;
  wire   [1:0] cell_1826_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1826_a_HPC2_and_mul;
  wire   [1:0] cell_1827_and_out;
  wire   [1:0] cell_1827_and_in;
  wire   [1:0] cell_1827_a_HPC2_and_a_reg;
  wire   [1:0] cell_1827_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1827_a_HPC2_and_mul;
  wire   [1:0] cell_1828_and_out;
  wire   [1:0] cell_1828_and_in;
  wire   [1:0] cell_1828_a_HPC2_and_a_reg;
  wire   [1:0] cell_1828_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1828_a_HPC2_and_mul;
  wire   [1:0] cell_1829_and_out;
  wire   [1:0] cell_1829_and_in;
  wire   [1:0] cell_1829_a_HPC2_and_a_reg;
  wire   [1:0] cell_1829_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1829_a_HPC2_and_mul;
  wire   [1:0] cell_1830_and_out;
  wire   [1:0] cell_1830_and_in;
  wire   [1:0] cell_1830_a_HPC2_and_a_reg;
  wire   [1:0] cell_1830_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1830_a_HPC2_and_mul;
  wire   [1:0] cell_1831_and_out;
  wire   [1:0] cell_1831_and_in;
  wire   [1:0] cell_1831_a_HPC2_and_a_reg;
  wire   [1:0] cell_1831_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1831_a_HPC2_and_mul;
  wire   [1:0] cell_1832_and_out;
  wire   [1:0] cell_1832_and_in;
  wire   [1:0] cell_1832_a_HPC2_and_a_reg;
  wire   [1:0] cell_1832_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1832_a_HPC2_and_mul;
  wire   [1:0] cell_1833_and_out;
  wire   [1:0] cell_1833_and_in;
  wire   [1:0] cell_1833_a_HPC2_and_a_reg;
  wire   [1:0] cell_1833_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1833_a_HPC2_and_mul;
  wire   [1:0] cell_1834_and_out;
  wire   [1:0] cell_1834_and_in;
  wire   [1:0] cell_1834_a_HPC2_and_a_reg;
  wire   [1:0] cell_1834_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1834_a_HPC2_and_mul;
  wire   [1:0] cell_1835_and_out;
  wire   [1:0] cell_1835_and_in;
  wire   [1:0] cell_1835_a_HPC2_and_a_reg;
  wire   [1:0] cell_1835_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1835_a_HPC2_and_mul;
  wire   [1:0] cell_1836_and_out;
  wire   [1:0] cell_1836_and_in;
  wire   [1:0] cell_1836_a_HPC2_and_a_reg;
  wire   [1:0] cell_1836_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1836_a_HPC2_and_mul;
  wire   [1:0] cell_1837_and_out;
  wire   [1:0] cell_1837_and_in;
  wire   [1:0] cell_1837_a_HPC2_and_a_reg;
  wire   [1:0] cell_1837_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1837_a_HPC2_and_mul;
  wire   [1:0] cell_1838_and_out;
  wire   [1:0] cell_1838_and_in;
  wire   [1:0] cell_1838_a_HPC2_and_a_reg;
  wire   [1:0] cell_1838_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1838_a_HPC2_and_mul;
  wire   [1:0] cell_1839_and_out;
  wire   [1:0] cell_1839_and_in;
  wire   [1:0] cell_1839_a_HPC2_and_a_reg;
  wire   [1:0] cell_1839_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1839_a_HPC2_and_mul;
  wire   [1:0] cell_1840_and_out;
  wire   [1:0] cell_1840_and_in;
  wire   [1:0] cell_1840_a_HPC2_and_a_reg;
  wire   [1:0] cell_1840_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1840_a_HPC2_and_mul;
  wire   [1:0] cell_1841_and_out;
  wire   [1:0] cell_1841_and_in;
  wire   [1:0] cell_1841_a_HPC2_and_a_reg;
  wire   [1:0] cell_1841_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1841_a_HPC2_and_mul;
  wire   [1:0] cell_1842_and_out;
  wire   [1:0] cell_1842_and_in;
  wire   [1:0] cell_1842_a_HPC2_and_a_reg;
  wire   [1:0] cell_1842_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1842_a_HPC2_and_mul;
  wire   [1:0] cell_1843_and_out;
  wire   [1:0] cell_1843_and_in;
  wire   [1:0] cell_1843_a_HPC2_and_a_reg;
  wire   [1:0] cell_1843_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1843_a_HPC2_and_mul;
  wire   [1:0] cell_1844_and_out;
  wire   [1:0] cell_1844_and_in;
  wire   [1:0] cell_1844_a_HPC2_and_a_reg;
  wire   [1:0] cell_1844_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1844_a_HPC2_and_mul;
  wire   [1:0] cell_1845_and_out;
  wire   [1:0] cell_1845_and_in;
  wire   [1:0] cell_1845_a_HPC2_and_a_reg;
  wire   [1:0] cell_1845_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1845_a_HPC2_and_mul;
  wire   [1:0] cell_1846_and_out;
  wire   [1:0] cell_1846_and_in;
  wire   [1:0] cell_1846_a_HPC2_and_a_reg;
  wire   [1:0] cell_1846_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1846_a_HPC2_and_mul;
  wire   [1:0] cell_1847_and_out;
  wire   [1:0] cell_1847_and_in;
  wire   [1:0] cell_1847_a_HPC2_and_a_reg;
  wire   [1:0] cell_1847_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1847_a_HPC2_and_mul;
  wire   [1:0] cell_1848_and_out;
  wire   [1:0] cell_1848_and_in;
  wire   [1:0] cell_1848_a_HPC2_and_a_reg;
  wire   [1:0] cell_1848_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1848_a_HPC2_and_mul;
  wire   [1:0] cell_1849_and_out;
  wire   [1:0] cell_1849_and_in;
  wire   [1:0] cell_1849_a_HPC2_and_a_reg;
  wire   [1:0] cell_1849_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1849_a_HPC2_and_mul;
  wire   [1:0] cell_1850_and_out;
  wire   [1:0] cell_1850_and_in;
  wire   [1:0] cell_1850_a_HPC2_and_a_reg;
  wire   [1:0] cell_1850_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1850_a_HPC2_and_mul;
  wire   [1:0] cell_1851_and_out;
  wire   [1:0] cell_1851_and_in;
  wire   [1:0] cell_1851_a_HPC2_and_a_reg;
  wire   [1:0] cell_1851_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1851_a_HPC2_and_mul;
  wire   [1:0] cell_1852_and_out;
  wire   [1:0] cell_1852_and_in;
  wire   [1:0] cell_1852_a_HPC2_and_a_reg;
  wire   [1:0] cell_1852_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1852_a_HPC2_and_mul;
  wire   [1:0] cell_1853_and_out;
  wire   [1:0] cell_1853_and_in;
  wire   [1:0] cell_1853_a_HPC2_and_a_reg;
  wire   [1:0] cell_1853_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1853_a_HPC2_and_mul;
  wire   [1:0] cell_1854_and_out;
  wire   [1:0] cell_1854_and_in;
  wire   [1:0] cell_1854_a_HPC2_and_a_reg;
  wire   [1:0] cell_1854_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1854_a_HPC2_and_mul;
  wire   [1:0] cell_1855_and_out;
  wire   [1:0] cell_1855_and_in;
  wire   [1:0] cell_1855_a_HPC2_and_a_reg;
  wire   [1:0] cell_1855_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1855_a_HPC2_and_mul;
  wire   [1:0] cell_1856_and_out;
  wire   [1:0] cell_1856_and_in;
  wire   [1:0] cell_1856_a_HPC2_and_a_reg;
  wire   [1:0] cell_1856_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1856_a_HPC2_and_mul;
  wire   [1:0] cell_1857_and_out;
  wire   [1:0] cell_1857_and_in;
  wire   [1:0] cell_1857_a_HPC2_and_a_reg;
  wire   [1:0] cell_1857_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1857_a_HPC2_and_mul;
  wire   [1:0] cell_1858_and_out;
  wire   [1:0] cell_1858_and_in;
  wire   [1:0] cell_1858_a_HPC2_and_a_reg;
  wire   [1:0] cell_1858_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1858_a_HPC2_and_mul;
  wire   [1:0] cell_1859_and_out;
  wire   [1:0] cell_1859_and_in;
  wire   [1:0] cell_1859_a_HPC2_and_a_reg;
  wire   [1:0] cell_1859_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1859_a_HPC2_and_mul;
  wire   [1:0] cell_1860_and_out;
  wire   [1:0] cell_1860_and_in;
  wire   [1:0] cell_1860_a_HPC2_and_a_reg;
  wire   [1:0] cell_1860_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1860_a_HPC2_and_mul;
  wire   [1:0] cell_1861_and_out;
  wire   [1:0] cell_1861_and_in;
  wire   [1:0] cell_1861_a_HPC2_and_a_reg;
  wire   [1:0] cell_1861_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1861_a_HPC2_and_mul;
  wire   [1:0] cell_1862_and_out;
  wire   [1:0] cell_1862_and_in;
  wire   [1:0] cell_1862_a_HPC2_and_a_reg;
  wire   [1:0] cell_1862_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1862_a_HPC2_and_mul;
  wire   [1:0] cell_1863_and_out;
  wire   [1:0] cell_1863_and_in;
  wire   [1:0] cell_1863_a_HPC2_and_a_reg;
  wire   [1:0] cell_1863_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1863_a_HPC2_and_mul;
  wire   [1:0] cell_1864_and_out;
  wire   [1:0] cell_1864_and_in;
  wire   [1:0] cell_1864_a_HPC2_and_a_reg;
  wire   [1:0] cell_1864_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1864_a_HPC2_and_mul;
  wire   [1:0] cell_1865_and_out;
  wire   [1:0] cell_1865_and_in;
  wire   [1:0] cell_1865_a_HPC2_and_a_reg;
  wire   [1:0] cell_1865_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1865_a_HPC2_and_mul;
  wire   [1:0] cell_1866_and_out;
  wire   [1:0] cell_1866_and_in;
  wire   [1:0] cell_1866_a_HPC2_and_a_reg;
  wire   [1:0] cell_1866_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1866_a_HPC2_and_mul;
  wire   [1:0] cell_1867_and_out;
  wire   [1:0] cell_1867_and_in;
  wire   [1:0] cell_1867_a_HPC2_and_a_reg;
  wire   [1:0] cell_1867_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1867_a_HPC2_and_mul;
  wire   [1:0] cell_1868_and_out;
  wire   [1:0] cell_1868_and_in;
  wire   [1:0] cell_1868_a_HPC2_and_a_reg;
  wire   [1:0] cell_1868_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1868_a_HPC2_and_mul;
  wire   [1:0] cell_1869_and_out;
  wire   [1:0] cell_1869_and_in;
  wire   [1:0] cell_1869_a_HPC2_and_a_reg;
  wire   [1:0] cell_1869_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1869_a_HPC2_and_mul;
  wire   [1:0] cell_1870_and_out;
  wire   [1:0] cell_1870_and_in;
  wire   [1:0] cell_1870_a_HPC2_and_a_reg;
  wire   [1:0] cell_1870_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1870_a_HPC2_and_mul;
  wire   [1:0] cell_1871_and_out;
  wire   [1:0] cell_1871_and_in;
  wire   [1:0] cell_1871_a_HPC2_and_a_reg;
  wire   [1:0] cell_1871_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1871_a_HPC2_and_mul;
  wire   [1:0] cell_1872_and_out;
  wire   [1:0] cell_1872_and_in;
  wire   [1:0] cell_1872_a_HPC2_and_a_reg;
  wire   [1:0] cell_1872_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1872_a_HPC2_and_mul;
  wire   [1:0] cell_1873_and_out;
  wire   [1:0] cell_1873_and_in;
  wire   [1:0] cell_1873_a_HPC2_and_a_reg;
  wire   [1:0] cell_1873_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1873_a_HPC2_and_mul;
  wire   [1:0] cell_1874_and_out;
  wire   [1:0] cell_1874_and_in;
  wire   [1:0] cell_1874_a_HPC2_and_a_reg;
  wire   [1:0] cell_1874_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1874_a_HPC2_and_mul;
  wire   [1:0] cell_1875_and_out;
  wire   [1:0] cell_1875_and_in;
  wire   [1:0] cell_1875_a_HPC2_and_a_reg;
  wire   [1:0] cell_1875_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1875_a_HPC2_and_mul;
  wire   [1:0] cell_1876_and_out;
  wire   [1:0] cell_1876_and_in;
  wire   [1:0] cell_1876_a_HPC2_and_a_reg;
  wire   [1:0] cell_1876_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1876_a_HPC2_and_mul;
  wire   [1:0] cell_1877_and_out;
  wire   [1:0] cell_1877_and_in;
  wire   [1:0] cell_1877_a_HPC2_and_a_reg;
  wire   [1:0] cell_1877_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1877_a_HPC2_and_mul;
  wire   [1:0] cell_1878_and_out;
  wire   [1:0] cell_1878_and_in;
  wire   [1:0] cell_1878_a_HPC2_and_a_reg;
  wire   [1:0] cell_1878_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1878_a_HPC2_and_mul;
  wire   [1:0] cell_1879_and_out;
  wire   [1:0] cell_1879_and_in;
  wire   [1:0] cell_1879_a_HPC2_and_a_reg;
  wire   [1:0] cell_1879_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1879_a_HPC2_and_mul;
  wire   [1:0] cell_1880_and_out;
  wire   [1:0] cell_1880_and_in;
  wire   [1:0] cell_1880_a_HPC2_and_a_reg;
  wire   [1:0] cell_1880_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1880_a_HPC2_and_mul;
  wire   [1:0] cell_1881_and_out;
  wire   [1:0] cell_1881_and_in;
  wire   [1:0] cell_1881_a_HPC2_and_a_reg;
  wire   [1:0] cell_1881_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1881_a_HPC2_and_mul;
  wire   [1:0] cell_1882_and_out;
  wire   [1:0] cell_1882_and_in;
  wire   [1:0] cell_1882_a_HPC2_and_a_reg;
  wire   [1:0] cell_1882_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1882_a_HPC2_and_mul;
  wire   [1:0] cell_1883_and_out;
  wire   [1:0] cell_1883_and_in;
  wire   [1:0] cell_1883_a_HPC2_and_a_reg;
  wire   [1:0] cell_1883_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1883_a_HPC2_and_mul;
  wire   [1:0] cell_1884_and_out;
  wire   [1:0] cell_1884_and_in;
  wire   [1:0] cell_1884_a_HPC2_and_a_reg;
  wire   [1:0] cell_1884_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1884_a_HPC2_and_mul;
  wire   [1:0] cell_1885_and_out;
  wire   [1:0] cell_1885_and_in;
  wire   [1:0] cell_1885_a_HPC2_and_a_reg;
  wire   [1:0] cell_1885_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1885_a_HPC2_and_mul;
  wire   [1:0] cell_1886_and_out;
  wire   [1:0] cell_1886_and_in;
  wire   [1:0] cell_1886_a_HPC2_and_a_reg;
  wire   [1:0] cell_1886_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1886_a_HPC2_and_mul;
  wire   [1:0] cell_1887_and_out;
  wire   [1:0] cell_1887_and_in;
  wire   [1:0] cell_1887_a_HPC2_and_a_reg;
  wire   [1:0] cell_1887_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1887_a_HPC2_and_mul;
  wire   [1:0] cell_1888_and_out;
  wire   [1:0] cell_1888_and_in;
  wire   [1:0] cell_1888_a_HPC2_and_a_reg;
  wire   [1:0] cell_1888_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1888_a_HPC2_and_mul;
  wire   [1:0] cell_1889_and_out;
  wire   [1:0] cell_1889_and_in;
  wire   [1:0] cell_1889_a_HPC2_and_a_reg;
  wire   [1:0] cell_1889_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1889_a_HPC2_and_mul;
  wire   [1:0] cell_1890_and_out;
  wire   [1:0] cell_1890_and_in;
  wire   [1:0] cell_1890_a_HPC2_and_a_reg;
  wire   [1:0] cell_1890_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1890_a_HPC2_and_mul;
  wire   [1:0] cell_1891_and_out;
  wire   [1:0] cell_1891_and_in;
  wire   [1:0] cell_1891_a_HPC2_and_a_reg;
  wire   [1:0] cell_1891_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1891_a_HPC2_and_mul;
  wire   [1:0] cell_1892_and_out;
  wire   [1:0] cell_1892_and_in;
  wire   [1:0] cell_1892_a_HPC2_and_a_reg;
  wire   [1:0] cell_1892_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1892_a_HPC2_and_mul;
  wire   [1:0] cell_1893_and_out;
  wire   [1:0] cell_1893_and_in;
  wire   [1:0] cell_1893_a_HPC2_and_a_reg;
  wire   [1:0] cell_1893_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1893_a_HPC2_and_mul;
  wire   [1:0] cell_1894_and_out;
  wire   [1:0] cell_1894_and_in;
  wire   [1:0] cell_1894_a_HPC2_and_a_reg;
  wire   [1:0] cell_1894_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1894_a_HPC2_and_mul;
  wire   [1:0] cell_1895_and_out;
  wire   [1:0] cell_1895_and_in;
  wire   [1:0] cell_1895_a_HPC2_and_a_reg;
  wire   [1:0] cell_1895_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1895_a_HPC2_and_mul;
  wire   [1:0] cell_1896_and_out;
  wire   [1:0] cell_1896_and_in;
  wire   [1:0] cell_1896_a_HPC2_and_a_reg;
  wire   [1:0] cell_1896_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1896_a_HPC2_and_mul;
  wire   [1:0] cell_1897_and_out;
  wire   [1:0] cell_1897_and_in;
  wire   [1:0] cell_1897_a_HPC2_and_a_reg;
  wire   [1:0] cell_1897_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1897_a_HPC2_and_mul;
  wire   [1:0] cell_1898_and_out;
  wire   [1:0] cell_1898_and_in;
  wire   [1:0] cell_1898_a_HPC2_and_a_reg;
  wire   [1:0] cell_1898_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1898_a_HPC2_and_mul;
  wire   [1:0] cell_1899_and_out;
  wire   [1:0] cell_1899_and_in;
  wire   [1:0] cell_1899_a_HPC2_and_a_reg;
  wire   [1:0] cell_1899_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1899_a_HPC2_and_mul;
  wire   [1:0] cell_1900_and_out;
  wire   [1:0] cell_1900_and_in;
  wire   [1:0] cell_1900_a_HPC2_and_a_reg;
  wire   [1:0] cell_1900_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1900_a_HPC2_and_mul;
  wire   [1:0] cell_1901_and_out;
  wire   [1:0] cell_1901_and_in;
  wire   [1:0] cell_1901_a_HPC2_and_a_reg;
  wire   [1:0] cell_1901_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1901_a_HPC2_and_mul;
  wire   [1:0] cell_1902_and_out;
  wire   [1:0] cell_1902_and_in;
  wire   [1:0] cell_1902_a_HPC2_and_a_reg;
  wire   [1:0] cell_1902_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1902_a_HPC2_and_mul;
  wire   [1:0] cell_1903_and_out;
  wire   [1:0] cell_1903_and_in;
  wire   [1:0] cell_1903_a_HPC2_and_a_reg;
  wire   [1:0] cell_1903_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1903_a_HPC2_and_mul;
  wire   [1:0] cell_1904_and_out;
  wire   [1:0] cell_1904_and_in;
  wire   [1:0] cell_1904_a_HPC2_and_a_reg;
  wire   [1:0] cell_1904_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1904_a_HPC2_and_mul;
  wire   [1:0] cell_1905_and_out;
  wire   [1:0] cell_1905_and_in;
  wire   [1:0] cell_1905_a_HPC2_and_a_reg;
  wire   [1:0] cell_1905_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1905_a_HPC2_and_mul;
  wire   [1:0] cell_1906_and_out;
  wire   [1:0] cell_1906_and_in;
  wire   [1:0] cell_1906_a_HPC2_and_a_reg;
  wire   [1:0] cell_1906_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1906_a_HPC2_and_mul;
  wire   [1:0] cell_1907_and_out;
  wire   [1:0] cell_1907_and_in;
  wire   [1:0] cell_1907_a_HPC2_and_a_reg;
  wire   [1:0] cell_1907_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1907_a_HPC2_and_mul;
  wire   [1:0] cell_1908_and_out;
  wire   [1:0] cell_1908_and_in;
  wire   [1:0] cell_1908_a_HPC2_and_a_reg;
  wire   [1:0] cell_1908_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1908_a_HPC2_and_mul;
  wire   [1:0] cell_1909_and_out;
  wire   [1:0] cell_1909_and_in;
  wire   [1:0] cell_1909_a_HPC2_and_a_reg;
  wire   [1:0] cell_1909_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1909_a_HPC2_and_mul;
  wire   [1:0] cell_1910_and_out;
  wire   [1:0] cell_1910_and_in;
  wire   [1:0] cell_1910_a_HPC2_and_a_reg;
  wire   [1:0] cell_1910_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1910_a_HPC2_and_mul;
  wire   [1:0] cell_1911_and_out;
  wire   [1:0] cell_1911_and_in;
  wire   [1:0] cell_1911_a_HPC2_and_a_reg;
  wire   [1:0] cell_1911_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1911_a_HPC2_and_mul;
  wire   [1:0] cell_1912_and_out;
  wire   [1:0] cell_1912_and_in;
  wire   [1:0] cell_1912_a_HPC2_and_a_reg;
  wire   [1:0] cell_1912_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1912_a_HPC2_and_mul;
  wire   [1:0] cell_1913_and_out;
  wire   [1:0] cell_1913_and_in;
  wire   [1:0] cell_1913_a_HPC2_and_a_reg;
  wire   [1:0] cell_1913_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1913_a_HPC2_and_mul;
  wire   [1:0] cell_1914_and_out;
  wire   [1:0] cell_1914_and_in;
  wire   [1:0] cell_1914_a_HPC2_and_a_reg;
  wire   [1:0] cell_1914_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1914_a_HPC2_and_mul;
  wire   [1:0] cell_1915_and_out;
  wire   [1:0] cell_1915_and_in;
  wire   [1:0] cell_1915_a_HPC2_and_a_reg;
  wire   [1:0] cell_1915_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1915_a_HPC2_and_mul;
  wire   [1:0] cell_1916_and_out;
  wire   [1:0] cell_1916_and_in;
  wire   [1:0] cell_1916_a_HPC2_and_a_reg;
  wire   [1:0] cell_1916_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1916_a_HPC2_and_mul;
  wire   [1:0] cell_1917_and_out;
  wire   [1:0] cell_1917_and_in;
  wire   [1:0] cell_1917_a_HPC2_and_a_reg;
  wire   [1:0] cell_1917_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1917_a_HPC2_and_mul;
  wire   [1:0] cell_1918_and_out;
  wire   [1:0] cell_1918_and_in;
  wire   [1:0] cell_1918_a_HPC2_and_a_reg;
  wire   [1:0] cell_1918_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1918_a_HPC2_and_mul;
  wire   [1:0] cell_1919_and_out;
  wire   [1:0] cell_1919_and_in;
  wire   [1:0] cell_1919_a_HPC2_and_a_reg;
  wire   [1:0] cell_1919_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1919_a_HPC2_and_mul;
  wire   [1:0] cell_1920_and_out;
  wire   [1:0] cell_1920_and_in;
  wire   [1:0] cell_1920_a_HPC2_and_a_reg;
  wire   [1:0] cell_1920_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1920_a_HPC2_and_mul;
  wire   [1:0] cell_1921_and_out;
  wire   [1:0] cell_1921_and_in;
  wire   [1:0] cell_1921_a_HPC2_and_a_reg;
  wire   [1:0] cell_1921_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1921_a_HPC2_and_mul;
  wire   [1:0] cell_1922_and_out;
  wire   [1:0] cell_1922_and_in;
  wire   [1:0] cell_1922_a_HPC2_and_a_reg;
  wire   [1:0] cell_1922_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1922_a_HPC2_and_mul;
  wire   [1:0] cell_1923_and_out;
  wire   [1:0] cell_1923_and_in;
  wire   [1:0] cell_1923_a_HPC2_and_a_reg;
  wire   [1:0] cell_1923_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1923_a_HPC2_and_mul;
  wire   [1:0] cell_1924_and_out;
  wire   [1:0] cell_1924_and_in;
  wire   [1:0] cell_1924_a_HPC2_and_a_reg;
  wire   [1:0] cell_1924_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1924_a_HPC2_and_mul;
  wire   [1:0] cell_1925_and_out;
  wire   [1:0] cell_1925_and_in;
  wire   [1:0] cell_1925_a_HPC2_and_a_reg;
  wire   [1:0] cell_1925_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1925_a_HPC2_and_mul;
  wire   [1:0] cell_1926_and_out;
  wire   [1:0] cell_1926_and_in;
  wire   [1:0] cell_1926_a_HPC2_and_a_reg;
  wire   [1:0] cell_1926_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1926_a_HPC2_and_mul;
  wire   [1:0] cell_1927_and_out;
  wire   [1:0] cell_1927_and_in;
  wire   [1:0] cell_1927_a_HPC2_and_a_reg;
  wire   [1:0] cell_1927_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1927_a_HPC2_and_mul;
  wire   [1:0] cell_1928_and_out;
  wire   [1:0] cell_1928_and_in;
  wire   [1:0] cell_1928_a_HPC2_and_a_reg;
  wire   [1:0] cell_1928_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1928_a_HPC2_and_mul;
  wire   [1:0] cell_1929_and_out;
  wire   [1:0] cell_1929_and_in;
  wire   [1:0] cell_1929_a_HPC2_and_a_reg;
  wire   [1:0] cell_1929_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1929_a_HPC2_and_mul;
  wire   [1:0] cell_1930_and_out;
  wire   [1:0] cell_1930_and_in;
  wire   [1:0] cell_1930_a_HPC2_and_a_reg;
  wire   [1:0] cell_1930_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1930_a_HPC2_and_mul;
  wire   [1:0] cell_1931_and_out;
  wire   [1:0] cell_1931_and_in;
  wire   [1:0] cell_1931_a_HPC2_and_a_reg;
  wire   [1:0] cell_1931_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1931_a_HPC2_and_mul;
  wire   [1:0] cell_1932_and_out;
  wire   [1:0] cell_1932_and_in;
  wire   [1:0] cell_1932_a_HPC2_and_a_reg;
  wire   [1:0] cell_1932_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1932_a_HPC2_and_mul;
  wire   [1:0] cell_1933_and_out;
  wire   [1:0] cell_1933_and_in;
  wire   [1:0] cell_1933_a_HPC2_and_a_reg;
  wire   [1:0] cell_1933_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1933_a_HPC2_and_mul;
  wire   [1:0] cell_1934_and_out;
  wire   [1:0] cell_1934_and_in;
  wire   [1:0] cell_1934_a_HPC2_and_a_reg;
  wire   [1:0] cell_1934_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1934_a_HPC2_and_mul;
  wire   [1:0] cell_1935_and_out;
  wire   [1:0] cell_1935_and_in;
  wire   [1:0] cell_1935_a_HPC2_and_a_reg;
  wire   [1:0] cell_1935_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1935_a_HPC2_and_mul;
  wire   [1:0] cell_1936_and_out;
  wire   [1:0] cell_1936_and_in;
  wire   [1:0] cell_1936_a_HPC2_and_a_reg;
  wire   [1:0] cell_1936_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1936_a_HPC2_and_mul;
  wire   [1:0] cell_1937_and_out;
  wire   [1:0] cell_1937_and_in;
  wire   [1:0] cell_1937_a_HPC2_and_a_reg;
  wire   [1:0] cell_1937_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1937_a_HPC2_and_mul;
  wire   [1:0] cell_1938_and_out;
  wire   [1:0] cell_1938_and_in;
  wire   [1:0] cell_1938_a_HPC2_and_a_reg;
  wire   [1:0] cell_1938_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1938_a_HPC2_and_mul;
  wire   [1:0] cell_1939_and_out;
  wire   [1:0] cell_1939_and_in;
  wire   [1:0] cell_1939_a_HPC2_and_a_reg;
  wire   [1:0] cell_1939_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1939_a_HPC2_and_mul;
  wire   [1:0] cell_1940_and_out;
  wire   [1:0] cell_1940_and_in;
  wire   [1:0] cell_1940_a_HPC2_and_a_reg;
  wire   [1:0] cell_1940_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1940_a_HPC2_and_mul;
  wire   [1:0] cell_1941_and_out;
  wire   [1:0] cell_1941_and_in;
  wire   [1:0] cell_1941_a_HPC2_and_a_reg;
  wire   [1:0] cell_1941_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1941_a_HPC2_and_mul;
  wire   [1:0] cell_1942_and_out;
  wire   [1:0] cell_1942_and_in;
  wire   [1:0] cell_1942_a_HPC2_and_a_reg;
  wire   [1:0] cell_1942_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1942_a_HPC2_and_mul;
  wire   [1:0] cell_1943_and_out;
  wire   [1:0] cell_1943_and_in;
  wire   [1:0] cell_1943_a_HPC2_and_a_reg;
  wire   [1:0] cell_1943_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1943_a_HPC2_and_mul;
  wire   [1:0] cell_1944_and_out;
  wire   [1:0] cell_1944_and_in;
  wire   [1:0] cell_1944_a_HPC2_and_a_reg;
  wire   [1:0] cell_1944_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1944_a_HPC2_and_mul;
  wire   [1:0] cell_1945_and_out;
  wire   [1:0] cell_1945_and_in;
  wire   [1:0] cell_1945_a_HPC2_and_a_reg;
  wire   [1:0] cell_1945_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1945_a_HPC2_and_mul;
  wire   [1:0] cell_1946_and_out;
  wire   [1:0] cell_1946_and_in;
  wire   [1:0] cell_1946_a_HPC2_and_a_reg;
  wire   [1:0] cell_1946_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1946_a_HPC2_and_mul;
  wire   [1:0] cell_1947_and_out;
  wire   [1:0] cell_1947_and_in;
  wire   [1:0] cell_1947_a_HPC2_and_a_reg;
  wire   [1:0] cell_1947_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1947_a_HPC2_and_mul;
  wire   [1:0] cell_1948_and_out;
  wire   [1:0] cell_1948_and_in;
  wire   [1:0] cell_1948_a_HPC2_and_a_reg;
  wire   [1:0] cell_1948_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1948_a_HPC2_and_mul;
  wire   [1:0] cell_1949_and_out;
  wire   [1:0] cell_1949_and_in;
  wire   [1:0] cell_1949_a_HPC2_and_a_reg;
  wire   [1:0] cell_1949_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1949_a_HPC2_and_mul;
  wire   [1:0] cell_1950_and_out;
  wire   [1:0] cell_1950_and_in;
  wire   [1:0] cell_1950_a_HPC2_and_a_reg;
  wire   [1:0] cell_1950_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1950_a_HPC2_and_mul;
  wire   [1:0] cell_1951_and_out;
  wire   [1:0] cell_1951_and_in;
  wire   [1:0] cell_1951_a_HPC2_and_a_reg;
  wire   [1:0] cell_1951_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1951_a_HPC2_and_mul;
  wire   [1:0] cell_1952_and_out;
  wire   [1:0] cell_1952_and_in;
  wire   [1:0] cell_1952_a_HPC2_and_a_reg;
  wire   [1:0] cell_1952_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1952_a_HPC2_and_mul;
  wire   [1:0] cell_1953_and_out;
  wire   [1:0] cell_1953_and_in;
  wire   [1:0] cell_1953_a_HPC2_and_a_reg;
  wire   [1:0] cell_1953_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1953_a_HPC2_and_mul;
  wire   [1:0] cell_1954_and_out;
  wire   [1:0] cell_1954_and_in;
  wire   [1:0] cell_1954_a_HPC2_and_a_reg;
  wire   [1:0] cell_1954_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1954_a_HPC2_and_mul;
  wire   [1:0] cell_1955_and_out;
  wire   [1:0] cell_1955_and_in;
  wire   [1:0] cell_1955_a_HPC2_and_a_reg;
  wire   [1:0] cell_1955_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1955_a_HPC2_and_mul;
  wire   [1:0] cell_1956_and_out;
  wire   [1:0] cell_1956_and_in;
  wire   [1:0] cell_1956_a_HPC2_and_a_reg;
  wire   [1:0] cell_1956_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1956_a_HPC2_and_mul;
  wire   [1:0] cell_1957_and_out;
  wire   [1:0] cell_1957_and_in;
  wire   [1:0] cell_1957_a_HPC2_and_a_reg;
  wire   [1:0] cell_1957_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1957_a_HPC2_and_mul;
  wire   [1:0] cell_1958_and_out;
  wire   [1:0] cell_1958_and_in;
  wire   [1:0] cell_1958_a_HPC2_and_a_reg;
  wire   [1:0] cell_1958_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1958_a_HPC2_and_mul;
  wire   [1:0] cell_1959_and_out;
  wire   [1:0] cell_1959_and_in;
  wire   [1:0] cell_1959_a_HPC2_and_a_reg;
  wire   [1:0] cell_1959_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1959_a_HPC2_and_mul;
  wire   [1:0] cell_1960_and_out;
  wire   [1:0] cell_1960_and_in;
  wire   [1:0] cell_1960_a_HPC2_and_a_reg;
  wire   [1:0] cell_1960_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1960_a_HPC2_and_mul;
  wire   [1:0] cell_1961_and_out;
  wire   [1:0] cell_1961_and_in;
  wire   [1:0] cell_1961_a_HPC2_and_a_reg;
  wire   [1:0] cell_1961_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1961_a_HPC2_and_mul;
  wire   [1:0] cell_1962_and_out;
  wire   [1:0] cell_1962_and_in;
  wire   [1:0] cell_1962_a_HPC2_and_a_reg;
  wire   [1:0] cell_1962_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1962_a_HPC2_and_mul;
  wire   [1:0] cell_1963_and_out;
  wire   [1:0] cell_1963_and_in;
  wire   [1:0] cell_1963_a_HPC2_and_a_reg;
  wire   [1:0] cell_1963_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1963_a_HPC2_and_mul;
  wire   [1:0] cell_1964_and_out;
  wire   [1:0] cell_1964_and_in;
  wire   [1:0] cell_1964_a_HPC2_and_a_reg;
  wire   [1:0] cell_1964_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1964_a_HPC2_and_mul;
  wire   [1:0] cell_1965_and_out;
  wire   [1:0] cell_1965_and_in;
  wire   [1:0] cell_1965_a_HPC2_and_a_reg;
  wire   [1:0] cell_1965_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1965_a_HPC2_and_mul;
  wire   [1:0] cell_1966_and_out;
  wire   [1:0] cell_1966_and_in;
  wire   [1:0] cell_1966_a_HPC2_and_a_reg;
  wire   [1:0] cell_1966_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1966_a_HPC2_and_mul;
  wire   [1:0] cell_1967_and_out;
  wire   [1:0] cell_1967_and_in;
  wire   [1:0] cell_1967_a_HPC2_and_a_reg;
  wire   [1:0] cell_1967_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1967_a_HPC2_and_mul;
  wire   [1:0] cell_1968_and_out;
  wire   [1:0] cell_1968_and_in;
  wire   [1:0] cell_1968_a_HPC2_and_a_reg;
  wire   [1:0] cell_1968_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1968_a_HPC2_and_mul;
  wire   [1:0] cell_1969_and_out;
  wire   [1:0] cell_1969_and_in;
  wire   [1:0] cell_1969_a_HPC2_and_a_reg;
  wire   [1:0] cell_1969_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1969_a_HPC2_and_mul;
  wire   [1:0] cell_1970_and_out;
  wire   [1:0] cell_1970_and_in;
  wire   [1:0] cell_1970_a_HPC2_and_a_reg;
  wire   [1:0] cell_1970_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1970_a_HPC2_and_mul;
  wire   [1:0] cell_1971_and_out;
  wire   [1:0] cell_1971_and_in;
  wire   [1:0] cell_1971_a_HPC2_and_a_reg;
  wire   [1:0] cell_1971_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1971_a_HPC2_and_mul;
  wire   [1:0] cell_1972_and_out;
  wire   [1:0] cell_1972_and_in;
  wire   [1:0] cell_1972_a_HPC2_and_a_reg;
  wire   [1:0] cell_1972_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1972_a_HPC2_and_mul;
  wire   [1:0] cell_1973_and_out;
  wire   [1:0] cell_1973_and_in;
  wire   [1:0] cell_1973_a_HPC2_and_a_reg;
  wire   [1:0] cell_1973_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1973_a_HPC2_and_mul;
  wire   [1:0] cell_1974_and_out;
  wire   [1:0] cell_1974_and_in;
  wire   [1:0] cell_1974_a_HPC2_and_a_reg;
  wire   [1:0] cell_1974_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1974_a_HPC2_and_mul;
  wire   [1:0] cell_1975_and_out;
  wire   [1:0] cell_1975_and_in;
  wire   [1:0] cell_1975_a_HPC2_and_a_reg;
  wire   [1:0] cell_1975_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1975_a_HPC2_and_mul;
  wire   [1:0] cell_1976_and_out;
  wire   [1:0] cell_1976_and_in;
  wire   [1:0] cell_1976_a_HPC2_and_a_reg;
  wire   [1:0] cell_1976_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1976_a_HPC2_and_mul;
  wire   [1:0] cell_1977_and_out;
  wire   [1:0] cell_1977_and_in;
  wire   [1:0] cell_1977_a_HPC2_and_a_reg;
  wire   [1:0] cell_1977_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1977_a_HPC2_and_mul;
  wire   [1:0] cell_1978_and_out;
  wire   [1:0] cell_1978_and_in;
  wire   [1:0] cell_1978_a_HPC2_and_a_reg;
  wire   [1:0] cell_1978_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1978_a_HPC2_and_mul;
  wire   [1:0] cell_1979_and_out;
  wire   [1:0] cell_1979_and_in;
  wire   [1:0] cell_1979_a_HPC2_and_a_reg;
  wire   [1:0] cell_1979_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1979_a_HPC2_and_mul;
  wire   [1:0] cell_1980_and_out;
  wire   [1:0] cell_1980_and_in;
  wire   [1:0] cell_1980_a_HPC2_and_a_reg;
  wire   [1:0] cell_1980_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1980_a_HPC2_and_mul;
  wire   [1:0] cell_1981_and_out;
  wire   [1:0] cell_1981_and_in;
  wire   [1:0] cell_1981_a_HPC2_and_a_reg;
  wire   [1:0] cell_1981_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1981_a_HPC2_and_mul;
  wire   [1:0] cell_1982_and_out;
  wire   [1:0] cell_1982_and_in;
  wire   [1:0] cell_1982_a_HPC2_and_a_reg;
  wire   [1:0] cell_1982_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1982_a_HPC2_and_mul;
  wire   [1:0] cell_1983_and_out;
  wire   [1:0] cell_1983_and_in;
  wire   [1:0] cell_1983_a_HPC2_and_a_reg;
  wire   [1:0] cell_1983_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1983_a_HPC2_and_mul;
  wire   [1:0] cell_1984_and_out;
  wire   [1:0] cell_1984_and_in;
  wire   [1:0] cell_1984_a_HPC2_and_a_reg;
  wire   [1:0] cell_1984_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1984_a_HPC2_and_mul;
  wire   [1:0] cell_1985_and_out;
  wire   [1:0] cell_1985_and_in;
  wire   [1:0] cell_1985_a_HPC2_and_a_reg;
  wire   [1:0] cell_1985_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1985_a_HPC2_and_mul;
  wire   [1:0] cell_1986_and_out;
  wire   [1:0] cell_1986_and_in;
  wire   [1:0] cell_1986_a_HPC2_and_a_reg;
  wire   [1:0] cell_1986_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1986_a_HPC2_and_mul;
  wire   [1:0] cell_1987_and_out;
  wire   [1:0] cell_1987_and_in;
  wire   [1:0] cell_1987_a_HPC2_and_a_reg;
  wire   [1:0] cell_1987_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1987_a_HPC2_and_mul;
  wire   [1:0] cell_1988_and_out;
  wire   [1:0] cell_1988_and_in;
  wire   [1:0] cell_1988_a_HPC2_and_a_reg;
  wire   [1:0] cell_1988_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1988_a_HPC2_and_mul;
  wire   [1:0] cell_1989_and_out;
  wire   [1:0] cell_1989_and_in;
  wire   [1:0] cell_1989_a_HPC2_and_a_reg;
  wire   [1:0] cell_1989_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1989_a_HPC2_and_mul;
  wire   [1:0] cell_1990_and_out;
  wire   [1:0] cell_1990_and_in;
  wire   [1:0] cell_1990_a_HPC2_and_a_reg;
  wire   [1:0] cell_1990_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1990_a_HPC2_and_mul;
  wire   [1:0] cell_1991_and_out;
  wire   [1:0] cell_1991_and_in;
  wire   [1:0] cell_1991_a_HPC2_and_a_reg;
  wire   [1:0] cell_1991_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1991_a_HPC2_and_mul;
  wire   [1:0] cell_1992_and_out;
  wire   [1:0] cell_1992_and_in;
  wire   [1:0] cell_1992_a_HPC2_and_a_reg;
  wire   [1:0] cell_1992_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1992_a_HPC2_and_mul;
  wire   [1:0] cell_1993_and_out;
  wire   [1:0] cell_1993_and_in;
  wire   [1:0] cell_1993_a_HPC2_and_a_reg;
  wire   [1:0] cell_1993_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1993_a_HPC2_and_mul;
  wire   [1:0] cell_1994_and_out;
  wire   [1:0] cell_1994_and_in;
  wire   [1:0] cell_1994_a_HPC2_and_a_reg;
  wire   [1:0] cell_1994_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1994_a_HPC2_and_mul;
  wire   [1:0] cell_1995_and_out;
  wire   [1:0] cell_1995_and_in;
  wire   [1:0] cell_1995_a_HPC2_and_a_reg;
  wire   [1:0] cell_1995_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1995_a_HPC2_and_mul;
  wire   [1:0] cell_1996_and_out;
  wire   [1:0] cell_1996_and_in;
  wire   [1:0] cell_1996_a_HPC2_and_a_reg;
  wire   [1:0] cell_1996_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1996_a_HPC2_and_mul;
  wire   [1:0] cell_1997_and_out;
  wire   [1:0] cell_1997_and_in;
  wire   [1:0] cell_1997_a_HPC2_and_a_reg;
  wire   [1:0] cell_1997_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1997_a_HPC2_and_mul;
  wire   [1:0] cell_1998_and_out;
  wire   [1:0] cell_1998_and_in;
  wire   [1:0] cell_1998_a_HPC2_and_a_reg;
  wire   [1:0] cell_1998_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1998_a_HPC2_and_mul;
  wire   [1:0] cell_1999_and_out;
  wire   [1:0] cell_1999_and_in;
  wire   [1:0] cell_1999_a_HPC2_and_a_reg;
  wire   [1:0] cell_1999_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_1999_a_HPC2_and_mul;
  wire   [1:0] cell_2000_and_out;
  wire   [1:0] cell_2000_and_in;
  wire   [1:0] cell_2000_a_HPC2_and_a_reg;
  wire   [1:0] cell_2000_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2000_a_HPC2_and_mul;
  wire   [1:0] cell_2001_and_out;
  wire   [1:0] cell_2001_and_in;
  wire   [1:0] cell_2001_a_HPC2_and_a_reg;
  wire   [1:0] cell_2001_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2001_a_HPC2_and_mul;
  wire   [1:0] cell_2002_and_out;
  wire   [1:0] cell_2002_and_in;
  wire   [1:0] cell_2002_a_HPC2_and_a_reg;
  wire   [1:0] cell_2002_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2002_a_HPC2_and_mul;
  wire   [1:0] cell_2003_and_out;
  wire   [1:0] cell_2003_and_in;
  wire   [1:0] cell_2003_a_HPC2_and_a_reg;
  wire   [1:0] cell_2003_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2003_a_HPC2_and_mul;
  wire   [1:0] cell_2004_and_out;
  wire   [1:0] cell_2004_and_in;
  wire   [1:0] cell_2004_a_HPC2_and_a_reg;
  wire   [1:0] cell_2004_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2004_a_HPC2_and_mul;
  wire   [1:0] cell_2005_and_out;
  wire   [1:0] cell_2005_and_in;
  wire   [1:0] cell_2005_a_HPC2_and_a_reg;
  wire   [1:0] cell_2005_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2005_a_HPC2_and_mul;
  wire   [1:0] cell_2006_and_out;
  wire   [1:0] cell_2006_and_in;
  wire   [1:0] cell_2006_a_HPC2_and_a_reg;
  wire   [1:0] cell_2006_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2006_a_HPC2_and_mul;
  wire   [1:0] cell_2007_and_out;
  wire   [1:0] cell_2007_and_in;
  wire   [1:0] cell_2007_a_HPC2_and_a_reg;
  wire   [1:0] cell_2007_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2007_a_HPC2_and_mul;
  wire   [1:0] cell_2008_and_out;
  wire   [1:0] cell_2008_and_in;
  wire   [1:0] cell_2008_a_HPC2_and_a_reg;
  wire   [1:0] cell_2008_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2008_a_HPC2_and_mul;
  wire   [1:0] cell_2009_and_out;
  wire   [1:0] cell_2009_and_in;
  wire   [1:0] cell_2009_a_HPC2_and_a_reg;
  wire   [1:0] cell_2009_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2009_a_HPC2_and_mul;
  wire   [1:0] cell_2010_and_out;
  wire   [1:0] cell_2010_and_in;
  wire   [1:0] cell_2010_a_HPC2_and_a_reg;
  wire   [1:0] cell_2010_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2010_a_HPC2_and_mul;
  wire   [1:0] cell_2011_and_out;
  wire   [1:0] cell_2011_and_in;
  wire   [1:0] cell_2011_a_HPC2_and_a_reg;
  wire   [1:0] cell_2011_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2011_a_HPC2_and_mul;
  wire   [1:0] cell_2012_and_out;
  wire   [1:0] cell_2012_and_in;
  wire   [1:0] cell_2012_a_HPC2_and_a_reg;
  wire   [1:0] cell_2012_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2012_a_HPC2_and_mul;
  wire   [1:0] cell_2013_and_out;
  wire   [1:0] cell_2013_and_in;
  wire   [1:0] cell_2013_a_HPC2_and_a_reg;
  wire   [1:0] cell_2013_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2013_a_HPC2_and_mul;
  wire   [1:0] cell_2014_and_out;
  wire   [1:0] cell_2014_and_in;
  wire   [1:0] cell_2014_a_HPC2_and_a_reg;
  wire   [1:0] cell_2014_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2014_a_HPC2_and_mul;
  wire   [1:0] cell_2015_and_out;
  wire   [1:0] cell_2015_and_in;
  wire   [1:0] cell_2015_a_HPC2_and_a_reg;
  wire   [1:0] cell_2015_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2015_a_HPC2_and_mul;
  wire   [1:0] cell_2016_and_out;
  wire   [1:0] cell_2016_and_in;
  wire   [1:0] cell_2016_a_HPC2_and_a_reg;
  wire   [1:0] cell_2016_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2016_a_HPC2_and_mul;
  wire   [1:0] cell_2017_and_out;
  wire   [1:0] cell_2017_and_in;
  wire   [1:0] cell_2017_a_HPC2_and_a_reg;
  wire   [1:0] cell_2017_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2017_a_HPC2_and_mul;
  wire   [1:0] cell_2018_and_out;
  wire   [1:0] cell_2018_and_in;
  wire   [1:0] cell_2018_a_HPC2_and_a_reg;
  wire   [1:0] cell_2018_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2018_a_HPC2_and_mul;
  wire   [1:0] cell_2019_and_out;
  wire   [1:0] cell_2019_and_in;
  wire   [1:0] cell_2019_a_HPC2_and_a_reg;
  wire   [1:0] cell_2019_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2019_a_HPC2_and_mul;
  wire   [1:0] cell_2020_and_out;
  wire   [1:0] cell_2020_and_in;
  wire   [1:0] cell_2020_a_HPC2_and_a_reg;
  wire   [1:0] cell_2020_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2020_a_HPC2_and_mul;
  wire   [1:0] cell_2021_and_out;
  wire   [1:0] cell_2021_and_in;
  wire   [1:0] cell_2021_a_HPC2_and_a_reg;
  wire   [1:0] cell_2021_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2021_a_HPC2_and_mul;
  wire   [1:0] cell_2022_and_out;
  wire   [1:0] cell_2022_and_in;
  wire   [1:0] cell_2022_a_HPC2_and_a_reg;
  wire   [1:0] cell_2022_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2022_a_HPC2_and_mul;
  wire   [1:0] cell_2023_and_out;
  wire   [1:0] cell_2023_and_in;
  wire   [1:0] cell_2023_a_HPC2_and_a_reg;
  wire   [1:0] cell_2023_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2023_a_HPC2_and_mul;
  wire   [1:0] cell_2024_and_out;
  wire   [1:0] cell_2024_and_in;
  wire   [1:0] cell_2024_a_HPC2_and_a_reg;
  wire   [1:0] cell_2024_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2024_a_HPC2_and_mul;
  wire   [1:0] cell_2025_and_out;
  wire   [1:0] cell_2025_and_in;
  wire   [1:0] cell_2025_a_HPC2_and_a_reg;
  wire   [1:0] cell_2025_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2025_a_HPC2_and_mul;
  wire   [1:0] cell_2026_and_out;
  wire   [1:0] cell_2026_and_in;
  wire   [1:0] cell_2026_a_HPC2_and_a_reg;
  wire   [1:0] cell_2026_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2026_a_HPC2_and_mul;
  wire   [1:0] cell_2027_and_out;
  wire   [1:0] cell_2027_and_in;
  wire   [1:0] cell_2027_a_HPC2_and_a_reg;
  wire   [1:0] cell_2027_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2027_a_HPC2_and_mul;
  wire   [1:0] cell_2028_and_out;
  wire   [1:0] cell_2028_and_in;
  wire   [1:0] cell_2028_a_HPC2_and_a_reg;
  wire   [1:0] cell_2028_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2028_a_HPC2_and_mul;
  wire   [1:0] cell_2029_and_out;
  wire   [1:0] cell_2029_and_in;
  wire   [1:0] cell_2029_a_HPC2_and_a_reg;
  wire   [1:0] cell_2029_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2029_a_HPC2_and_mul;
  wire   [1:0] cell_2030_and_out;
  wire   [1:0] cell_2030_and_in;
  wire   [1:0] cell_2030_a_HPC2_and_a_reg;
  wire   [1:0] cell_2030_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2030_a_HPC2_and_mul;
  wire   [1:0] cell_2031_and_out;
  wire   [1:0] cell_2031_and_in;
  wire   [1:0] cell_2031_a_HPC2_and_a_reg;
  wire   [1:0] cell_2031_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2031_a_HPC2_and_mul;
  wire   [1:0] cell_2032_and_out;
  wire   [1:0] cell_2032_and_in;
  wire   [1:0] cell_2032_a_HPC2_and_a_reg;
  wire   [1:0] cell_2032_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2032_a_HPC2_and_mul;
  wire   [1:0] cell_2033_and_out;
  wire   [1:0] cell_2033_and_in;
  wire   [1:0] cell_2033_a_HPC2_and_a_reg;
  wire   [1:0] cell_2033_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2033_a_HPC2_and_mul;
  wire   [1:0] cell_2034_and_out;
  wire   [1:0] cell_2034_and_in;
  wire   [1:0] cell_2034_a_HPC2_and_a_reg;
  wire   [1:0] cell_2034_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2034_a_HPC2_and_mul;
  wire   [1:0] cell_2035_and_out;
  wire   [1:0] cell_2035_and_in;
  wire   [1:0] cell_2035_a_HPC2_and_a_reg;
  wire   [1:0] cell_2035_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2035_a_HPC2_and_mul;
  wire   [1:0] cell_2036_and_out;
  wire   [1:0] cell_2036_and_in;
  wire   [1:0] cell_2036_a_HPC2_and_a_reg;
  wire   [1:0] cell_2036_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2036_a_HPC2_and_mul;
  wire   [1:0] cell_2037_and_out;
  wire   [1:0] cell_2037_and_in;
  wire   [1:0] cell_2037_a_HPC2_and_a_reg;
  wire   [1:0] cell_2037_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2037_a_HPC2_and_mul;
  wire   [1:0] cell_2038_and_out;
  wire   [1:0] cell_2038_and_in;
  wire   [1:0] cell_2038_a_HPC2_and_a_reg;
  wire   [1:0] cell_2038_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2038_a_HPC2_and_mul;
  wire   [1:0] cell_2039_and_out;
  wire   [1:0] cell_2039_and_in;
  wire   [1:0] cell_2039_a_HPC2_and_a_reg;
  wire   [1:0] cell_2039_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2039_a_HPC2_and_mul;
  wire   [1:0] cell_2040_and_out;
  wire   [1:0] cell_2040_and_in;
  wire   [1:0] cell_2040_a_HPC2_and_a_reg;
  wire   [1:0] cell_2040_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2040_a_HPC2_and_mul;
  wire   [1:0] cell_2041_and_out;
  wire   [1:0] cell_2041_and_in;
  wire   [1:0] cell_2041_a_HPC2_and_a_reg;
  wire   [1:0] cell_2041_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2041_a_HPC2_and_mul;
  wire   [1:0] cell_2042_and_out;
  wire   [1:0] cell_2042_and_in;
  wire   [1:0] cell_2042_a_HPC2_and_a_reg;
  wire   [1:0] cell_2042_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2042_a_HPC2_and_mul;
  wire   [1:0] cell_2043_and_out;
  wire   [1:0] cell_2043_and_in;
  wire   [1:0] cell_2043_a_HPC2_and_a_reg;
  wire   [1:0] cell_2043_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2043_a_HPC2_and_mul;
  wire   [1:0] cell_2044_and_out;
  wire   [1:0] cell_2044_and_in;
  wire   [1:0] cell_2044_a_HPC2_and_a_reg;
  wire   [1:0] cell_2044_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2044_a_HPC2_and_mul;
  wire   [1:0] cell_2045_and_out;
  wire   [1:0] cell_2045_and_in;
  wire   [1:0] cell_2045_a_HPC2_and_a_reg;
  wire   [1:0] cell_2045_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2045_a_HPC2_and_mul;
  wire   [1:0] cell_2046_and_out;
  wire   [1:0] cell_2046_and_in;
  wire   [1:0] cell_2046_a_HPC2_and_a_reg;
  wire   [1:0] cell_2046_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2046_a_HPC2_and_mul;
  wire   [1:0] cell_2047_and_out;
  wire   [1:0] cell_2047_and_in;
  wire   [1:0] cell_2047_a_HPC2_and_a_reg;
  wire   [1:0] cell_2047_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2047_a_HPC2_and_mul;
  wire   [1:0] cell_2048_and_out;
  wire   [1:0] cell_2048_and_in;
  wire   [1:0] cell_2048_a_HPC2_and_a_reg;
  wire   [1:0] cell_2048_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2048_a_HPC2_and_mul;
  wire   [1:0] cell_2049_and_out;
  wire   [1:0] cell_2049_and_in;
  wire   [1:0] cell_2049_a_HPC2_and_a_reg;
  wire   [1:0] cell_2049_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2049_a_HPC2_and_mul;
  wire   [1:0] cell_2050_and_out;
  wire   [1:0] cell_2050_and_in;
  wire   [1:0] cell_2050_a_HPC2_and_a_reg;
  wire   [1:0] cell_2050_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2050_a_HPC2_and_mul;
  wire   [1:0] cell_2051_and_out;
  wire   [1:0] cell_2051_and_in;
  wire   [1:0] cell_2051_a_HPC2_and_a_reg;
  wire   [1:0] cell_2051_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2051_a_HPC2_and_mul;
  wire   [1:0] cell_2052_and_out;
  wire   [1:0] cell_2052_and_in;
  wire   [1:0] cell_2052_a_HPC2_and_a_reg;
  wire   [1:0] cell_2052_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2052_a_HPC2_and_mul;
  wire   [1:0] cell_2053_and_out;
  wire   [1:0] cell_2053_and_in;
  wire   [1:0] cell_2053_a_HPC2_and_a_reg;
  wire   [1:0] cell_2053_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2053_a_HPC2_and_mul;
  wire   [1:0] cell_2054_and_out;
  wire   [1:0] cell_2054_and_in;
  wire   [1:0] cell_2054_a_HPC2_and_a_reg;
  wire   [1:0] cell_2054_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2054_a_HPC2_and_mul;
  wire   [1:0] cell_2055_and_out;
  wire   [1:0] cell_2055_and_in;
  wire   [1:0] cell_2055_a_HPC2_and_a_reg;
  wire   [1:0] cell_2055_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2055_a_HPC2_and_mul;
  wire   [1:0] cell_2056_and_out;
  wire   [1:0] cell_2056_and_in;
  wire   [1:0] cell_2056_a_HPC2_and_a_reg;
  wire   [1:0] cell_2056_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2056_a_HPC2_and_mul;
  wire   [1:0] cell_2057_and_out;
  wire   [1:0] cell_2057_and_in;
  wire   [1:0] cell_2057_a_HPC2_and_a_reg;
  wire   [1:0] cell_2057_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2057_a_HPC2_and_mul;
  wire   [1:0] cell_2058_and_out;
  wire   [1:0] cell_2058_and_in;
  wire   [1:0] cell_2058_a_HPC2_and_a_reg;
  wire   [1:0] cell_2058_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2058_a_HPC2_and_mul;
  wire   [1:0] cell_2059_and_out;
  wire   [1:0] cell_2059_and_in;
  wire   [1:0] cell_2059_a_HPC2_and_a_reg;
  wire   [1:0] cell_2059_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2059_a_HPC2_and_mul;
  wire   [1:0] cell_2060_and_out;
  wire   [1:0] cell_2060_and_in;
  wire   [1:0] cell_2060_a_HPC2_and_a_reg;
  wire   [1:0] cell_2060_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2060_a_HPC2_and_mul;
  wire   [1:0] cell_2061_and_out;
  wire   [1:0] cell_2061_and_in;
  wire   [1:0] cell_2061_a_HPC2_and_a_reg;
  wire   [1:0] cell_2061_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2061_a_HPC2_and_mul;
  wire   [1:0] cell_2062_and_out;
  wire   [1:0] cell_2062_and_in;
  wire   [1:0] cell_2062_a_HPC2_and_a_reg;
  wire   [1:0] cell_2062_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2062_a_HPC2_and_mul;
  wire   [1:0] cell_2063_and_out;
  wire   [1:0] cell_2063_and_in;
  wire   [1:0] cell_2063_a_HPC2_and_a_reg;
  wire   [1:0] cell_2063_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2063_a_HPC2_and_mul;
  wire   [1:0] cell_2064_and_out;
  wire   [1:0] cell_2064_and_in;
  wire   [1:0] cell_2064_a_HPC2_and_a_reg;
  wire   [1:0] cell_2064_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2064_a_HPC2_and_mul;
  wire   [1:0] cell_2065_and_out;
  wire   [1:0] cell_2065_and_in;
  wire   [1:0] cell_2065_a_HPC2_and_a_reg;
  wire   [1:0] cell_2065_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2065_a_HPC2_and_mul;
  wire   [1:0] cell_2066_and_out;
  wire   [1:0] cell_2066_and_in;
  wire   [1:0] cell_2066_a_HPC2_and_a_reg;
  wire   [1:0] cell_2066_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2066_a_HPC2_and_mul;
  wire   [1:0] cell_2067_and_out;
  wire   [1:0] cell_2067_and_in;
  wire   [1:0] cell_2067_a_HPC2_and_a_reg;
  wire   [1:0] cell_2067_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2067_a_HPC2_and_mul;
  wire   [1:0] cell_2068_and_out;
  wire   [1:0] cell_2068_and_in;
  wire   [1:0] cell_2068_a_HPC2_and_a_reg;
  wire   [1:0] cell_2068_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2068_a_HPC2_and_mul;
  wire   [1:0] cell_2069_and_out;
  wire   [1:0] cell_2069_and_in;
  wire   [1:0] cell_2069_a_HPC2_and_a_reg;
  wire   [1:0] cell_2069_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2069_a_HPC2_and_mul;
  wire   [1:0] cell_2070_and_out;
  wire   [1:0] cell_2070_and_in;
  wire   [1:0] cell_2070_a_HPC2_and_a_reg;
  wire   [1:0] cell_2070_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2070_a_HPC2_and_mul;
  wire   [1:0] cell_2071_and_out;
  wire   [1:0] cell_2071_and_in;
  wire   [1:0] cell_2071_a_HPC2_and_a_reg;
  wire   [1:0] cell_2071_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2071_a_HPC2_and_mul;
  wire   [1:0] cell_2072_and_out;
  wire   [1:0] cell_2072_and_in;
  wire   [1:0] cell_2072_a_HPC2_and_a_reg;
  wire   [1:0] cell_2072_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2072_a_HPC2_and_mul;
  wire   [1:0] cell_2073_and_out;
  wire   [1:0] cell_2073_and_in;
  wire   [1:0] cell_2073_a_HPC2_and_a_reg;
  wire   [1:0] cell_2073_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2073_a_HPC2_and_mul;
  wire   [1:0] cell_2074_and_out;
  wire   [1:0] cell_2074_and_in;
  wire   [1:0] cell_2074_a_HPC2_and_a_reg;
  wire   [1:0] cell_2074_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2074_a_HPC2_and_mul;
  wire   [1:0] cell_2075_and_out;
  wire   [1:0] cell_2075_and_in;
  wire   [1:0] cell_2075_a_HPC2_and_a_reg;
  wire   [1:0] cell_2075_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2075_a_HPC2_and_mul;
  wire   [1:0] cell_2076_and_out;
  wire   [1:0] cell_2076_and_in;
  wire   [1:0] cell_2076_a_HPC2_and_a_reg;
  wire   [1:0] cell_2076_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2076_a_HPC2_and_mul;
  wire   [1:0] cell_2077_and_out;
  wire   [1:0] cell_2077_and_in;
  wire   [1:0] cell_2077_a_HPC2_and_a_reg;
  wire   [1:0] cell_2077_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2077_a_HPC2_and_mul;
  wire   [1:0] cell_2078_and_out;
  wire   [1:0] cell_2078_and_in;
  wire   [1:0] cell_2078_a_HPC2_and_a_reg;
  wire   [1:0] cell_2078_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2078_a_HPC2_and_mul;
  wire   [1:0] cell_2079_and_out;
  wire   [1:0] cell_2079_and_in;
  wire   [1:0] cell_2079_a_HPC2_and_a_reg;
  wire   [1:0] cell_2079_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2079_a_HPC2_and_mul;
  wire   [1:0] cell_2080_and_out;
  wire   [1:0] cell_2080_and_in;
  wire   [1:0] cell_2080_a_HPC2_and_a_reg;
  wire   [1:0] cell_2080_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2080_a_HPC2_and_mul;
  wire   [1:0] cell_2081_and_out;
  wire   [1:0] cell_2081_and_in;
  wire   [1:0] cell_2081_a_HPC2_and_a_reg;
  wire   [1:0] cell_2081_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2081_a_HPC2_and_mul;
  wire   [1:0] cell_2082_and_out;
  wire   [1:0] cell_2082_and_in;
  wire   [1:0] cell_2082_a_HPC2_and_a_reg;
  wire   [1:0] cell_2082_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2082_a_HPC2_and_mul;
  wire   [1:0] cell_2083_and_out;
  wire   [1:0] cell_2083_and_in;
  wire   [1:0] cell_2083_a_HPC2_and_a_reg;
  wire   [1:0] cell_2083_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2083_a_HPC2_and_mul;
  wire   [1:0] cell_2084_and_out;
  wire   [1:0] cell_2084_and_in;
  wire   [1:0] cell_2084_a_HPC2_and_a_reg;
  wire   [1:0] cell_2084_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2084_a_HPC2_and_mul;
  wire   [1:0] cell_2085_and_out;
  wire   [1:0] cell_2085_and_in;
  wire   [1:0] cell_2085_a_HPC2_and_a_reg;
  wire   [1:0] cell_2085_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2085_a_HPC2_and_mul;
  wire   [1:0] cell_2086_and_out;
  wire   [1:0] cell_2086_and_in;
  wire   [1:0] cell_2086_a_HPC2_and_a_reg;
  wire   [1:0] cell_2086_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2086_a_HPC2_and_mul;
  wire   [1:0] cell_2087_and_out;
  wire   [1:0] cell_2087_and_in;
  wire   [1:0] cell_2087_a_HPC2_and_a_reg;
  wire   [1:0] cell_2087_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2087_a_HPC2_and_mul;
  wire   [1:0] cell_2088_and_out;
  wire   [1:0] cell_2088_and_in;
  wire   [1:0] cell_2088_a_HPC2_and_a_reg;
  wire   [1:0] cell_2088_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2088_a_HPC2_and_mul;
  wire   [1:0] cell_2089_and_out;
  wire   [1:0] cell_2089_and_in;
  wire   [1:0] cell_2089_a_HPC2_and_a_reg;
  wire   [1:0] cell_2089_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2089_a_HPC2_and_mul;
  wire   [1:0] cell_2090_and_out;
  wire   [1:0] cell_2090_and_in;
  wire   [1:0] cell_2090_a_HPC2_and_a_reg;
  wire   [1:0] cell_2090_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2090_a_HPC2_and_mul;
  wire   [1:0] cell_2091_and_out;
  wire   [1:0] cell_2091_and_in;
  wire   [1:0] cell_2091_a_HPC2_and_a_reg;
  wire   [1:0] cell_2091_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2091_a_HPC2_and_mul;
  wire   [1:0] cell_2092_and_out;
  wire   [1:0] cell_2092_and_in;
  wire   [1:0] cell_2092_a_HPC2_and_a_reg;
  wire   [1:0] cell_2092_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2092_a_HPC2_and_mul;
  wire   [1:0] cell_2093_and_out;
  wire   [1:0] cell_2093_and_in;
  wire   [1:0] cell_2093_a_HPC2_and_a_reg;
  wire   [1:0] cell_2093_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2093_a_HPC2_and_mul;
  wire   [1:0] cell_2094_and_out;
  wire   [1:0] cell_2094_and_in;
  wire   [1:0] cell_2094_a_HPC2_and_a_reg;
  wire   [1:0] cell_2094_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2094_a_HPC2_and_mul;
  wire   [1:0] cell_2095_and_out;
  wire   [1:0] cell_2095_and_in;
  wire   [1:0] cell_2095_a_HPC2_and_a_reg;
  wire   [1:0] cell_2095_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2095_a_HPC2_and_mul;
  wire   [1:0] cell_2096_and_out;
  wire   [1:0] cell_2096_and_in;
  wire   [1:0] cell_2096_a_HPC2_and_a_reg;
  wire   [1:0] cell_2096_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2096_a_HPC2_and_mul;
  wire   [1:0] cell_2097_and_out;
  wire   [1:0] cell_2097_and_in;
  wire   [1:0] cell_2097_a_HPC2_and_a_reg;
  wire   [1:0] cell_2097_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2097_a_HPC2_and_mul;
  wire   [1:0] cell_2098_and_out;
  wire   [1:0] cell_2098_and_in;
  wire   [1:0] cell_2098_a_HPC2_and_a_reg;
  wire   [1:0] cell_2098_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2098_a_HPC2_and_mul;
  wire   [1:0] cell_2099_and_out;
  wire   [1:0] cell_2099_and_in;
  wire   [1:0] cell_2099_a_HPC2_and_a_reg;
  wire   [1:0] cell_2099_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2099_a_HPC2_and_mul;
  wire   [1:0] cell_2100_and_out;
  wire   [1:0] cell_2100_and_in;
  wire   [1:0] cell_2100_a_HPC2_and_a_reg;
  wire   [1:0] cell_2100_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2100_a_HPC2_and_mul;
  wire   [1:0] cell_2101_and_out;
  wire   [1:0] cell_2101_and_in;
  wire   [1:0] cell_2101_a_HPC2_and_a_reg;
  wire   [1:0] cell_2101_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2101_a_HPC2_and_mul;
  wire   [1:0] cell_2102_and_out;
  wire   [1:0] cell_2102_and_in;
  wire   [1:0] cell_2102_a_HPC2_and_a_reg;
  wire   [1:0] cell_2102_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2102_a_HPC2_and_mul;
  wire   [1:0] cell_2103_and_out;
  wire   [1:0] cell_2103_and_in;
  wire   [1:0] cell_2103_a_HPC2_and_a_reg;
  wire   [1:0] cell_2103_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2103_a_HPC2_and_mul;
  wire   [1:0] cell_2104_and_out;
  wire   [1:0] cell_2104_and_in;
  wire   [1:0] cell_2104_a_HPC2_and_a_reg;
  wire   [1:0] cell_2104_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2104_a_HPC2_and_mul;
  wire   [1:0] cell_2105_and_out;
  wire   [1:0] cell_2105_and_in;
  wire   [1:0] cell_2105_a_HPC2_and_a_reg;
  wire   [1:0] cell_2105_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2105_a_HPC2_and_mul;
  wire   [1:0] cell_2106_and_out;
  wire   [1:0] cell_2106_and_in;
  wire   [1:0] cell_2106_a_HPC2_and_a_reg;
  wire   [1:0] cell_2106_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2106_a_HPC2_and_mul;
  wire   [1:0] cell_2107_and_out;
  wire   [1:0] cell_2107_and_in;
  wire   [1:0] cell_2107_a_HPC2_and_a_reg;
  wire   [1:0] cell_2107_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2107_a_HPC2_and_mul;
  wire   [1:0] cell_2108_and_out;
  wire   [1:0] cell_2108_and_in;
  wire   [1:0] cell_2108_a_HPC2_and_a_reg;
  wire   [1:0] cell_2108_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2108_a_HPC2_and_mul;
  wire   [1:0] cell_2109_and_out;
  wire   [1:0] cell_2109_and_in;
  wire   [1:0] cell_2109_a_HPC2_and_a_reg;
  wire   [1:0] cell_2109_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2109_a_HPC2_and_mul;
  wire   [1:0] cell_2110_and_out;
  wire   [1:0] cell_2110_and_in;
  wire   [1:0] cell_2110_a_HPC2_and_a_reg;
  wire   [1:0] cell_2110_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2110_a_HPC2_and_mul;
  wire   [1:0] cell_2111_and_out;
  wire   [1:0] cell_2111_and_in;
  wire   [1:0] cell_2111_a_HPC2_and_a_reg;
  wire   [1:0] cell_2111_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2111_a_HPC2_and_mul;
  wire   [1:0] cell_2112_and_out;
  wire   [1:0] cell_2112_and_in;
  wire   [1:0] cell_2112_a_HPC2_and_a_reg;
  wire   [1:0] cell_2112_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2112_a_HPC2_and_mul;
  wire   [1:0] cell_2113_and_out;
  wire   [1:0] cell_2113_and_in;
  wire   [1:0] cell_2113_a_HPC2_and_a_reg;
  wire   [1:0] cell_2113_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2113_a_HPC2_and_mul;
  wire   [1:0] cell_2114_and_out;
  wire   [1:0] cell_2114_and_in;
  wire   [1:0] cell_2114_a_HPC2_and_a_reg;
  wire   [1:0] cell_2114_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2114_a_HPC2_and_mul;
  wire   [1:0] cell_2115_and_out;
  wire   [1:0] cell_2115_and_in;
  wire   [1:0] cell_2115_a_HPC2_and_a_reg;
  wire   [1:0] cell_2115_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2115_a_HPC2_and_mul;
  wire   [1:0] cell_2116_and_out;
  wire   [1:0] cell_2116_and_in;
  wire   [1:0] cell_2116_a_HPC2_and_a_reg;
  wire   [1:0] cell_2116_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2116_a_HPC2_and_mul;
  wire   [1:0] cell_2117_and_out;
  wire   [1:0] cell_2117_and_in;
  wire   [1:0] cell_2117_a_HPC2_and_a_reg;
  wire   [1:0] cell_2117_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2117_a_HPC2_and_mul;
  wire   [1:0] cell_2118_and_out;
  wire   [1:0] cell_2118_and_in;
  wire   [1:0] cell_2118_a_HPC2_and_a_reg;
  wire   [1:0] cell_2118_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2118_a_HPC2_and_mul;
  wire   [1:0] cell_2119_and_out;
  wire   [1:0] cell_2119_and_in;
  wire   [1:0] cell_2119_a_HPC2_and_a_reg;
  wire   [1:0] cell_2119_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2119_a_HPC2_and_mul;
  wire   [1:0] cell_2120_and_out;
  wire   [1:0] cell_2120_and_in;
  wire   [1:0] cell_2120_a_HPC2_and_a_reg;
  wire   [1:0] cell_2120_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2120_a_HPC2_and_mul;
  wire   [1:0] cell_2121_and_out;
  wire   [1:0] cell_2121_and_in;
  wire   [1:0] cell_2121_a_HPC2_and_a_reg;
  wire   [1:0] cell_2121_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2121_a_HPC2_and_mul;
  wire   [1:0] cell_2122_and_out;
  wire   [1:0] cell_2122_and_in;
  wire   [1:0] cell_2122_a_HPC2_and_a_reg;
  wire   [1:0] cell_2122_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2122_a_HPC2_and_mul;
  wire   [1:0] cell_2123_and_out;
  wire   [1:0] cell_2123_and_in;
  wire   [1:0] cell_2123_a_HPC2_and_a_reg;
  wire   [1:0] cell_2123_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2123_a_HPC2_and_mul;
  wire   [1:0] cell_2124_and_out;
  wire   [1:0] cell_2124_and_in;
  wire   [1:0] cell_2124_a_HPC2_and_a_reg;
  wire   [1:0] cell_2124_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2124_a_HPC2_and_mul;
  wire   [1:0] cell_2125_and_out;
  wire   [1:0] cell_2125_and_in;
  wire   [1:0] cell_2125_a_HPC2_and_a_reg;
  wire   [1:0] cell_2125_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2125_a_HPC2_and_mul;
  wire   [1:0] cell_2126_and_out;
  wire   [1:0] cell_2126_and_in;
  wire   [1:0] cell_2126_a_HPC2_and_a_reg;
  wire   [1:0] cell_2126_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2126_a_HPC2_and_mul;
  wire   [1:0] cell_2127_and_out;
  wire   [1:0] cell_2127_and_in;
  wire   [1:0] cell_2127_a_HPC2_and_a_reg;
  wire   [1:0] cell_2127_a_HPC2_and_mul_s1_out;
  wire   [1:0] cell_2127_a_HPC2_and_mul;

  DFF_X1 cell_33 ( .D(signal_429), .CK(signal_4640), .Q(), .QN(n273) );
  DFF_X1 cell_36 ( .D(signal_431), .CK(signal_4640), .Q(n265), .QN() );
  DFF_X1 cell_39 ( .D(signal_433), .CK(signal_4640), .Q(n267), .QN() );
  DFF_X1 cell_42 ( .D(signal_435), .CK(signal_4640), .Q(n266), .QN() );
  DFF_X1 cell_45 ( .D(signal_437), .CK(signal_4640), .Q(), .QN(n279) );
  DFF_X1 cell_48 ( .D(signal_439), .CK(signal_4640), .Q(signal_421), .QN(n278)
         );
  DFF_X1 cell_51 ( .D(signal_441), .CK(signal_4640), .Q(signal_420), .QN() );
  DFF_X1 cell_53 ( .D(signal_419), .CK(signal_4640), .Q(signal_418), .QN() );
  DFF_X1 cell_55 ( .D(n340), .CK(signal_4640), .Q(), .QN(n268) );
  DFF_X1 cell_1561 ( .D(signal_1275), .CK(signal_4640), .Q(signal_1268), .QN(
        n270) );
  DFF_X1 cell_1563 ( .D(signal_1266), .CK(signal_4640), .Q(signal_1269), .QN(
        n276) );
  DFF_X1 cell_1565 ( .D(signal_1264), .CK(signal_4640), .Q(signal_1270), .QN(
        n269) );
  DFF_X1 cell_1567 ( .D(signal_1262), .CK(signal_4640), .Q(signal_1271), .QN(
        n277) );
  DFF_X1 cell_1569 ( .D(signal_1260), .CK(signal_4640), .Q(signal_1272), .QN(
        n275) );
  DFF_X1 cell_1571 ( .D(signal_1259), .CK(signal_4640), .Q(signal_1273), .QN(
        n271) );
  DFF_X1 cell_1573 ( .D(signal_1258), .CK(signal_4640), .Q(signal_1274), .QN(
        n274) );
  DFF_X1 cell_1575 ( .D(signal_1256), .CK(signal_4640), .Q(signal_1254), .QN(
        n272) );
  DFF_X1 cell_1713 ( .D(n253), .CK(signal_4640), .Q(n35), .QN(n42) );
  BUF_X4 U113 ( .A(signal_1987), .Z(n380) );
  BUF_X4 U114 ( .A(signal_3261), .Z(n381) );
  BUF_X4 U115 ( .A(signal_1999), .Z(n366) );
  BUF_X4 U116 ( .A(signal_3413), .Z(n367) );
  BUF_X4 U117 ( .A(signal_1982), .Z(n388) );
  BUF_X4 U118 ( .A(signal_3256), .Z(n389) );
  INV_X1 U119 ( .A(n487), .ZN(n242) );
  BUF_X1 U120 ( .A(n29), .Z(n347) );
  BUF_X1 U121 ( .A(n29), .Z(n344) );
  BUF_X1 U122 ( .A(signal_3407), .Z(n379) );
  BUF_X1 U123 ( .A(signal_1993), .Z(n377) );
  BUF_X1 U124 ( .A(signal_1996), .Z(n373) );
  BUF_X1 U125 ( .A(signal_3410), .Z(n375) );
  BUF_X1 U126 ( .A(n309), .Z(n314) );
  BUF_X1 U127 ( .A(n29), .Z(n340) );
  BUF_X1 U128 ( .A(signal_3424), .Z(n360) );
  BUF_X1 U129 ( .A(signal_2010), .Z(n358) );
  BUF_X1 U130 ( .A(signal_2015), .Z(n353) );
  BUF_X1 U131 ( .A(signal_3429), .Z(n355) );
  BUF_X1 U132 ( .A(signal_3414), .Z(n365) );
  BUF_X1 U133 ( .A(signal_2000), .Z(n363) );
  BUF_X1 U134 ( .A(signal_1514), .Z(n441) );
  BUF_X1 U135 ( .A(signal_3235), .Z(n455) );
  BUF_X1 U136 ( .A(n242), .Z(n307) );
  BUF_X1 U137 ( .A(n242), .Z(n309) );
  BUF_X1 U138 ( .A(signal_2015), .Z(n352) );
  BUF_X1 U139 ( .A(n242), .Z(n319) );
  BUF_X1 U140 ( .A(signal_3429), .Z(n354) );
  BUF_X1 U141 ( .A(signal_1996), .Z(n372) );
  BUF_X1 U142 ( .A(n242), .Z(n317) );
  BUF_X1 U143 ( .A(signal_3410), .Z(n374) );
  BUF_X1 U144 ( .A(n29), .Z(n351) );
  BUF_X1 U145 ( .A(n242), .Z(n308) );
  BUF_X1 U146 ( .A(n344), .Z(n341) );
  BUF_X1 U147 ( .A(n344), .Z(n342) );
  BUF_X1 U148 ( .A(n285), .Z(n296) );
  BUF_X1 U149 ( .A(n284), .Z(n300) );
  BUF_X1 U150 ( .A(n284), .Z(n304) );
  BUF_X1 U151 ( .A(n286), .Z(n295) );
  BUF_X1 U152 ( .A(n284), .Z(n297) );
  INV_X1 U153 ( .A(n343), .ZN(n331) );
  INV_X1 U154 ( .A(n348), .ZN(n337) );
  BUF_X1 U155 ( .A(n348), .Z(n350) );
  BUF_X1 U156 ( .A(n344), .Z(n349) );
  BUF_X1 U157 ( .A(n343), .Z(n345) );
  BUF_X1 U158 ( .A(n286), .Z(n302) );
  BUF_X1 U159 ( .A(n285), .Z(n306) );
  BUF_X1 U160 ( .A(n285), .Z(n301) );
  BUF_X1 U161 ( .A(n35), .Z(n285) );
  BUF_X2 U162 ( .A(signal_1511), .Z(n392) );
  BUF_X2 U163 ( .A(signal_3238), .Z(n393) );
  BUF_X1 U164 ( .A(n282), .Z(n293) );
  BUF_X1 U165 ( .A(signal_3235), .Z(n442) );
  BUF_X1 U166 ( .A(signal_1514), .Z(n428) );
  BUF_X1 U167 ( .A(n281), .Z(n287) );
  INV_X1 U168 ( .A(n347), .ZN(n330) );
  BUF_X1 U169 ( .A(n283), .Z(n289) );
  INV_X1 U170 ( .A(n348), .ZN(n328) );
  INV_X1 U171 ( .A(n339), .ZN(n334) );
  INV_X1 U172 ( .A(n343), .ZN(n327) );
  BUF_X1 U173 ( .A(n29), .Z(n343) );
  BUF_X1 U174 ( .A(n281), .Z(n290) );
  BUF_X1 U175 ( .A(n282), .Z(n291) );
  INV_X1 U176 ( .A(n347), .ZN(n326) );
  INV_X1 U177 ( .A(n340), .ZN(n329) );
  BUF_X1 U178 ( .A(n282), .Z(n288) );
  BUF_X1 U179 ( .A(n317), .Z(n322) );
  INV_X1 U180 ( .A(n340), .ZN(n335) );
  BUF_X1 U181 ( .A(n319), .Z(n313) );
  BUF_X1 U182 ( .A(n309), .Z(n312) );
  INV_X1 U183 ( .A(n344), .ZN(n325) );
  BUF_X1 U184 ( .A(n316), .Z(n320) );
  INV_X1 U185 ( .A(n348), .ZN(n336) );
  BUF_X1 U186 ( .A(n29), .Z(n348) );
  INV_X1 U187 ( .A(n347), .ZN(n324) );
  BUF_X1 U188 ( .A(n309), .Z(n311) );
  BUF_X1 U189 ( .A(n281), .Z(n294) );
  BUF_X1 U190 ( .A(signal_1514), .Z(n434) );
  BUF_X1 U191 ( .A(signal_3235), .Z(n448) );
  INV_X1 U192 ( .A(n344), .ZN(n332) );
  INV_X1 U193 ( .A(n340), .ZN(n333) );
  BUF_X1 U194 ( .A(n35), .Z(n284) );
  BUF_X1 U195 ( .A(n283), .Z(n299) );
  BUF_X1 U196 ( .A(n286), .Z(n298) );
  BUF_X1 U197 ( .A(n35), .Z(n286) );
  BUF_X1 U198 ( .A(signal_1514), .Z(n438) );
  BUF_X1 U199 ( .A(signal_3235), .Z(n452) );
  BUF_X1 U200 ( .A(signal_3237), .Z(n413) );
  BUF_X1 U201 ( .A(signal_1512), .Z(n396) );
  BUF_X1 U202 ( .A(signal_3237), .Z(n427) );
  BUF_X1 U203 ( .A(signal_1512), .Z(n410) );
  BUF_X1 U204 ( .A(signal_3237), .Z(n412) );
  BUF_X1 U205 ( .A(signal_1512), .Z(n395) );
  BUF_X1 U206 ( .A(signal_1512), .Z(n407) );
  BUF_X1 U207 ( .A(signal_3237), .Z(n424) );
  BUF_X1 U208 ( .A(signal_1512), .Z(n408) );
  BUF_X1 U209 ( .A(signal_3237), .Z(n425) );
  BUF_X1 U210 ( .A(signal_1512), .Z(n409) );
  BUF_X1 U211 ( .A(signal_3237), .Z(n426) );
  BUF_X1 U212 ( .A(signal_3237), .Z(n411) );
  BUF_X1 U213 ( .A(signal_1512), .Z(n394) );
  BUF_X1 U214 ( .A(signal_3237), .Z(n416) );
  BUF_X1 U215 ( .A(signal_1512), .Z(n399) );
  BUF_X1 U216 ( .A(signal_1512), .Z(n400) );
  BUF_X1 U217 ( .A(signal_3237), .Z(n417) );
  BUF_X1 U218 ( .A(signal_3237), .Z(n421) );
  BUF_X1 U219 ( .A(signal_1512), .Z(n404) );
  BUF_X1 U220 ( .A(signal_1512), .Z(n401) );
  BUF_X1 U221 ( .A(signal_3237), .Z(n418) );
  BUF_X1 U222 ( .A(signal_3237), .Z(n420) );
  BUF_X1 U223 ( .A(signal_1512), .Z(n403) );
  BUF_X1 U224 ( .A(signal_1512), .Z(n402) );
  BUF_X1 U225 ( .A(signal_3237), .Z(n419) );
  BUF_X1 U226 ( .A(signal_1512), .Z(n397) );
  BUF_X1 U227 ( .A(signal_3237), .Z(n414) );
  BUF_X1 U228 ( .A(signal_3237), .Z(n423) );
  BUF_X1 U229 ( .A(signal_1512), .Z(n406) );
  BUF_X1 U230 ( .A(signal_3411), .Z(n371) );
  BUF_X1 U231 ( .A(signal_1997), .Z(n369) );
  BUF_X1 U232 ( .A(signal_1512), .Z(n405) );
  BUF_X1 U233 ( .A(signal_3237), .Z(n415) );
  BUF_X1 U234 ( .A(signal_3237), .Z(n422) );
  BUF_X1 U235 ( .A(signal_1512), .Z(n398) );
  BUF_X1 U236 ( .A(signal_1514), .Z(n437) );
  BUF_X1 U237 ( .A(signal_3235), .Z(n451) );
  BUF_X1 U238 ( .A(signal_1514), .Z(n430) );
  BUF_X1 U239 ( .A(signal_3235), .Z(n444) );
  BUF_X1 U240 ( .A(signal_1514), .Z(n429) );
  BUF_X1 U241 ( .A(signal_3235), .Z(n445) );
  BUF_X1 U242 ( .A(signal_3235), .Z(n443) );
  BUF_X1 U243 ( .A(signal_1514), .Z(n431) );
  BUF_X1 U244 ( .A(n340), .Z(n338) );
  BUF_X1 U245 ( .A(signal_1514), .Z(n432) );
  BUF_X1 U246 ( .A(signal_3235), .Z(n446) );
  BUF_X1 U247 ( .A(n455), .Z(n454) );
  BUF_X1 U248 ( .A(n309), .Z(n318) );
  BUF_X1 U249 ( .A(n441), .Z(n439) );
  BUF_X1 U250 ( .A(n441), .Z(n440) );
  BUF_X1 U251 ( .A(n455), .Z(n453) );
  BUF_X2 U252 ( .A(signal_1516), .Z(n465) );
  BUF_X2 U253 ( .A(signal_3233), .Z(n469) );
  BUF_X1 U254 ( .A(signal_3411), .Z(n370) );
  BUF_X1 U255 ( .A(signal_1997), .Z(n368) );
  BUF_X2 U256 ( .A(signal_1516), .Z(n463) );
  BUF_X2 U257 ( .A(signal_3233), .Z(n467) );
  BUF_X1 U258 ( .A(signal_3235), .Z(n449) );
  BUF_X1 U259 ( .A(signal_1514), .Z(n436) );
  BUF_X1 U260 ( .A(signal_3235), .Z(n450) );
  BUF_X1 U261 ( .A(signal_1514), .Z(n435) );
  BUF_X1 U262 ( .A(signal_3235), .Z(n447) );
  BUF_X1 U263 ( .A(signal_1514), .Z(n433) );
  BUF_X1 U264 ( .A(signal_2010), .Z(n359) );
  BUF_X1 U265 ( .A(signal_3424), .Z(n361) );
  BUF_X1 U266 ( .A(signal_1515), .Z(n458) );
  BUF_X1 U267 ( .A(signal_3234), .Z(n461) );
  BUF_X2 U268 ( .A(signal_1516), .Z(n462) );
  BUF_X1 U269 ( .A(signal_1993), .Z(n376) );
  BUF_X2 U270 ( .A(signal_3233), .Z(n466) );
  BUF_X1 U271 ( .A(signal_3407), .Z(n378) );
  BUF_X1 U272 ( .A(signal_1515), .Z(n456) );
  BUF_X2 U273 ( .A(signal_1516), .Z(n464) );
  BUF_X1 U274 ( .A(signal_3234), .Z(n459) );
  BUF_X2 U275 ( .A(signal_3233), .Z(n468) );
  BUF_X1 U276 ( .A(signal_3239), .Z(n391) );
  BUF_X2 U277 ( .A(signal_3427), .Z(n357) );
  BUF_X1 U278 ( .A(signal_1510), .Z(n390) );
  BUF_X2 U279 ( .A(signal_2013), .Z(n356) );
  BUF_X1 U280 ( .A(signal_3234), .Z(n460) );
  BUF_X1 U281 ( .A(signal_1515), .Z(n457) );
  BUF_X1 U282 ( .A(signal_1983), .Z(n385) );
  BUF_X1 U283 ( .A(signal_3257), .Z(n387) );
  BUF_X1 U284 ( .A(signal_3414), .Z(n364) );
  BUF_X1 U285 ( .A(signal_2000), .Z(n362) );
  BUF_X1 U286 ( .A(n242), .Z(n321) );
  BUF_X1 U287 ( .A(signal_399), .Z(n471) );
  BUF_X1 U288 ( .A(signal_3257), .Z(n386) );
  BUF_X1 U289 ( .A(signal_1983), .Z(n384) );
  BUF_X2 U290 ( .A(signal_1984), .Z(n382) );
  BUF_X2 U291 ( .A(signal_3258), .Z(n383) );
  BUF_X1 U292 ( .A(n29), .Z(n339) );
  BUF_X1 U293 ( .A(n242), .Z(n315) );
  BUF_X1 U294 ( .A(signal_399), .Z(n472) );
  BUF_X1 U295 ( .A(n242), .Z(n310) );
  BUF_X1 U296 ( .A(n283), .Z(n292) );
  BUF_X1 U297 ( .A(n308), .Z(n323) );
  BUF_X1 U298 ( .A(signal_399), .Z(n470) );
  BUF_X1 U299 ( .A(signal_399), .Z(n473) );
  INV_X1 U300 ( .A(n474), .ZN(signal_399) );
  NOR2_X1 U301 ( .A1(n42), .A2(n475), .ZN(n29) );
  OR4_X1 U302 ( .A1(n265), .A2(n267), .A3(n266), .A4(n484), .ZN(n475) );
  BUF_X1 U303 ( .A(n242), .Z(n316) );
  NAND2_X1 U304 ( .A1(signal_418), .A2(n280), .ZN(n487) );
  BUF_X1 U305 ( .A(n35), .Z(n280) );
  BUF_X1 U306 ( .A(n35), .Z(n303) );
  BUF_X1 U307 ( .A(n35), .Z(n305) );
  AOI211_X4 U308 ( .C1(n482), .C2(n481), .A(n42), .B(n483), .ZN(signal_400) );
  BUF_X1 U309 ( .A(n35), .Z(n282) );
  BUF_X1 U310 ( .A(n35), .Z(n281) );
  BUF_X1 U311 ( .A(n35), .Z(n283) );
  NAND2_X1 U312 ( .A1(n273), .A2(n279), .ZN(n484) );
  BUF_X1 U313 ( .A(n29), .Z(n346) );
  NAND4_X1 U314 ( .A1(signal_1272), .A2(signal_1270), .A3(signal_1269), .A4(
        signal_1273), .ZN(n474) );
  NOR4_X1 U315 ( .A1(signal_420), .A2(n278), .A3(n336), .A4(n474), .ZN(done)
         );
  OAI221_X1 U316 ( .B1(n343), .B2(n272), .C1(n337), .C2(n274), .A(n280), .ZN(
        signal_1256) );
  NAND2_X1 U317 ( .A1(n283), .A2(n475), .ZN(n486) );
  OAI22_X1 U318 ( .A1(n337), .A2(n271), .B1(n486), .B2(n274), .ZN(signal_1258)
         );
  OAI22_X1 U319 ( .A1(n336), .A2(n275), .B1(n486), .B2(n271), .ZN(signal_1259)
         );
  NAND2_X1 U320 ( .A1(n347), .A2(signal_1254), .ZN(n480) );
  NOR2_X1 U321 ( .A1(signal_1254), .A2(n325), .ZN(n478) );
  INV_X1 U322 ( .A(n486), .ZN(n485) );
  AOI22_X1 U323 ( .A1(signal_1271), .A2(n478), .B1(n485), .B2(signal_1272), 
        .ZN(n476) );
  OAI21_X1 U324 ( .B1(signal_1271), .B2(n480), .A(n476), .ZN(signal_1260) );
  AOI22_X1 U325 ( .A1(signal_1271), .A2(n332), .B1(n478), .B2(signal_1270), 
        .ZN(n477) );
  OAI211_X1 U326 ( .C1(signal_1270), .C2(n480), .A(n477), .B(n294), .ZN(
        signal_1262) );
  OAI221_X1 U327 ( .B1(n339), .B2(n269), .C1(n328), .C2(n276), .A(n298), .ZN(
        signal_1264) );
  AOI22_X1 U328 ( .A1(n478), .A2(signal_1268), .B1(n485), .B2(signal_1269), 
        .ZN(n479) );
  OAI21_X1 U329 ( .B1(signal_1268), .B2(n480), .A(n479), .ZN(signal_1266) );
  OAI211_X1 U330 ( .C1(n347), .C2(n270), .A(n291), .B(n480), .ZN(signal_1275)
         );
  NOR2_X1 U331 ( .A1(n272), .A2(n268), .ZN(signal_1494) );
  NOR2_X1 U332 ( .A1(n274), .A2(n268), .ZN(signal_1495) );
  NOR2_X1 U333 ( .A1(n271), .A2(n268), .ZN(signal_1496) );
  NOR2_X1 U334 ( .A1(n275), .A2(n268), .ZN(signal_1497) );
  NOR2_X1 U335 ( .A1(n277), .A2(n268), .ZN(signal_1498) );
  NOR2_X1 U336 ( .A1(n269), .A2(n268), .ZN(signal_1499) );
  NOR2_X1 U337 ( .A1(n276), .A2(n268), .ZN(signal_1500) );
  NOR2_X1 U338 ( .A1(n270), .A2(n268), .ZN(signal_1501) );
  NOR4_X1 U339 ( .A1(n277), .A2(n272), .A3(n269), .A4(n270), .ZN(n482) );
  NOR4_X1 U340 ( .A1(signal_1272), .A2(signal_1269), .A3(signal_1274), .A4(
        signal_1273), .ZN(n481) );
  NOR2_X1 U341 ( .A1(signal_421), .A2(signal_420), .ZN(n483) );
  OAI21_X1 U342 ( .B1(n483), .B2(n487), .A(n328), .ZN(signal_419) );
  OAI211_X1 U343 ( .C1(n273), .C2(n279), .A(n299), .B(n484), .ZN(signal_429)
         );
  NOR2_X1 U344 ( .A1(n42), .A2(n273), .ZN(signal_431) );
  OR2_X1 U345 ( .A1(n42), .A2(n265), .ZN(signal_433) );
  AND2_X1 U346 ( .A1(n267), .A2(n290), .ZN(signal_435) );
  OR2_X1 U347 ( .A1(n42), .A2(n266), .ZN(signal_437) );
  NAND2_X1 U348 ( .A1(n485), .A2(signal_420), .ZN(signal_439) );
  NOR2_X1 U349 ( .A1(n486), .A2(n278), .ZN(signal_441) );
  INV_X1 U350 ( .A(start), .ZN(n253) );
  XOR2_X1 cell_1_Ins_0_U1 ( .A(ciphertext_s0[120]), .B(signal_1493), .Z(
        signal_1413) );
  XOR2_X1 cell_1_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(signal_2389), .Z(
        signal_2390) );
  XOR2_X1 cell_2_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(signal_1492), .Z(
        signal_1412) );
  XOR2_X1 cell_2_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(signal_2392), .Z(
        signal_2393) );
  XOR2_X1 cell_3_Ins_0_U1 ( .A(ciphertext_s0[122]), .B(signal_1491), .Z(
        signal_1411) );
  XOR2_X1 cell_3_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(signal_2395), .Z(
        signal_2396) );
  XOR2_X1 cell_4_Ins_0_U1 ( .A(ciphertext_s0[123]), .B(signal_1490), .Z(
        signal_1410) );
  XOR2_X1 cell_4_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(signal_2398), .Z(
        signal_2399) );
  XOR2_X1 cell_5_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(signal_1489), .Z(
        signal_1409) );
  XOR2_X1 cell_5_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(signal_2401), .Z(
        signal_2402) );
  XOR2_X1 cell_6_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(signal_1488), .Z(
        signal_1408) );
  XOR2_X1 cell_6_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(signal_2404), .Z(
        signal_2405) );
  XOR2_X1 cell_7_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(signal_1487), .Z(
        signal_1407) );
  XOR2_X1 cell_7_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(signal_2407), .Z(
        signal_2408) );
  XOR2_X1 cell_8_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(signal_1486), .Z(
        signal_1406) );
  XOR2_X1 cell_8_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(signal_2410), .Z(
        signal_2411) );
  MUX2_X1 cell_85_Ins_0_U1 ( .A(signal_1677), .B(ciphertext_s0[120]), .S(n338), 
        .Z(signal_465) );
  MUX2_X1 cell_85_Ins_1_U1 ( .A(signal_2562), .B(ciphertext_s1[120]), .S(n338), 
        .Z(signal_3786) );
  MUX2_X1 cell_88_Ins_0_U1 ( .A(signal_1676), .B(ciphertext_s0[121]), .S(n348), 
        .Z(signal_467) );
  MUX2_X1 cell_88_Ins_1_U1 ( .A(signal_2565), .B(ciphertext_s1[121]), .S(n348), 
        .Z(signal_3787) );
  MUX2_X1 cell_91_Ins_0_U1 ( .A(signal_1675), .B(ciphertext_s0[122]), .S(n340), 
        .Z(signal_469) );
  MUX2_X1 cell_91_Ins_1_U1 ( .A(signal_2568), .B(ciphertext_s1[122]), .S(n340), 
        .Z(signal_3788) );
  MUX2_X1 cell_94_Ins_0_U1 ( .A(signal_1674), .B(ciphertext_s0[123]), .S(n339), 
        .Z(signal_471) );
  MUX2_X1 cell_94_Ins_1_U1 ( .A(signal_2571), .B(ciphertext_s1[123]), .S(n339), 
        .Z(signal_3789) );
  MUX2_X1 cell_97_Ins_0_U1 ( .A(signal_1673), .B(ciphertext_s0[124]), .S(n344), 
        .Z(signal_473) );
  MUX2_X1 cell_97_Ins_1_U1 ( .A(signal_2574), .B(ciphertext_s1[124]), .S(n344), 
        .Z(signal_3790) );
  MUX2_X1 cell_100_Ins_0_U1 ( .A(signal_1672), .B(ciphertext_s0[125]), .S(n347), .Z(signal_475) );
  MUX2_X1 cell_100_Ins_1_U1 ( .A(signal_2577), .B(ciphertext_s1[125]), .S(n347), .Z(signal_3791) );
  MUX2_X1 cell_103_Ins_0_U1 ( .A(signal_1671), .B(ciphertext_s0[126]), .S(n348), .Z(signal_477) );
  MUX2_X1 cell_103_Ins_1_U1 ( .A(signal_2580), .B(ciphertext_s1[126]), .S(n348), .Z(signal_3792) );
  MUX2_X1 cell_106_Ins_0_U1 ( .A(signal_1670), .B(ciphertext_s0[127]), .S(n343), .Z(signal_479) );
  MUX2_X1 cell_106_Ins_1_U1 ( .A(signal_2583), .B(ciphertext_s1[127]), .S(n343), .Z(signal_3793) );
  MUX2_X1 cell_109_Ins_0_U1 ( .A(signal_1669), .B(ciphertext_s0[112]), .S(n347), .Z(signal_481) );
  MUX2_X1 cell_109_Ins_1_U1 ( .A(signal_2586), .B(ciphertext_s1[112]), .S(n347), .Z(signal_3794) );
  MUX2_X1 cell_112_Ins_0_U1 ( .A(signal_1668), .B(ciphertext_s0[113]), .S(n343), .Z(signal_483) );
  MUX2_X1 cell_112_Ins_1_U1 ( .A(signal_2589), .B(ciphertext_s1[113]), .S(n343), .Z(signal_3795) );
  MUX2_X1 cell_115_Ins_0_U1 ( .A(signal_1667), .B(ciphertext_s0[114]), .S(n339), .Z(signal_485) );
  MUX2_X1 cell_115_Ins_1_U1 ( .A(signal_2592), .B(ciphertext_s1[114]), .S(n339), .Z(signal_3796) );
  MUX2_X1 cell_118_Ins_0_U1 ( .A(signal_1666), .B(ciphertext_s0[115]), .S(n343), .Z(signal_487) );
  MUX2_X1 cell_118_Ins_1_U1 ( .A(signal_2595), .B(ciphertext_s1[115]), .S(n343), .Z(signal_3797) );
  MUX2_X1 cell_121_Ins_0_U1 ( .A(signal_1665), .B(ciphertext_s0[116]), .S(n349), .Z(signal_489) );
  MUX2_X1 cell_121_Ins_1_U1 ( .A(signal_2598), .B(ciphertext_s1[116]), .S(n349), .Z(signal_3798) );
  MUX2_X1 cell_124_Ins_0_U1 ( .A(signal_1664), .B(ciphertext_s0[117]), .S(n348), .Z(signal_491) );
  MUX2_X1 cell_124_Ins_1_U1 ( .A(signal_2601), .B(ciphertext_s1[117]), .S(n348), .Z(signal_3799) );
  MUX2_X1 cell_127_Ins_0_U1 ( .A(signal_1663), .B(ciphertext_s0[118]), .S(n340), .Z(signal_493) );
  MUX2_X1 cell_127_Ins_1_U1 ( .A(signal_2604), .B(ciphertext_s1[118]), .S(n340), .Z(signal_3800) );
  MUX2_X1 cell_130_Ins_0_U1 ( .A(signal_1662), .B(ciphertext_s0[119]), .S(n344), .Z(signal_495) );
  MUX2_X1 cell_130_Ins_1_U1 ( .A(signal_2607), .B(ciphertext_s1[119]), .S(n344), .Z(signal_3801) );
  MUX2_X1 cell_133_Ins_0_U1 ( .A(signal_1661), .B(ciphertext_s0[104]), .S(n339), .Z(signal_497) );
  MUX2_X1 cell_133_Ins_1_U1 ( .A(signal_2610), .B(ciphertext_s1[104]), .S(n339), .Z(signal_3802) );
  MUX2_X1 cell_136_Ins_0_U1 ( .A(signal_1660), .B(ciphertext_s0[105]), .S(n343), .Z(signal_499) );
  MUX2_X1 cell_136_Ins_1_U1 ( .A(signal_2613), .B(ciphertext_s1[105]), .S(n343), .Z(signal_3803) );
  MUX2_X1 cell_139_Ins_0_U1 ( .A(signal_1659), .B(ciphertext_s0[106]), .S(n347), .Z(signal_501) );
  MUX2_X1 cell_139_Ins_1_U1 ( .A(signal_2616), .B(ciphertext_s1[106]), .S(n347), .Z(signal_3804) );
  MUX2_X1 cell_142_Ins_0_U1 ( .A(signal_1658), .B(ciphertext_s0[107]), .S(n344), .Z(signal_503) );
  MUX2_X1 cell_142_Ins_1_U1 ( .A(signal_2619), .B(ciphertext_s1[107]), .S(n344), .Z(signal_3805) );
  MUX2_X1 cell_145_Ins_0_U1 ( .A(signal_1657), .B(ciphertext_s0[108]), .S(n347), .Z(signal_505) );
  MUX2_X1 cell_145_Ins_1_U1 ( .A(signal_2622), .B(ciphertext_s1[108]), .S(n347), .Z(signal_3806) );
  MUX2_X1 cell_148_Ins_0_U1 ( .A(signal_1656), .B(ciphertext_s0[109]), .S(n339), .Z(signal_507) );
  MUX2_X1 cell_148_Ins_1_U1 ( .A(signal_2625), .B(ciphertext_s1[109]), .S(n339), .Z(signal_3807) );
  MUX2_X1 cell_151_Ins_0_U1 ( .A(signal_1655), .B(ciphertext_s0[110]), .S(n340), .Z(signal_509) );
  MUX2_X1 cell_151_Ins_1_U1 ( .A(signal_2628), .B(ciphertext_s1[110]), .S(n340), .Z(signal_3808) );
  MUX2_X1 cell_154_Ins_0_U1 ( .A(signal_1654), .B(ciphertext_s0[111]), .S(n348), .Z(signal_511) );
  MUX2_X1 cell_154_Ins_1_U1 ( .A(signal_2631), .B(ciphertext_s1[111]), .S(n348), .Z(signal_3809) );
  MUX2_X1 cell_157_Ins_0_U1 ( .A(signal_1653), .B(ciphertext_s0[96]), .S(n346), 
        .Z(signal_513) );
  MUX2_X1 cell_157_Ins_1_U1 ( .A(signal_3592), .B(ciphertext_s1[96]), .S(n346), 
        .Z(signal_3810) );
  MUX2_X1 cell_160_Ins_0_U1 ( .A(signal_1652), .B(ciphertext_s0[97]), .S(n343), 
        .Z(signal_515) );
  MUX2_X1 cell_160_Ins_1_U1 ( .A(signal_3594), .B(ciphertext_s1[97]), .S(n343), 
        .Z(signal_3811) );
  MUX2_X1 cell_163_Ins_0_U1 ( .A(signal_1651), .B(ciphertext_s0[98]), .S(n345), 
        .Z(signal_517) );
  MUX2_X1 cell_163_Ins_1_U1 ( .A(signal_3596), .B(ciphertext_s1[98]), .S(n345), 
        .Z(signal_3812) );
  MUX2_X1 cell_166_Ins_0_U1 ( .A(signal_1650), .B(ciphertext_s0[99]), .S(n350), 
        .Z(signal_519) );
  MUX2_X1 cell_166_Ins_1_U1 ( .A(signal_3598), .B(ciphertext_s1[99]), .S(n350), 
        .Z(signal_3813) );
  MUX2_X1 cell_169_Ins_0_U1 ( .A(signal_1649), .B(ciphertext_s0[100]), .S(n351), .Z(signal_521) );
  MUX2_X1 cell_169_Ins_1_U1 ( .A(signal_3600), .B(ciphertext_s1[100]), .S(n351), .Z(signal_3814) );
  MUX2_X1 cell_172_Ins_0_U1 ( .A(signal_1648), .B(ciphertext_s0[101]), .S(n339), .Z(signal_523) );
  MUX2_X1 cell_172_Ins_1_U1 ( .A(signal_3602), .B(ciphertext_s1[101]), .S(n339), .Z(signal_3815) );
  MUX2_X1 cell_175_Ins_0_U1 ( .A(signal_1647), .B(ciphertext_s0[102]), .S(n351), .Z(signal_525) );
  MUX2_X1 cell_175_Ins_1_U1 ( .A(signal_3604), .B(ciphertext_s1[102]), .S(n351), .Z(signal_3816) );
  MUX2_X1 cell_178_Ins_0_U1 ( .A(signal_1646), .B(ciphertext_s0[103]), .S(n346), .Z(signal_527) );
  MUX2_X1 cell_178_Ins_1_U1 ( .A(signal_3606), .B(ciphertext_s1[103]), .S(n346), .Z(signal_3817) );
  MUX2_X1 cell_181_Ins_0_U1 ( .A(signal_1645), .B(ciphertext_s0[80]), .S(n351), 
        .Z(signal_529) );
  MUX2_X1 cell_181_Ins_1_U1 ( .A(signal_2634), .B(ciphertext_s1[80]), .S(n351), 
        .Z(signal_3818) );
  MUX2_X1 cell_184_Ins_0_U1 ( .A(signal_1644), .B(ciphertext_s0[81]), .S(n345), 
        .Z(signal_531) );
  MUX2_X1 cell_184_Ins_1_U1 ( .A(signal_2637), .B(ciphertext_s1[81]), .S(n345), 
        .Z(signal_3819) );
  MUX2_X1 cell_187_Ins_0_U1 ( .A(signal_1643), .B(ciphertext_s0[82]), .S(n351), 
        .Z(signal_533) );
  MUX2_X1 cell_187_Ins_1_U1 ( .A(signal_2640), .B(ciphertext_s1[82]), .S(n351), 
        .Z(signal_3820) );
  MUX2_X1 cell_190_Ins_0_U1 ( .A(signal_1642), .B(ciphertext_s0[83]), .S(n346), 
        .Z(signal_535) );
  MUX2_X1 cell_190_Ins_1_U1 ( .A(signal_2643), .B(ciphertext_s1[83]), .S(n346), 
        .Z(signal_3821) );
  MUX2_X1 cell_193_Ins_0_U1 ( .A(signal_1641), .B(ciphertext_s0[84]), .S(n346), 
        .Z(signal_537) );
  MUX2_X1 cell_193_Ins_1_U1 ( .A(signal_2646), .B(ciphertext_s1[84]), .S(n346), 
        .Z(signal_3822) );
  MUX2_X1 cell_196_Ins_0_U1 ( .A(signal_1640), .B(ciphertext_s0[85]), .S(n338), 
        .Z(signal_539) );
  MUX2_X1 cell_196_Ins_1_U1 ( .A(signal_2649), .B(ciphertext_s1[85]), .S(n338), 
        .Z(signal_3823) );
  MUX2_X1 cell_199_Ins_0_U1 ( .A(signal_1639), .B(ciphertext_s0[86]), .S(n346), 
        .Z(signal_541) );
  MUX2_X1 cell_199_Ins_1_U1 ( .A(signal_2652), .B(ciphertext_s1[86]), .S(n346), 
        .Z(signal_3824) );
  MUX2_X1 cell_202_Ins_0_U1 ( .A(signal_1638), .B(ciphertext_s0[87]), .S(n346), 
        .Z(signal_543) );
  MUX2_X1 cell_202_Ins_1_U1 ( .A(signal_2655), .B(ciphertext_s1[87]), .S(n346), 
        .Z(signal_3825) );
  MUX2_X1 cell_205_Ins_0_U1 ( .A(signal_1637), .B(ciphertext_s0[72]), .S(n351), 
        .Z(signal_545) );
  MUX2_X1 cell_205_Ins_1_U1 ( .A(signal_2658), .B(ciphertext_s1[72]), .S(n351), 
        .Z(signal_3826) );
  MUX2_X1 cell_208_Ins_0_U1 ( .A(signal_1636), .B(ciphertext_s0[73]), .S(n349), 
        .Z(signal_547) );
  MUX2_X1 cell_208_Ins_1_U1 ( .A(signal_2661), .B(ciphertext_s1[73]), .S(n349), 
        .Z(signal_3827) );
  MUX2_X1 cell_211_Ins_0_U1 ( .A(signal_1635), .B(ciphertext_s0[74]), .S(n351), 
        .Z(signal_549) );
  MUX2_X1 cell_211_Ins_1_U1 ( .A(signal_2664), .B(ciphertext_s1[74]), .S(n351), 
        .Z(signal_3828) );
  MUX2_X1 cell_214_Ins_0_U1 ( .A(signal_1634), .B(ciphertext_s0[75]), .S(n351), 
        .Z(signal_551) );
  MUX2_X1 cell_214_Ins_1_U1 ( .A(signal_2667), .B(ciphertext_s1[75]), .S(n351), 
        .Z(signal_3829) );
  MUX2_X1 cell_217_Ins_0_U1 ( .A(signal_1633), .B(ciphertext_s0[76]), .S(n346), 
        .Z(signal_553) );
  MUX2_X1 cell_217_Ins_1_U1 ( .A(signal_2670), .B(ciphertext_s1[76]), .S(n346), 
        .Z(signal_3830) );
  MUX2_X1 cell_220_Ins_0_U1 ( .A(signal_1632), .B(ciphertext_s0[77]), .S(n338), 
        .Z(signal_555) );
  MUX2_X1 cell_220_Ins_1_U1 ( .A(signal_2673), .B(ciphertext_s1[77]), .S(n338), 
        .Z(signal_3831) );
  MUX2_X1 cell_223_Ins_0_U1 ( .A(signal_1631), .B(ciphertext_s0[78]), .S(n351), 
        .Z(signal_557) );
  MUX2_X1 cell_223_Ins_1_U1 ( .A(signal_2676), .B(ciphertext_s1[78]), .S(n351), 
        .Z(signal_3832) );
  MUX2_X1 cell_226_Ins_0_U1 ( .A(signal_1630), .B(ciphertext_s0[79]), .S(n349), 
        .Z(signal_559) );
  MUX2_X1 cell_226_Ins_1_U1 ( .A(signal_2679), .B(ciphertext_s1[79]), .S(n349), 
        .Z(signal_3833) );
  MUX2_X1 cell_229_Ins_0_U1 ( .A(signal_1629), .B(ciphertext_s0[64]), .S(n351), 
        .Z(signal_561) );
  MUX2_X1 cell_229_Ins_1_U1 ( .A(signal_2682), .B(ciphertext_s1[64]), .S(n351), 
        .Z(signal_3834) );
  MUX2_X1 cell_232_Ins_0_U1 ( .A(signal_1628), .B(ciphertext_s0[65]), .S(n351), 
        .Z(signal_563) );
  MUX2_X1 cell_232_Ins_1_U1 ( .A(signal_2685), .B(ciphertext_s1[65]), .S(n351), 
        .Z(signal_3835) );
  MUX2_X1 cell_235_Ins_0_U1 ( .A(signal_1627), .B(ciphertext_s0[66]), .S(n350), 
        .Z(signal_565) );
  MUX2_X1 cell_235_Ins_1_U1 ( .A(signal_2688), .B(ciphertext_s1[66]), .S(n350), 
        .Z(signal_3836) );
  MUX2_X1 cell_238_Ins_0_U1 ( .A(signal_1626), .B(ciphertext_s0[67]), .S(n340), 
        .Z(signal_567) );
  MUX2_X1 cell_238_Ins_1_U1 ( .A(signal_2691), .B(ciphertext_s1[67]), .S(n340), 
        .Z(signal_3837) );
  MUX2_X1 cell_241_Ins_0_U1 ( .A(signal_1625), .B(ciphertext_s0[68]), .S(n341), 
        .Z(signal_569) );
  MUX2_X1 cell_241_Ins_1_U1 ( .A(signal_2694), .B(ciphertext_s1[68]), .S(n341), 
        .Z(signal_3838) );
  MUX2_X1 cell_244_Ins_0_U1 ( .A(signal_1624), .B(ciphertext_s0[69]), .S(n342), 
        .Z(signal_571) );
  MUX2_X1 cell_244_Ins_1_U1 ( .A(signal_2697), .B(ciphertext_s1[69]), .S(n342), 
        .Z(signal_3839) );
  MUX2_X1 cell_247_Ins_0_U1 ( .A(signal_1623), .B(ciphertext_s0[70]), .S(n341), 
        .Z(signal_573) );
  MUX2_X1 cell_247_Ins_1_U1 ( .A(signal_2700), .B(ciphertext_s1[70]), .S(n341), 
        .Z(signal_3840) );
  MUX2_X1 cell_250_Ins_0_U1 ( .A(signal_1622), .B(ciphertext_s0[71]), .S(n341), 
        .Z(signal_575) );
  MUX2_X1 cell_250_Ins_1_U1 ( .A(signal_2703), .B(ciphertext_s1[71]), .S(n341), 
        .Z(signal_3841) );
  MUX2_X1 cell_253_Ins_0_U1 ( .A(signal_1621), .B(ciphertext_s0[88]), .S(n350), 
        .Z(signal_577) );
  MUX2_X1 cell_253_Ins_1_U1 ( .A(signal_3608), .B(ciphertext_s1[88]), .S(n350), 
        .Z(signal_3842) );
  MUX2_X1 cell_256_Ins_0_U1 ( .A(signal_1620), .B(ciphertext_s0[89]), .S(n341), 
        .Z(signal_579) );
  MUX2_X1 cell_256_Ins_1_U1 ( .A(signal_3610), .B(ciphertext_s1[89]), .S(n341), 
        .Z(signal_3843) );
  MUX2_X1 cell_259_Ins_0_U1 ( .A(signal_1619), .B(ciphertext_s0[90]), .S(n342), 
        .Z(signal_581) );
  MUX2_X1 cell_259_Ins_1_U1 ( .A(signal_3612), .B(ciphertext_s1[90]), .S(n342), 
        .Z(signal_3844) );
  MUX2_X1 cell_262_Ins_0_U1 ( .A(signal_1618), .B(ciphertext_s0[91]), .S(n350), 
        .Z(signal_583) );
  MUX2_X1 cell_262_Ins_1_U1 ( .A(signal_3614), .B(ciphertext_s1[91]), .S(n350), 
        .Z(signal_3845) );
  MUX2_X1 cell_265_Ins_0_U1 ( .A(signal_1617), .B(ciphertext_s0[92]), .S(n350), 
        .Z(signal_585) );
  MUX2_X1 cell_265_Ins_1_U1 ( .A(signal_3616), .B(ciphertext_s1[92]), .S(n350), 
        .Z(signal_3846) );
  MUX2_X1 cell_268_Ins_0_U1 ( .A(signal_1616), .B(ciphertext_s0[93]), .S(n350), 
        .Z(signal_587) );
  MUX2_X1 cell_268_Ins_1_U1 ( .A(signal_3618), .B(ciphertext_s1[93]), .S(n350), 
        .Z(signal_3847) );
  MUX2_X1 cell_271_Ins_0_U1 ( .A(signal_1615), .B(ciphertext_s0[94]), .S(n349), 
        .Z(signal_589) );
  MUX2_X1 cell_271_Ins_1_U1 ( .A(signal_3620), .B(ciphertext_s1[94]), .S(n349), 
        .Z(signal_3848) );
  MUX2_X1 cell_274_Ins_0_U1 ( .A(signal_1614), .B(ciphertext_s0[95]), .S(n349), 
        .Z(signal_591) );
  MUX2_X1 cell_274_Ins_1_U1 ( .A(signal_3622), .B(ciphertext_s1[95]), .S(n349), 
        .Z(signal_3849) );
  MUX2_X1 cell_277_Ins_0_U1 ( .A(signal_1613), .B(ciphertext_s0[40]), .S(n349), 
        .Z(signal_593) );
  MUX2_X1 cell_277_Ins_1_U1 ( .A(signal_2706), .B(ciphertext_s1[40]), .S(n349), 
        .Z(signal_3850) );
  MUX2_X1 cell_280_Ins_0_U1 ( .A(signal_1612), .B(ciphertext_s0[41]), .S(n342), 
        .Z(signal_595) );
  MUX2_X1 cell_280_Ins_1_U1 ( .A(signal_2709), .B(ciphertext_s1[41]), .S(n342), 
        .Z(signal_3851) );
  MUX2_X1 cell_283_Ins_0_U1 ( .A(signal_1611), .B(ciphertext_s0[42]), .S(n342), 
        .Z(signal_597) );
  MUX2_X1 cell_283_Ins_1_U1 ( .A(signal_2712), .B(ciphertext_s1[42]), .S(n342), 
        .Z(signal_3852) );
  MUX2_X1 cell_286_Ins_0_U1 ( .A(signal_1610), .B(ciphertext_s0[43]), .S(n342), 
        .Z(signal_599) );
  MUX2_X1 cell_286_Ins_1_U1 ( .A(signal_2715), .B(ciphertext_s1[43]), .S(n342), 
        .Z(signal_3853) );
  MUX2_X1 cell_289_Ins_0_U1 ( .A(signal_1609), .B(ciphertext_s0[44]), .S(n341), 
        .Z(signal_601) );
  MUX2_X1 cell_289_Ins_1_U1 ( .A(signal_2718), .B(ciphertext_s1[44]), .S(n341), 
        .Z(signal_3854) );
  MUX2_X1 cell_292_Ins_0_U1 ( .A(signal_1608), .B(ciphertext_s0[45]), .S(n341), 
        .Z(signal_603) );
  MUX2_X1 cell_292_Ins_1_U1 ( .A(signal_2721), .B(ciphertext_s1[45]), .S(n341), 
        .Z(signal_3855) );
  MUX2_X1 cell_295_Ins_0_U1 ( .A(signal_1607), .B(ciphertext_s0[46]), .S(n341), 
        .Z(signal_605) );
  MUX2_X1 cell_295_Ins_1_U1 ( .A(signal_2724), .B(ciphertext_s1[46]), .S(n341), 
        .Z(signal_3856) );
  MUX2_X1 cell_298_Ins_0_U1 ( .A(signal_1606), .B(ciphertext_s0[47]), .S(n348), 
        .Z(signal_607) );
  MUX2_X1 cell_298_Ins_1_U1 ( .A(signal_2727), .B(ciphertext_s1[47]), .S(n348), 
        .Z(signal_3857) );
  MUX2_X1 cell_301_Ins_0_U1 ( .A(signal_1605), .B(ciphertext_s0[32]), .S(n348), 
        .Z(signal_609) );
  MUX2_X1 cell_301_Ins_1_U1 ( .A(signal_2730), .B(ciphertext_s1[32]), .S(n348), 
        .Z(signal_3858) );
  MUX2_X1 cell_304_Ins_0_U1 ( .A(signal_1604), .B(ciphertext_s0[33]), .S(n348), 
        .Z(signal_611) );
  MUX2_X1 cell_304_Ins_1_U1 ( .A(signal_2733), .B(ciphertext_s1[33]), .S(n348), 
        .Z(signal_3859) );
  MUX2_X1 cell_307_Ins_0_U1 ( .A(signal_1603), .B(ciphertext_s0[34]), .S(n338), 
        .Z(signal_613) );
  MUX2_X1 cell_307_Ins_1_U1 ( .A(signal_2736), .B(ciphertext_s1[34]), .S(n338), 
        .Z(signal_3860) );
  MUX2_X1 cell_310_Ins_0_U1 ( .A(signal_1602), .B(ciphertext_s0[35]), .S(n348), 
        .Z(signal_615) );
  MUX2_X1 cell_310_Ins_1_U1 ( .A(signal_2739), .B(ciphertext_s1[35]), .S(n348), 
        .Z(signal_3861) );
  MUX2_X1 cell_313_Ins_0_U1 ( .A(signal_1601), .B(ciphertext_s0[36]), .S(n345), 
        .Z(signal_617) );
  MUX2_X1 cell_313_Ins_1_U1 ( .A(signal_2742), .B(ciphertext_s1[36]), .S(n345), 
        .Z(signal_3862) );
  MUX2_X1 cell_316_Ins_0_U1 ( .A(signal_1600), .B(ciphertext_s0[37]), .S(n347), 
        .Z(signal_619) );
  MUX2_X1 cell_316_Ins_1_U1 ( .A(signal_2745), .B(ciphertext_s1[37]), .S(n347), 
        .Z(signal_3863) );
  MUX2_X1 cell_319_Ins_0_U1 ( .A(signal_1599), .B(ciphertext_s0[38]), .S(n347), 
        .Z(signal_621) );
  MUX2_X1 cell_319_Ins_1_U1 ( .A(signal_2748), .B(ciphertext_s1[38]), .S(n347), 
        .Z(signal_3864) );
  MUX2_X1 cell_322_Ins_0_U1 ( .A(signal_1598), .B(ciphertext_s0[39]), .S(n347), 
        .Z(signal_623) );
  MUX2_X1 cell_322_Ins_1_U1 ( .A(signal_2751), .B(ciphertext_s1[39]), .S(n347), 
        .Z(signal_3865) );
  MUX2_X1 cell_325_Ins_0_U1 ( .A(signal_1597), .B(ciphertext_s0[56]), .S(n350), 
        .Z(signal_625) );
  MUX2_X1 cell_325_Ins_1_U1 ( .A(signal_2754), .B(ciphertext_s1[56]), .S(n350), 
        .Z(signal_3866) );
  MUX2_X1 cell_328_Ins_0_U1 ( .A(signal_1596), .B(ciphertext_s0[57]), .S(n349), 
        .Z(signal_627) );
  MUX2_X1 cell_328_Ins_1_U1 ( .A(signal_2757), .B(ciphertext_s1[57]), .S(n349), 
        .Z(signal_3867) );
  MUX2_X1 cell_331_Ins_0_U1 ( .A(signal_1595), .B(ciphertext_s0[58]), .S(n338), 
        .Z(signal_629) );
  MUX2_X1 cell_331_Ins_1_U1 ( .A(signal_2760), .B(ciphertext_s1[58]), .S(n338), 
        .Z(signal_3868) );
  MUX2_X1 cell_334_Ins_0_U1 ( .A(signal_1594), .B(ciphertext_s0[59]), .S(n346), 
        .Z(signal_631) );
  MUX2_X1 cell_334_Ins_1_U1 ( .A(signal_2763), .B(ciphertext_s1[59]), .S(n346), 
        .Z(signal_3869) );
  MUX2_X1 cell_337_Ins_0_U1 ( .A(signal_1593), .B(ciphertext_s0[60]), .S(n346), 
        .Z(signal_633) );
  MUX2_X1 cell_337_Ins_1_U1 ( .A(signal_2766), .B(ciphertext_s1[60]), .S(n346), 
        .Z(signal_3870) );
  MUX2_X1 cell_340_Ins_0_U1 ( .A(signal_1592), .B(ciphertext_s0[61]), .S(n346), 
        .Z(signal_635) );
  MUX2_X1 cell_340_Ins_1_U1 ( .A(signal_2769), .B(ciphertext_s1[61]), .S(n346), 
        .Z(signal_3871) );
  MUX2_X1 cell_343_Ins_0_U1 ( .A(signal_1591), .B(ciphertext_s0[62]), .S(n345), 
        .Z(signal_637) );
  MUX2_X1 cell_343_Ins_1_U1 ( .A(signal_2772), .B(ciphertext_s1[62]), .S(n345), 
        .Z(signal_3872) );
  MUX2_X1 cell_346_Ins_0_U1 ( .A(signal_1590), .B(ciphertext_s0[63]), .S(n345), 
        .Z(signal_639) );
  MUX2_X1 cell_346_Ins_1_U1 ( .A(signal_2775), .B(ciphertext_s1[63]), .S(n345), 
        .Z(signal_3873) );
  MUX2_X1 cell_349_Ins_0_U1 ( .A(signal_1589), .B(ciphertext_s0[48]), .S(n345), 
        .Z(signal_641) );
  MUX2_X1 cell_349_Ins_1_U1 ( .A(signal_3624), .B(ciphertext_s1[48]), .S(n345), 
        .Z(signal_3874) );
  MUX2_X1 cell_352_Ins_0_U1 ( .A(signal_1588), .B(ciphertext_s0[49]), .S(n344), 
        .Z(signal_643) );
  MUX2_X1 cell_352_Ins_1_U1 ( .A(signal_3626), .B(ciphertext_s1[49]), .S(n344), 
        .Z(signal_3875) );
  MUX2_X1 cell_355_Ins_0_U1 ( .A(signal_1587), .B(ciphertext_s0[50]), .S(n344), 
        .Z(signal_645) );
  MUX2_X1 cell_355_Ins_1_U1 ( .A(signal_3628), .B(ciphertext_s1[50]), .S(n344), 
        .Z(signal_3876) );
  MUX2_X1 cell_358_Ins_0_U1 ( .A(signal_1586), .B(ciphertext_s0[51]), .S(n344), 
        .Z(signal_647) );
  MUX2_X1 cell_358_Ins_1_U1 ( .A(signal_3630), .B(ciphertext_s1[51]), .S(n344), 
        .Z(signal_3877) );
  MUX2_X1 cell_361_Ins_0_U1 ( .A(signal_1585), .B(ciphertext_s0[52]), .S(n343), 
        .Z(signal_649) );
  MUX2_X1 cell_361_Ins_1_U1 ( .A(signal_3632), .B(ciphertext_s1[52]), .S(n343), 
        .Z(signal_3878) );
  MUX2_X1 cell_364_Ins_0_U1 ( .A(signal_1584), .B(ciphertext_s0[53]), .S(n343), 
        .Z(signal_651) );
  MUX2_X1 cell_364_Ins_1_U1 ( .A(signal_3634), .B(ciphertext_s1[53]), .S(n343), 
        .Z(signal_3879) );
  MUX2_X1 cell_367_Ins_0_U1 ( .A(signal_1583), .B(ciphertext_s0[54]), .S(n343), 
        .Z(signal_653) );
  MUX2_X1 cell_367_Ins_1_U1 ( .A(signal_3636), .B(ciphertext_s1[54]), .S(n343), 
        .Z(signal_3880) );
  MUX2_X1 cell_370_Ins_0_U1 ( .A(signal_1582), .B(ciphertext_s0[55]), .S(n342), 
        .Z(signal_655) );
  MUX2_X1 cell_370_Ins_1_U1 ( .A(signal_3638), .B(ciphertext_s1[55]), .S(n342), 
        .Z(signal_3881) );
  MUX2_X1 cell_373_Ins_0_U1 ( .A(signal_1581), .B(ciphertext_s0[0]), .S(n338), 
        .Z(signal_657) );
  MUX2_X1 cell_373_Ins_1_U1 ( .A(signal_2778), .B(ciphertext_s1[0]), .S(n338), 
        .Z(signal_3882) );
  MUX2_X1 cell_376_Ins_0_U1 ( .A(signal_1580), .B(ciphertext_s0[1]), .S(n345), 
        .Z(signal_659) );
  MUX2_X1 cell_376_Ins_1_U1 ( .A(signal_2781), .B(ciphertext_s1[1]), .S(n345), 
        .Z(signal_3883) );
  MUX2_X1 cell_379_Ins_0_U1 ( .A(signal_1579), .B(ciphertext_s0[2]), .S(n349), 
        .Z(signal_661) );
  MUX2_X1 cell_379_Ins_1_U1 ( .A(signal_2784), .B(ciphertext_s1[2]), .S(n349), 
        .Z(signal_3884) );
  MUX2_X1 cell_382_Ins_0_U1 ( .A(signal_1578), .B(ciphertext_s0[3]), .S(n339), 
        .Z(signal_663) );
  MUX2_X1 cell_382_Ins_1_U1 ( .A(signal_2787), .B(ciphertext_s1[3]), .S(n339), 
        .Z(signal_3885) );
  MUX2_X1 cell_385_Ins_0_U1 ( .A(signal_1577), .B(ciphertext_s0[4]), .S(n350), 
        .Z(signal_665) );
  MUX2_X1 cell_385_Ins_1_U1 ( .A(signal_2790), .B(ciphertext_s1[4]), .S(n350), 
        .Z(signal_3886) );
  MUX2_X1 cell_388_Ins_0_U1 ( .A(signal_1576), .B(ciphertext_s0[5]), .S(n349), 
        .Z(signal_667) );
  MUX2_X1 cell_388_Ins_1_U1 ( .A(signal_2793), .B(ciphertext_s1[5]), .S(n349), 
        .Z(signal_3887) );
  MUX2_X1 cell_391_Ins_0_U1 ( .A(signal_1575), .B(ciphertext_s0[6]), .S(n342), 
        .Z(signal_669) );
  MUX2_X1 cell_391_Ins_1_U1 ( .A(signal_2796), .B(ciphertext_s1[6]), .S(n342), 
        .Z(signal_3888) );
  MUX2_X1 cell_394_Ins_0_U1 ( .A(signal_1574), .B(ciphertext_s0[7]), .S(n342), 
        .Z(signal_671) );
  MUX2_X1 cell_394_Ins_1_U1 ( .A(signal_2799), .B(ciphertext_s1[7]), .S(n342), 
        .Z(signal_3889) );
  MUX2_X1 cell_397_Ins_0_U1 ( .A(signal_1573), .B(ciphertext_s0[24]), .S(n342), 
        .Z(signal_673) );
  MUX2_X1 cell_397_Ins_1_U1 ( .A(signal_2802), .B(ciphertext_s1[24]), .S(n342), 
        .Z(signal_3890) );
  MUX2_X1 cell_400_Ins_0_U1 ( .A(signal_1572), .B(ciphertext_s0[25]), .S(n341), 
        .Z(signal_675) );
  MUX2_X1 cell_400_Ins_1_U1 ( .A(signal_2805), .B(ciphertext_s1[25]), .S(n341), 
        .Z(signal_3891) );
  MUX2_X1 cell_403_Ins_0_U1 ( .A(signal_1571), .B(ciphertext_s0[26]), .S(n341), 
        .Z(signal_677) );
  MUX2_X1 cell_403_Ins_1_U1 ( .A(signal_2808), .B(ciphertext_s1[26]), .S(n341), 
        .Z(signal_3892) );
  MUX2_X1 cell_406_Ins_0_U1 ( .A(signal_1570), .B(ciphertext_s0[27]), .S(n341), 
        .Z(signal_679) );
  MUX2_X1 cell_406_Ins_1_U1 ( .A(signal_2811), .B(ciphertext_s1[27]), .S(n341), 
        .Z(signal_3893) );
  MUX2_X1 cell_409_Ins_0_U1 ( .A(signal_1569), .B(ciphertext_s0[28]), .S(n340), 
        .Z(signal_681) );
  MUX2_X1 cell_409_Ins_1_U1 ( .A(signal_2814), .B(ciphertext_s1[28]), .S(n340), 
        .Z(signal_3894) );
  MUX2_X1 cell_412_Ins_0_U1 ( .A(signal_1568), .B(ciphertext_s0[29]), .S(n340), 
        .Z(signal_683) );
  MUX2_X1 cell_412_Ins_1_U1 ( .A(signal_2817), .B(ciphertext_s1[29]), .S(n340), 
        .Z(signal_3895) );
  MUX2_X1 cell_415_Ins_0_U1 ( .A(signal_1567), .B(ciphertext_s0[30]), .S(n340), 
        .Z(signal_685) );
  MUX2_X1 cell_415_Ins_1_U1 ( .A(signal_2820), .B(ciphertext_s1[30]), .S(n340), 
        .Z(signal_3896) );
  MUX2_X1 cell_418_Ins_0_U1 ( .A(signal_1566), .B(ciphertext_s0[31]), .S(n338), 
        .Z(signal_687) );
  MUX2_X1 cell_418_Ins_1_U1 ( .A(signal_2823), .B(ciphertext_s1[31]), .S(n338), 
        .Z(signal_3897) );
  MUX2_X1 cell_421_Ins_0_U1 ( .A(signal_1565), .B(ciphertext_s0[16]), .S(n345), 
        .Z(signal_689) );
  MUX2_X1 cell_421_Ins_1_U1 ( .A(signal_2826), .B(ciphertext_s1[16]), .S(n345), 
        .Z(signal_3898) );
  MUX2_X1 cell_424_Ins_0_U1 ( .A(signal_1564), .B(ciphertext_s0[17]), .S(n342), 
        .Z(signal_691) );
  MUX2_X1 cell_424_Ins_1_U1 ( .A(signal_2829), .B(ciphertext_s1[17]), .S(n342), 
        .Z(signal_3899) );
  MUX2_X1 cell_427_Ins_0_U1 ( .A(signal_1563), .B(ciphertext_s0[18]), .S(n340), 
        .Z(signal_693) );
  MUX2_X1 cell_427_Ins_1_U1 ( .A(signal_2832), .B(ciphertext_s1[18]), .S(n340), 
        .Z(signal_3900) );
  MUX2_X1 cell_430_Ins_0_U1 ( .A(signal_1562), .B(ciphertext_s0[19]), .S(n344), 
        .Z(signal_695) );
  MUX2_X1 cell_430_Ins_1_U1 ( .A(signal_2835), .B(ciphertext_s1[19]), .S(n344), 
        .Z(signal_3901) );
  MUX2_X1 cell_433_Ins_0_U1 ( .A(signal_1561), .B(ciphertext_s0[20]), .S(n29), 
        .Z(signal_697) );
  MUX2_X1 cell_433_Ins_1_U1 ( .A(signal_2838), .B(ciphertext_s1[20]), .S(n29), 
        .Z(signal_3902) );
  MUX2_X1 cell_436_Ins_0_U1 ( .A(signal_1560), .B(ciphertext_s0[21]), .S(n350), 
        .Z(signal_699) );
  MUX2_X1 cell_436_Ins_1_U1 ( .A(signal_2841), .B(ciphertext_s1[21]), .S(n350), 
        .Z(signal_3903) );
  MUX2_X1 cell_439_Ins_0_U1 ( .A(signal_1559), .B(ciphertext_s0[22]), .S(n345), 
        .Z(signal_701) );
  MUX2_X1 cell_439_Ins_1_U1 ( .A(signal_2844), .B(ciphertext_s1[22]), .S(n345), 
        .Z(signal_3904) );
  MUX2_X1 cell_442_Ins_0_U1 ( .A(signal_1558), .B(ciphertext_s0[23]), .S(n350), 
        .Z(signal_703) );
  MUX2_X1 cell_442_Ins_1_U1 ( .A(signal_2847), .B(ciphertext_s1[23]), .S(n350), 
        .Z(signal_3905) );
  MUX2_X1 cell_469_Ins_0_U1 ( .A(plaintext_s0[120]), .B(ciphertext_s0[112]), 
        .S(n280), .Z(signal_1677) );
  MUX2_X1 cell_469_Ins_1_U1 ( .A(plaintext_s1[120]), .B(ciphertext_s1[112]), 
        .S(n280), .Z(signal_2562) );
  MUX2_X1 cell_470_Ins_0_U1 ( .A(plaintext_s0[121]), .B(ciphertext_s0[113]), 
        .S(n302), .Z(signal_1676) );
  MUX2_X1 cell_470_Ins_1_U1 ( .A(plaintext_s1[121]), .B(ciphertext_s1[113]), 
        .S(n302), .Z(signal_2565) );
  MUX2_X1 cell_471_Ins_0_U1 ( .A(plaintext_s0[122]), .B(ciphertext_s0[114]), 
        .S(n295), .Z(signal_1675) );
  MUX2_X1 cell_471_Ins_1_U1 ( .A(plaintext_s1[122]), .B(ciphertext_s1[114]), 
        .S(n295), .Z(signal_2568) );
  MUX2_X1 cell_472_Ins_0_U1 ( .A(plaintext_s0[123]), .B(ciphertext_s0[115]), 
        .S(n295), .Z(signal_1674) );
  MUX2_X1 cell_472_Ins_1_U1 ( .A(plaintext_s1[123]), .B(ciphertext_s1[115]), 
        .S(n295), .Z(signal_2571) );
  MUX2_X1 cell_473_Ins_0_U1 ( .A(plaintext_s0[124]), .B(ciphertext_s0[116]), 
        .S(n295), .Z(signal_1673) );
  MUX2_X1 cell_473_Ins_1_U1 ( .A(plaintext_s1[124]), .B(ciphertext_s1[116]), 
        .S(n295), .Z(signal_2574) );
  MUX2_X1 cell_474_Ins_0_U1 ( .A(plaintext_s0[125]), .B(ciphertext_s0[117]), 
        .S(n295), .Z(signal_1672) );
  MUX2_X1 cell_474_Ins_1_U1 ( .A(plaintext_s1[125]), .B(ciphertext_s1[117]), 
        .S(n295), .Z(signal_2577) );
  MUX2_X1 cell_475_Ins_0_U1 ( .A(plaintext_s0[126]), .B(ciphertext_s0[118]), 
        .S(n295), .Z(signal_1671) );
  MUX2_X1 cell_475_Ins_1_U1 ( .A(plaintext_s1[126]), .B(ciphertext_s1[118]), 
        .S(n295), .Z(signal_2580) );
  MUX2_X1 cell_476_Ins_0_U1 ( .A(plaintext_s0[127]), .B(ciphertext_s0[119]), 
        .S(n295), .Z(signal_1670) );
  MUX2_X1 cell_476_Ins_1_U1 ( .A(plaintext_s1[127]), .B(ciphertext_s1[119]), 
        .S(n295), .Z(signal_2583) );
  MUX2_X1 cell_477_Ins_0_U1 ( .A(plaintext_s0[112]), .B(ciphertext_s0[104]), 
        .S(n295), .Z(signal_1669) );
  MUX2_X1 cell_477_Ins_1_U1 ( .A(plaintext_s1[112]), .B(ciphertext_s1[104]), 
        .S(n295), .Z(signal_2586) );
  MUX2_X1 cell_478_Ins_0_U1 ( .A(plaintext_s0[113]), .B(ciphertext_s0[105]), 
        .S(n296), .Z(signal_1668) );
  MUX2_X1 cell_478_Ins_1_U1 ( .A(plaintext_s1[113]), .B(ciphertext_s1[105]), 
        .S(n296), .Z(signal_2589) );
  MUX2_X1 cell_479_Ins_0_U1 ( .A(plaintext_s0[114]), .B(ciphertext_s0[106]), 
        .S(n296), .Z(signal_1667) );
  MUX2_X1 cell_479_Ins_1_U1 ( .A(plaintext_s1[114]), .B(ciphertext_s1[106]), 
        .S(n296), .Z(signal_2592) );
  MUX2_X1 cell_480_Ins_0_U1 ( .A(plaintext_s0[115]), .B(ciphertext_s0[107]), 
        .S(n296), .Z(signal_1666) );
  MUX2_X1 cell_480_Ins_1_U1 ( .A(plaintext_s1[115]), .B(ciphertext_s1[107]), 
        .S(n296), .Z(signal_2595) );
  MUX2_X1 cell_481_Ins_0_U1 ( .A(plaintext_s0[116]), .B(ciphertext_s0[108]), 
        .S(n296), .Z(signal_1665) );
  MUX2_X1 cell_481_Ins_1_U1 ( .A(plaintext_s1[116]), .B(ciphertext_s1[108]), 
        .S(n296), .Z(signal_2598) );
  MUX2_X1 cell_482_Ins_0_U1 ( .A(plaintext_s0[117]), .B(ciphertext_s0[109]), 
        .S(n296), .Z(signal_1664) );
  MUX2_X1 cell_482_Ins_1_U1 ( .A(plaintext_s1[117]), .B(ciphertext_s1[109]), 
        .S(n296), .Z(signal_2601) );
  MUX2_X1 cell_483_Ins_0_U1 ( .A(plaintext_s0[118]), .B(ciphertext_s0[110]), 
        .S(n296), .Z(signal_1663) );
  MUX2_X1 cell_483_Ins_1_U1 ( .A(plaintext_s1[118]), .B(ciphertext_s1[110]), 
        .S(n296), .Z(signal_2604) );
  MUX2_X1 cell_484_Ins_0_U1 ( .A(plaintext_s0[119]), .B(ciphertext_s0[111]), 
        .S(n296), .Z(signal_1662) );
  MUX2_X1 cell_484_Ins_1_U1 ( .A(plaintext_s1[119]), .B(ciphertext_s1[111]), 
        .S(n296), .Z(signal_2607) );
  MUX2_X1 cell_485_Ins_0_U1 ( .A(plaintext_s0[104]), .B(ciphertext_s0[96]), 
        .S(n297), .Z(signal_1661) );
  MUX2_X1 cell_485_Ins_1_U1 ( .A(plaintext_s1[104]), .B(ciphertext_s1[96]), 
        .S(n297), .Z(signal_2610) );
  MUX2_X1 cell_486_Ins_0_U1 ( .A(plaintext_s0[105]), .B(ciphertext_s0[97]), 
        .S(n297), .Z(signal_1660) );
  MUX2_X1 cell_486_Ins_1_U1 ( .A(plaintext_s1[105]), .B(ciphertext_s1[97]), 
        .S(n297), .Z(signal_2613) );
  MUX2_X1 cell_487_Ins_0_U1 ( .A(plaintext_s0[106]), .B(ciphertext_s0[98]), 
        .S(n297), .Z(signal_1659) );
  MUX2_X1 cell_487_Ins_1_U1 ( .A(plaintext_s1[106]), .B(ciphertext_s1[98]), 
        .S(n297), .Z(signal_2616) );
  MUX2_X1 cell_488_Ins_0_U1 ( .A(plaintext_s0[107]), .B(ciphertext_s0[99]), 
        .S(n297), .Z(signal_1658) );
  MUX2_X1 cell_488_Ins_1_U1 ( .A(plaintext_s1[107]), .B(ciphertext_s1[99]), 
        .S(n297), .Z(signal_2619) );
  MUX2_X1 cell_489_Ins_0_U1 ( .A(plaintext_s0[108]), .B(ciphertext_s0[100]), 
        .S(n297), .Z(signal_1657) );
  MUX2_X1 cell_489_Ins_1_U1 ( .A(plaintext_s1[108]), .B(ciphertext_s1[100]), 
        .S(n297), .Z(signal_2622) );
  MUX2_X1 cell_490_Ins_0_U1 ( .A(plaintext_s0[109]), .B(ciphertext_s0[101]), 
        .S(n297), .Z(signal_1656) );
  MUX2_X1 cell_490_Ins_1_U1 ( .A(plaintext_s1[109]), .B(ciphertext_s1[101]), 
        .S(n297), .Z(signal_2625) );
  MUX2_X1 cell_491_Ins_0_U1 ( .A(plaintext_s0[110]), .B(ciphertext_s0[102]), 
        .S(n297), .Z(signal_1655) );
  MUX2_X1 cell_491_Ins_1_U1 ( .A(plaintext_s1[110]), .B(ciphertext_s1[102]), 
        .S(n297), .Z(signal_2628) );
  MUX2_X1 cell_492_Ins_0_U1 ( .A(plaintext_s0[111]), .B(ciphertext_s0[103]), 
        .S(n298), .Z(signal_1654) );
  MUX2_X1 cell_492_Ins_1_U1 ( .A(plaintext_s1[111]), .B(ciphertext_s1[103]), 
        .S(n298), .Z(signal_2631) );
  MUX2_X1 cell_493_Ins_0_U1 ( .A(ciphertext_s0[88]), .B(signal_1429), .S(n312), 
        .Z(signal_1549) );
  MUX2_X1 cell_493_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(signal_3282), .S(n312), 
        .Z(signal_3434) );
  MUX2_X1 cell_494_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(signal_1428), .S(n308), 
        .Z(signal_1548) );
  MUX2_X1 cell_494_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(signal_3283), .S(n308), 
        .Z(signal_3435) );
  MUX2_X1 cell_495_Ins_0_U1 ( .A(ciphertext_s0[90]), .B(signal_1427), .S(n320), 
        .Z(signal_1547) );
  MUX2_X1 cell_495_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(signal_3284), .S(n320), 
        .Z(signal_3436) );
  MUX2_X1 cell_496_Ins_0_U1 ( .A(ciphertext_s0[91]), .B(signal_1426), .S(n323), 
        .Z(signal_1546) );
  MUX2_X1 cell_496_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(signal_3285), .S(n323), 
        .Z(signal_3437) );
  MUX2_X1 cell_497_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(signal_1425), .S(n313), 
        .Z(signal_1545) );
  MUX2_X1 cell_497_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(signal_3286), .S(n313), 
        .Z(signal_3438) );
  MUX2_X1 cell_498_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(signal_1424), .S(n323), 
        .Z(signal_1544) );
  MUX2_X1 cell_498_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(signal_3287), .S(n323), 
        .Z(signal_3439) );
  MUX2_X1 cell_499_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(signal_1423), .S(n322), 
        .Z(signal_1543) );
  MUX2_X1 cell_499_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(signal_3288), .S(n322), 
        .Z(signal_3440) );
  MUX2_X1 cell_500_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(signal_1422), .S(n307), 
        .Z(signal_1542) );
  MUX2_X1 cell_500_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(signal_3289), .S(n307), 
        .Z(signal_3441) );
  MUX2_X1 cell_501_Ins_0_U1 ( .A(plaintext_s0[96]), .B(signal_1549), .S(n298), 
        .Z(signal_1653) );
  MUX2_X1 cell_501_Ins_1_U1 ( .A(plaintext_s1[96]), .B(signal_3434), .S(n298), 
        .Z(signal_3592) );
  MUX2_X1 cell_502_Ins_0_U1 ( .A(plaintext_s0[97]), .B(signal_1548), .S(n298), 
        .Z(signal_1652) );
  MUX2_X1 cell_502_Ins_1_U1 ( .A(plaintext_s1[97]), .B(signal_3435), .S(n298), 
        .Z(signal_3594) );
  MUX2_X1 cell_503_Ins_0_U1 ( .A(plaintext_s0[98]), .B(signal_1547), .S(n298), 
        .Z(signal_1651) );
  MUX2_X1 cell_503_Ins_1_U1 ( .A(plaintext_s1[98]), .B(signal_3436), .S(n298), 
        .Z(signal_3596) );
  MUX2_X1 cell_504_Ins_0_U1 ( .A(plaintext_s0[99]), .B(signal_1546), .S(n298), 
        .Z(signal_1650) );
  MUX2_X1 cell_504_Ins_1_U1 ( .A(plaintext_s1[99]), .B(signal_3437), .S(n298), 
        .Z(signal_3598) );
  MUX2_X1 cell_505_Ins_0_U1 ( .A(plaintext_s0[100]), .B(signal_1545), .S(n298), 
        .Z(signal_1649) );
  MUX2_X1 cell_505_Ins_1_U1 ( .A(plaintext_s1[100]), .B(signal_3438), .S(n298), 
        .Z(signal_3600) );
  MUX2_X1 cell_506_Ins_0_U1 ( .A(plaintext_s0[101]), .B(signal_1544), .S(n298), 
        .Z(signal_1648) );
  MUX2_X1 cell_506_Ins_1_U1 ( .A(plaintext_s1[101]), .B(signal_3439), .S(n298), 
        .Z(signal_3602) );
  MUX2_X1 cell_507_Ins_0_U1 ( .A(plaintext_s0[102]), .B(signal_1543), .S(n299), 
        .Z(signal_1647) );
  MUX2_X1 cell_507_Ins_1_U1 ( .A(plaintext_s1[102]), .B(signal_3440), .S(n299), 
        .Z(signal_3604) );
  MUX2_X1 cell_508_Ins_0_U1 ( .A(plaintext_s0[103]), .B(signal_1542), .S(n299), 
        .Z(signal_1646) );
  MUX2_X1 cell_508_Ins_1_U1 ( .A(plaintext_s1[103]), .B(signal_3441), .S(n299), 
        .Z(signal_3606) );
  MUX2_X1 cell_509_Ins_0_U1 ( .A(plaintext_s0[88]), .B(ciphertext_s0[80]), .S(
        n299), .Z(signal_1645) );
  MUX2_X1 cell_509_Ins_1_U1 ( .A(plaintext_s1[88]), .B(ciphertext_s1[80]), .S(
        n299), .Z(signal_2634) );
  MUX2_X1 cell_510_Ins_0_U1 ( .A(plaintext_s0[89]), .B(ciphertext_s0[81]), .S(
        n299), .Z(signal_1644) );
  MUX2_X1 cell_510_Ins_1_U1 ( .A(plaintext_s1[89]), .B(ciphertext_s1[81]), .S(
        n299), .Z(signal_2637) );
  MUX2_X1 cell_511_Ins_0_U1 ( .A(plaintext_s0[90]), .B(ciphertext_s0[82]), .S(
        n299), .Z(signal_1643) );
  MUX2_X1 cell_511_Ins_1_U1 ( .A(plaintext_s1[90]), .B(ciphertext_s1[82]), .S(
        n299), .Z(signal_2640) );
  MUX2_X1 cell_512_Ins_0_U1 ( .A(plaintext_s0[91]), .B(ciphertext_s0[83]), .S(
        n299), .Z(signal_1642) );
  MUX2_X1 cell_512_Ins_1_U1 ( .A(plaintext_s1[91]), .B(ciphertext_s1[83]), .S(
        n299), .Z(signal_2643) );
  MUX2_X1 cell_513_Ins_0_U1 ( .A(plaintext_s0[92]), .B(ciphertext_s0[84]), .S(
        n299), .Z(signal_1641) );
  MUX2_X1 cell_513_Ins_1_U1 ( .A(plaintext_s1[92]), .B(ciphertext_s1[84]), .S(
        n299), .Z(signal_2646) );
  MUX2_X1 cell_514_Ins_0_U1 ( .A(plaintext_s0[93]), .B(ciphertext_s0[85]), .S(
        n288), .Z(signal_1640) );
  MUX2_X1 cell_514_Ins_1_U1 ( .A(plaintext_s1[93]), .B(ciphertext_s1[85]), .S(
        n288), .Z(signal_2649) );
  MUX2_X1 cell_515_Ins_0_U1 ( .A(plaintext_s0[94]), .B(ciphertext_s0[86]), .S(
        n293), .Z(signal_1639) );
  MUX2_X1 cell_515_Ins_1_U1 ( .A(plaintext_s1[94]), .B(ciphertext_s1[86]), .S(
        n293), .Z(signal_2652) );
  MUX2_X1 cell_516_Ins_0_U1 ( .A(plaintext_s0[95]), .B(ciphertext_s0[87]), .S(
        n291), .Z(signal_1638) );
  MUX2_X1 cell_516_Ins_1_U1 ( .A(plaintext_s1[95]), .B(ciphertext_s1[87]), .S(
        n291), .Z(signal_2655) );
  MUX2_X1 cell_517_Ins_0_U1 ( .A(plaintext_s0[80]), .B(ciphertext_s0[72]), .S(
        n288), .Z(signal_1637) );
  MUX2_X1 cell_517_Ins_1_U1 ( .A(plaintext_s1[80]), .B(ciphertext_s1[72]), .S(
        n288), .Z(signal_2658) );
  MUX2_X1 cell_518_Ins_0_U1 ( .A(plaintext_s0[81]), .B(ciphertext_s0[73]), .S(
        n293), .Z(signal_1636) );
  MUX2_X1 cell_518_Ins_1_U1 ( .A(plaintext_s1[81]), .B(ciphertext_s1[73]), .S(
        n293), .Z(signal_2661) );
  MUX2_X1 cell_519_Ins_0_U1 ( .A(plaintext_s0[82]), .B(ciphertext_s0[74]), .S(
        n291), .Z(signal_1635) );
  MUX2_X1 cell_519_Ins_1_U1 ( .A(plaintext_s1[82]), .B(ciphertext_s1[74]), .S(
        n291), .Z(signal_2664) );
  MUX2_X1 cell_520_Ins_0_U1 ( .A(plaintext_s0[83]), .B(ciphertext_s0[75]), .S(
        n282), .Z(signal_1634) );
  MUX2_X1 cell_520_Ins_1_U1 ( .A(plaintext_s1[83]), .B(ciphertext_s1[75]), .S(
        n282), .Z(signal_2667) );
  MUX2_X1 cell_521_Ins_0_U1 ( .A(plaintext_s0[84]), .B(ciphertext_s0[76]), .S(
        n300), .Z(signal_1633) );
  MUX2_X1 cell_521_Ins_1_U1 ( .A(plaintext_s1[84]), .B(ciphertext_s1[76]), .S(
        n300), .Z(signal_2670) );
  MUX2_X1 cell_522_Ins_0_U1 ( .A(plaintext_s0[85]), .B(ciphertext_s0[77]), .S(
        n300), .Z(signal_1632) );
  MUX2_X1 cell_522_Ins_1_U1 ( .A(plaintext_s1[85]), .B(ciphertext_s1[77]), .S(
        n300), .Z(signal_2673) );
  MUX2_X1 cell_523_Ins_0_U1 ( .A(plaintext_s0[86]), .B(ciphertext_s0[78]), .S(
        n300), .Z(signal_1631) );
  MUX2_X1 cell_523_Ins_1_U1 ( .A(plaintext_s1[86]), .B(ciphertext_s1[78]), .S(
        n300), .Z(signal_2676) );
  MUX2_X1 cell_524_Ins_0_U1 ( .A(plaintext_s0[87]), .B(ciphertext_s0[79]), .S(
        n300), .Z(signal_1630) );
  MUX2_X1 cell_524_Ins_1_U1 ( .A(plaintext_s1[87]), .B(ciphertext_s1[79]), .S(
        n300), .Z(signal_2679) );
  MUX2_X1 cell_525_Ins_0_U1 ( .A(plaintext_s0[72]), .B(ciphertext_s0[64]), .S(
        n300), .Z(signal_1629) );
  MUX2_X1 cell_525_Ins_1_U1 ( .A(plaintext_s1[72]), .B(ciphertext_s1[64]), .S(
        n300), .Z(signal_2682) );
  MUX2_X1 cell_526_Ins_0_U1 ( .A(plaintext_s0[73]), .B(ciphertext_s0[65]), .S(
        n300), .Z(signal_1628) );
  MUX2_X1 cell_526_Ins_1_U1 ( .A(plaintext_s1[73]), .B(ciphertext_s1[65]), .S(
        n300), .Z(signal_2685) );
  MUX2_X1 cell_527_Ins_0_U1 ( .A(plaintext_s0[74]), .B(ciphertext_s0[66]), .S(
        n300), .Z(signal_1627) );
  MUX2_X1 cell_527_Ins_1_U1 ( .A(plaintext_s1[74]), .B(ciphertext_s1[66]), .S(
        n300), .Z(signal_2688) );
  MUX2_X1 cell_528_Ins_0_U1 ( .A(plaintext_s0[75]), .B(ciphertext_s0[67]), .S(
        n301), .Z(signal_1626) );
  MUX2_X1 cell_528_Ins_1_U1 ( .A(plaintext_s1[75]), .B(ciphertext_s1[67]), .S(
        n301), .Z(signal_2691) );
  MUX2_X1 cell_529_Ins_0_U1 ( .A(plaintext_s0[76]), .B(ciphertext_s0[68]), .S(
        n301), .Z(signal_1625) );
  MUX2_X1 cell_529_Ins_1_U1 ( .A(plaintext_s1[76]), .B(ciphertext_s1[68]), .S(
        n301), .Z(signal_2694) );
  MUX2_X1 cell_530_Ins_0_U1 ( .A(plaintext_s0[77]), .B(ciphertext_s0[69]), .S(
        n301), .Z(signal_1624) );
  MUX2_X1 cell_530_Ins_1_U1 ( .A(plaintext_s1[77]), .B(ciphertext_s1[69]), .S(
        n301), .Z(signal_2697) );
  MUX2_X1 cell_531_Ins_0_U1 ( .A(plaintext_s0[78]), .B(ciphertext_s0[70]), .S(
        n301), .Z(signal_1623) );
  MUX2_X1 cell_531_Ins_1_U1 ( .A(plaintext_s1[78]), .B(ciphertext_s1[70]), .S(
        n301), .Z(signal_2700) );
  MUX2_X1 cell_532_Ins_0_U1 ( .A(plaintext_s0[79]), .B(ciphertext_s0[71]), .S(
        n301), .Z(signal_1622) );
  MUX2_X1 cell_532_Ins_1_U1 ( .A(plaintext_s1[79]), .B(ciphertext_s1[71]), .S(
        n301), .Z(signal_2703) );
  MUX2_X1 cell_533_Ins_0_U1 ( .A(ciphertext_s0[56]), .B(signal_1437), .S(n307), 
        .Z(signal_1541) );
  MUX2_X1 cell_533_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(signal_3274), .S(n307), 
        .Z(signal_3442) );
  MUX2_X1 cell_534_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(signal_1436), .S(n307), 
        .Z(signal_1540) );
  MUX2_X1 cell_534_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(signal_3275), .S(n307), 
        .Z(signal_3443) );
  MUX2_X1 cell_535_Ins_0_U1 ( .A(ciphertext_s0[58]), .B(signal_1435), .S(n307), 
        .Z(signal_1539) );
  MUX2_X1 cell_535_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(signal_3276), .S(n307), 
        .Z(signal_3444) );
  MUX2_X1 cell_536_Ins_0_U1 ( .A(ciphertext_s0[59]), .B(signal_1434), .S(n307), 
        .Z(signal_1538) );
  MUX2_X1 cell_536_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(signal_3277), .S(n307), 
        .Z(signal_3445) );
  MUX2_X1 cell_537_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(signal_1433), .S(n307), 
        .Z(signal_1537) );
  MUX2_X1 cell_537_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(signal_3278), .S(n307), 
        .Z(signal_3446) );
  MUX2_X1 cell_538_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(signal_1432), .S(n307), 
        .Z(signal_1536) );
  MUX2_X1 cell_538_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(signal_3279), .S(n307), 
        .Z(signal_3447) );
  MUX2_X1 cell_539_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(signal_1431), .S(n308), 
        .Z(signal_1535) );
  MUX2_X1 cell_539_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(signal_3280), .S(n308), 
        .Z(signal_3448) );
  MUX2_X1 cell_540_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(signal_1430), .S(n308), 
        .Z(signal_1534) );
  MUX2_X1 cell_540_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(signal_3281), .S(n308), 
        .Z(signal_3449) );
  MUX2_X1 cell_541_Ins_0_U1 ( .A(plaintext_s0[64]), .B(signal_1541), .S(n301), 
        .Z(signal_1621) );
  MUX2_X1 cell_541_Ins_1_U1 ( .A(plaintext_s1[64]), .B(signal_3442), .S(n301), 
        .Z(signal_3608) );
  MUX2_X1 cell_542_Ins_0_U1 ( .A(plaintext_s0[65]), .B(signal_1540), .S(n301), 
        .Z(signal_1620) );
  MUX2_X1 cell_542_Ins_1_U1 ( .A(plaintext_s1[65]), .B(signal_3443), .S(n301), 
        .Z(signal_3610) );
  MUX2_X1 cell_543_Ins_0_U1 ( .A(plaintext_s0[66]), .B(signal_1539), .S(n302), 
        .Z(signal_1619) );
  MUX2_X1 cell_543_Ins_1_U1 ( .A(plaintext_s1[66]), .B(signal_3444), .S(n302), 
        .Z(signal_3612) );
  MUX2_X1 cell_544_Ins_0_U1 ( .A(plaintext_s0[67]), .B(signal_1538), .S(n302), 
        .Z(signal_1618) );
  MUX2_X1 cell_544_Ins_1_U1 ( .A(plaintext_s1[67]), .B(signal_3445), .S(n302), 
        .Z(signal_3614) );
  MUX2_X1 cell_545_Ins_0_U1 ( .A(plaintext_s0[68]), .B(signal_1537), .S(n302), 
        .Z(signal_1617) );
  MUX2_X1 cell_545_Ins_1_U1 ( .A(plaintext_s1[68]), .B(signal_3446), .S(n302), 
        .Z(signal_3616) );
  MUX2_X1 cell_546_Ins_0_U1 ( .A(plaintext_s0[69]), .B(signal_1536), .S(n302), 
        .Z(signal_1616) );
  MUX2_X1 cell_546_Ins_1_U1 ( .A(plaintext_s1[69]), .B(signal_3447), .S(n302), 
        .Z(signal_3618) );
  MUX2_X1 cell_547_Ins_0_U1 ( .A(plaintext_s0[70]), .B(signal_1535), .S(n302), 
        .Z(signal_1615) );
  MUX2_X1 cell_547_Ins_1_U1 ( .A(plaintext_s1[70]), .B(signal_3448), .S(n302), 
        .Z(signal_3620) );
  MUX2_X1 cell_548_Ins_0_U1 ( .A(plaintext_s0[71]), .B(signal_1534), .S(n302), 
        .Z(signal_1614) );
  MUX2_X1 cell_548_Ins_1_U1 ( .A(plaintext_s1[71]), .B(signal_3449), .S(n302), 
        .Z(signal_3622) );
  MUX2_X1 cell_549_Ins_0_U1 ( .A(plaintext_s0[56]), .B(ciphertext_s0[48]), .S(
        n303), .Z(signal_1613) );
  MUX2_X1 cell_549_Ins_1_U1 ( .A(plaintext_s1[56]), .B(ciphertext_s1[48]), .S(
        n303), .Z(signal_2706) );
  MUX2_X1 cell_550_Ins_0_U1 ( .A(plaintext_s0[57]), .B(ciphertext_s0[49]), .S(
        n303), .Z(signal_1612) );
  MUX2_X1 cell_550_Ins_1_U1 ( .A(plaintext_s1[57]), .B(ciphertext_s1[49]), .S(
        n303), .Z(signal_2709) );
  MUX2_X1 cell_551_Ins_0_U1 ( .A(plaintext_s0[58]), .B(ciphertext_s0[50]), .S(
        n303), .Z(signal_1611) );
  MUX2_X1 cell_551_Ins_1_U1 ( .A(plaintext_s1[58]), .B(ciphertext_s1[50]), .S(
        n303), .Z(signal_2712) );
  MUX2_X1 cell_552_Ins_0_U1 ( .A(plaintext_s0[59]), .B(ciphertext_s0[51]), .S(
        n303), .Z(signal_1610) );
  MUX2_X1 cell_552_Ins_1_U1 ( .A(plaintext_s1[59]), .B(ciphertext_s1[51]), .S(
        n303), .Z(signal_2715) );
  MUX2_X1 cell_553_Ins_0_U1 ( .A(plaintext_s0[60]), .B(ciphertext_s0[52]), .S(
        n303), .Z(signal_1609) );
  MUX2_X1 cell_553_Ins_1_U1 ( .A(plaintext_s1[60]), .B(ciphertext_s1[52]), .S(
        n303), .Z(signal_2718) );
  MUX2_X1 cell_554_Ins_0_U1 ( .A(plaintext_s0[61]), .B(ciphertext_s0[53]), .S(
        n303), .Z(signal_1608) );
  MUX2_X1 cell_554_Ins_1_U1 ( .A(plaintext_s1[61]), .B(ciphertext_s1[53]), .S(
        n303), .Z(signal_2721) );
  MUX2_X1 cell_555_Ins_0_U1 ( .A(plaintext_s0[62]), .B(ciphertext_s0[54]), .S(
        n303), .Z(signal_1607) );
  MUX2_X1 cell_555_Ins_1_U1 ( .A(plaintext_s1[62]), .B(ciphertext_s1[54]), .S(
        n303), .Z(signal_2724) );
  MUX2_X1 cell_556_Ins_0_U1 ( .A(plaintext_s0[63]), .B(ciphertext_s0[55]), .S(
        n304), .Z(signal_1606) );
  MUX2_X1 cell_556_Ins_1_U1 ( .A(plaintext_s1[63]), .B(ciphertext_s1[55]), .S(
        n304), .Z(signal_2727) );
  MUX2_X1 cell_557_Ins_0_U1 ( .A(plaintext_s0[48]), .B(ciphertext_s0[40]), .S(
        n304), .Z(signal_1605) );
  MUX2_X1 cell_557_Ins_1_U1 ( .A(plaintext_s1[48]), .B(ciphertext_s1[40]), .S(
        n304), .Z(signal_2730) );
  MUX2_X1 cell_558_Ins_0_U1 ( .A(plaintext_s0[49]), .B(ciphertext_s0[41]), .S(
        n304), .Z(signal_1604) );
  MUX2_X1 cell_558_Ins_1_U1 ( .A(plaintext_s1[49]), .B(ciphertext_s1[41]), .S(
        n304), .Z(signal_2733) );
  MUX2_X1 cell_559_Ins_0_U1 ( .A(plaintext_s0[50]), .B(ciphertext_s0[42]), .S(
        n304), .Z(signal_1603) );
  MUX2_X1 cell_559_Ins_1_U1 ( .A(plaintext_s1[50]), .B(ciphertext_s1[42]), .S(
        n304), .Z(signal_2736) );
  MUX2_X1 cell_560_Ins_0_U1 ( .A(plaintext_s0[51]), .B(ciphertext_s0[43]), .S(
        n304), .Z(signal_1602) );
  MUX2_X1 cell_560_Ins_1_U1 ( .A(plaintext_s1[51]), .B(ciphertext_s1[43]), .S(
        n304), .Z(signal_2739) );
  MUX2_X1 cell_561_Ins_0_U1 ( .A(plaintext_s0[52]), .B(ciphertext_s0[44]), .S(
        n304), .Z(signal_1601) );
  MUX2_X1 cell_561_Ins_1_U1 ( .A(plaintext_s1[52]), .B(ciphertext_s1[44]), .S(
        n304), .Z(signal_2742) );
  MUX2_X1 cell_562_Ins_0_U1 ( .A(plaintext_s0[53]), .B(ciphertext_s0[45]), .S(
        n305), .Z(signal_1600) );
  MUX2_X1 cell_562_Ins_1_U1 ( .A(plaintext_s1[53]), .B(ciphertext_s1[45]), .S(
        n305), .Z(signal_2745) );
  MUX2_X1 cell_563_Ins_0_U1 ( .A(plaintext_s0[54]), .B(ciphertext_s0[46]), .S(
        n304), .Z(signal_1599) );
  MUX2_X1 cell_563_Ins_1_U1 ( .A(plaintext_s1[54]), .B(ciphertext_s1[46]), .S(
        n304), .Z(signal_2748) );
  MUX2_X1 cell_564_Ins_0_U1 ( .A(plaintext_s0[55]), .B(ciphertext_s0[47]), .S(
        n305), .Z(signal_1598) );
  MUX2_X1 cell_564_Ins_1_U1 ( .A(plaintext_s1[55]), .B(ciphertext_s1[47]), .S(
        n305), .Z(signal_2751) );
  MUX2_X1 cell_565_Ins_0_U1 ( .A(plaintext_s0[40]), .B(ciphertext_s0[32]), .S(
        n305), .Z(signal_1597) );
  MUX2_X1 cell_565_Ins_1_U1 ( .A(plaintext_s1[40]), .B(ciphertext_s1[32]), .S(
        n305), .Z(signal_2754) );
  MUX2_X1 cell_566_Ins_0_U1 ( .A(plaintext_s0[41]), .B(ciphertext_s0[33]), .S(
        n305), .Z(signal_1596) );
  MUX2_X1 cell_566_Ins_1_U1 ( .A(plaintext_s1[41]), .B(ciphertext_s1[33]), .S(
        n305), .Z(signal_2757) );
  MUX2_X1 cell_567_Ins_0_U1 ( .A(plaintext_s0[42]), .B(ciphertext_s0[34]), .S(
        n305), .Z(signal_1595) );
  MUX2_X1 cell_567_Ins_1_U1 ( .A(plaintext_s1[42]), .B(ciphertext_s1[34]), .S(
        n305), .Z(signal_2760) );
  MUX2_X1 cell_568_Ins_0_U1 ( .A(plaintext_s0[43]), .B(ciphertext_s0[35]), .S(
        n305), .Z(signal_1594) );
  MUX2_X1 cell_568_Ins_1_U1 ( .A(plaintext_s1[43]), .B(ciphertext_s1[35]), .S(
        n305), .Z(signal_2763) );
  MUX2_X1 cell_569_Ins_0_U1 ( .A(plaintext_s0[44]), .B(ciphertext_s0[36]), .S(
        n305), .Z(signal_1593) );
  MUX2_X1 cell_569_Ins_1_U1 ( .A(plaintext_s1[44]), .B(ciphertext_s1[36]), .S(
        n305), .Z(signal_2766) );
  MUX2_X1 cell_570_Ins_0_U1 ( .A(plaintext_s0[45]), .B(ciphertext_s0[37]), .S(
        n306), .Z(signal_1592) );
  MUX2_X1 cell_570_Ins_1_U1 ( .A(plaintext_s1[45]), .B(ciphertext_s1[37]), .S(
        n306), .Z(signal_2769) );
  MUX2_X1 cell_571_Ins_0_U1 ( .A(plaintext_s0[46]), .B(ciphertext_s0[38]), .S(
        n306), .Z(signal_1591) );
  MUX2_X1 cell_571_Ins_1_U1 ( .A(plaintext_s1[46]), .B(ciphertext_s1[38]), .S(
        n306), .Z(signal_2772) );
  MUX2_X1 cell_572_Ins_0_U1 ( .A(plaintext_s0[47]), .B(ciphertext_s0[39]), .S(
        n306), .Z(signal_1590) );
  MUX2_X1 cell_572_Ins_1_U1 ( .A(plaintext_s1[47]), .B(ciphertext_s1[39]), .S(
        n306), .Z(signal_2775) );
  MUX2_X1 cell_573_Ins_0_U1 ( .A(ciphertext_s0[24]), .B(signal_1445), .S(n308), 
        .Z(signal_1533) );
  MUX2_X1 cell_573_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(signal_3266), .S(n308), 
        .Z(signal_3450) );
  MUX2_X1 cell_574_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(signal_1444), .S(n308), 
        .Z(signal_1532) );
  MUX2_X1 cell_574_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(signal_3267), .S(n308), 
        .Z(signal_3451) );
  MUX2_X1 cell_575_Ins_0_U1 ( .A(ciphertext_s0[26]), .B(signal_1443), .S(n308), 
        .Z(signal_1531) );
  MUX2_X1 cell_575_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(signal_3268), .S(n308), 
        .Z(signal_3452) );
  MUX2_X1 cell_576_Ins_0_U1 ( .A(ciphertext_s0[27]), .B(signal_1442), .S(n308), 
        .Z(signal_1530) );
  MUX2_X1 cell_576_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(signal_3269), .S(n308), 
        .Z(signal_3453) );
  MUX2_X1 cell_577_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(signal_1441), .S(n308), 
        .Z(signal_1529) );
  MUX2_X1 cell_577_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(signal_3270), .S(n308), 
        .Z(signal_3454) );
  MUX2_X1 cell_578_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(signal_1440), .S(n309), 
        .Z(signal_1528) );
  MUX2_X1 cell_578_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(signal_3271), .S(n309), 
        .Z(signal_3455) );
  MUX2_X1 cell_579_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(signal_1439), .S(n309), 
        .Z(signal_1527) );
  MUX2_X1 cell_579_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(signal_3272), .S(n309), 
        .Z(signal_3456) );
  MUX2_X1 cell_580_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(signal_1438), .S(n309), 
        .Z(signal_1526) );
  MUX2_X1 cell_580_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(signal_3273), .S(n309), 
        .Z(signal_3457) );
  MUX2_X1 cell_581_Ins_0_U1 ( .A(plaintext_s0[32]), .B(signal_1533), .S(n306), 
        .Z(signal_1589) );
  MUX2_X1 cell_581_Ins_1_U1 ( .A(plaintext_s1[32]), .B(signal_3450), .S(n306), 
        .Z(signal_3624) );
  MUX2_X1 cell_582_Ins_0_U1 ( .A(plaintext_s0[33]), .B(signal_1532), .S(n306), 
        .Z(signal_1588) );
  MUX2_X1 cell_582_Ins_1_U1 ( .A(plaintext_s1[33]), .B(signal_3451), .S(n306), 
        .Z(signal_3626) );
  MUX2_X1 cell_583_Ins_0_U1 ( .A(plaintext_s0[34]), .B(signal_1531), .S(n306), 
        .Z(signal_1587) );
  MUX2_X1 cell_583_Ins_1_U1 ( .A(plaintext_s1[34]), .B(signal_3452), .S(n306), 
        .Z(signal_3628) );
  MUX2_X1 cell_584_Ins_0_U1 ( .A(plaintext_s0[35]), .B(signal_1530), .S(n287), 
        .Z(signal_1586) );
  MUX2_X1 cell_584_Ins_1_U1 ( .A(plaintext_s1[35]), .B(signal_3453), .S(n287), 
        .Z(signal_3630) );
  MUX2_X1 cell_585_Ins_0_U1 ( .A(plaintext_s0[36]), .B(signal_1529), .S(n306), 
        .Z(signal_1585) );
  MUX2_X1 cell_585_Ins_1_U1 ( .A(plaintext_s1[36]), .B(signal_3454), .S(n306), 
        .Z(signal_3632) );
  MUX2_X1 cell_586_Ins_0_U1 ( .A(plaintext_s0[37]), .B(signal_1528), .S(n290), 
        .Z(signal_1584) );
  MUX2_X1 cell_586_Ins_1_U1 ( .A(plaintext_s1[37]), .B(signal_3455), .S(n290), 
        .Z(signal_3634) );
  MUX2_X1 cell_587_Ins_0_U1 ( .A(plaintext_s0[38]), .B(signal_1527), .S(n294), 
        .Z(signal_1583) );
  MUX2_X1 cell_587_Ins_1_U1 ( .A(plaintext_s1[38]), .B(signal_3456), .S(n294), 
        .Z(signal_3636) );
  MUX2_X1 cell_588_Ins_0_U1 ( .A(plaintext_s0[39]), .B(signal_1526), .S(n294), 
        .Z(signal_1582) );
  MUX2_X1 cell_588_Ins_1_U1 ( .A(plaintext_s1[39]), .B(signal_3457), .S(n294), 
        .Z(signal_3638) );
  MUX2_X1 cell_589_Ins_0_U1 ( .A(plaintext_s0[24]), .B(ciphertext_s0[16]), .S(
        n287), .Z(signal_1581) );
  MUX2_X1 cell_589_Ins_1_U1 ( .A(plaintext_s1[24]), .B(ciphertext_s1[16]), .S(
        n287), .Z(signal_2778) );
  MUX2_X1 cell_590_Ins_0_U1 ( .A(plaintext_s0[25]), .B(ciphertext_s0[17]), .S(
        n281), .Z(signal_1580) );
  MUX2_X1 cell_590_Ins_1_U1 ( .A(plaintext_s1[25]), .B(ciphertext_s1[17]), .S(
        n281), .Z(signal_2781) );
  MUX2_X1 cell_591_Ins_0_U1 ( .A(plaintext_s0[26]), .B(ciphertext_s0[18]), .S(
        n290), .Z(signal_1579) );
  MUX2_X1 cell_591_Ins_1_U1 ( .A(plaintext_s1[26]), .B(ciphertext_s1[18]), .S(
        n290), .Z(signal_2784) );
  MUX2_X1 cell_592_Ins_0_U1 ( .A(plaintext_s0[27]), .B(ciphertext_s0[19]), .S(
        n35), .Z(signal_1578) );
  MUX2_X1 cell_592_Ins_1_U1 ( .A(plaintext_s1[27]), .B(ciphertext_s1[19]), .S(
        n35), .Z(signal_2787) );
  MUX2_X1 cell_593_Ins_0_U1 ( .A(plaintext_s0[28]), .B(ciphertext_s0[20]), .S(
        n295), .Z(signal_1577) );
  MUX2_X1 cell_593_Ins_1_U1 ( .A(plaintext_s1[28]), .B(ciphertext_s1[20]), .S(
        n295), .Z(signal_2790) );
  MUX2_X1 cell_594_Ins_0_U1 ( .A(plaintext_s0[29]), .B(ciphertext_s0[21]), .S(
        n297), .Z(signal_1576) );
  MUX2_X1 cell_594_Ins_1_U1 ( .A(plaintext_s1[29]), .B(ciphertext_s1[21]), .S(
        n297), .Z(signal_2793) );
  MUX2_X1 cell_595_Ins_0_U1 ( .A(plaintext_s0[30]), .B(ciphertext_s0[22]), .S(
        n298), .Z(signal_1575) );
  MUX2_X1 cell_595_Ins_1_U1 ( .A(plaintext_s1[30]), .B(ciphertext_s1[22]), .S(
        n298), .Z(signal_2796) );
  MUX2_X1 cell_596_Ins_0_U1 ( .A(plaintext_s0[31]), .B(ciphertext_s0[23]), .S(
        n296), .Z(signal_1574) );
  MUX2_X1 cell_596_Ins_1_U1 ( .A(plaintext_s1[31]), .B(ciphertext_s1[23]), .S(
        n296), .Z(signal_2799) );
  MUX2_X1 cell_597_Ins_0_U1 ( .A(plaintext_s0[16]), .B(ciphertext_s0[8]), .S(
        n295), .Z(signal_1573) );
  MUX2_X1 cell_597_Ins_1_U1 ( .A(plaintext_s1[16]), .B(ciphertext_s1[8]), .S(
        n295), .Z(signal_2802) );
  MUX2_X1 cell_598_Ins_0_U1 ( .A(plaintext_s0[17]), .B(ciphertext_s0[9]), .S(
        n303), .Z(signal_1572) );
  MUX2_X1 cell_598_Ins_1_U1 ( .A(plaintext_s1[17]), .B(ciphertext_s1[9]), .S(
        n303), .Z(signal_2805) );
  MUX2_X1 cell_599_Ins_0_U1 ( .A(plaintext_s0[18]), .B(ciphertext_s0[10]), .S(
        n35), .Z(signal_1571) );
  MUX2_X1 cell_599_Ins_1_U1 ( .A(plaintext_s1[18]), .B(ciphertext_s1[10]), .S(
        n35), .Z(signal_2808) );
  MUX2_X1 cell_600_Ins_0_U1 ( .A(plaintext_s0[19]), .B(ciphertext_s0[11]), .S(
        n303), .Z(signal_1570) );
  MUX2_X1 cell_600_Ins_1_U1 ( .A(plaintext_s1[19]), .B(ciphertext_s1[11]), .S(
        n303), .Z(signal_2811) );
  MUX2_X1 cell_601_Ins_0_U1 ( .A(plaintext_s0[20]), .B(ciphertext_s0[12]), .S(
        n305), .Z(signal_1569) );
  MUX2_X1 cell_601_Ins_1_U1 ( .A(plaintext_s1[20]), .B(ciphertext_s1[12]), .S(
        n305), .Z(signal_2814) );
  MUX2_X1 cell_602_Ins_0_U1 ( .A(plaintext_s0[21]), .B(ciphertext_s0[13]), .S(
        n303), .Z(signal_1568) );
  MUX2_X1 cell_602_Ins_1_U1 ( .A(plaintext_s1[21]), .B(ciphertext_s1[13]), .S(
        n303), .Z(signal_2817) );
  MUX2_X1 cell_603_Ins_0_U1 ( .A(plaintext_s0[22]), .B(ciphertext_s0[14]), .S(
        n305), .Z(signal_1567) );
  MUX2_X1 cell_603_Ins_1_U1 ( .A(plaintext_s1[22]), .B(ciphertext_s1[14]), .S(
        n305), .Z(signal_2820) );
  MUX2_X1 cell_604_Ins_0_U1 ( .A(plaintext_s0[23]), .B(ciphertext_s0[15]), .S(
        n305), .Z(signal_1566) );
  MUX2_X1 cell_604_Ins_1_U1 ( .A(plaintext_s1[23]), .B(ciphertext_s1[15]), .S(
        n305), .Z(signal_2823) );
  MUX2_X1 cell_605_Ins_0_U1 ( .A(plaintext_s0[8]), .B(ciphertext_s0[0]), .S(
        n296), .Z(signal_1565) );
  MUX2_X1 cell_605_Ins_1_U1 ( .A(plaintext_s1[8]), .B(ciphertext_s1[0]), .S(
        n296), .Z(signal_2826) );
  MUX2_X1 cell_606_Ins_0_U1 ( .A(plaintext_s0[9]), .B(ciphertext_s0[1]), .S(
        n285), .Z(signal_1564) );
  MUX2_X1 cell_606_Ins_1_U1 ( .A(plaintext_s1[9]), .B(ciphertext_s1[1]), .S(
        n285), .Z(signal_2829) );
  MUX2_X1 cell_607_Ins_0_U1 ( .A(plaintext_s0[10]), .B(ciphertext_s0[2]), .S(
        n284), .Z(signal_1563) );
  MUX2_X1 cell_607_Ins_1_U1 ( .A(plaintext_s1[10]), .B(ciphertext_s1[2]), .S(
        n284), .Z(signal_2832) );
  MUX2_X1 cell_608_Ins_0_U1 ( .A(plaintext_s0[11]), .B(ciphertext_s0[3]), .S(
        n280), .Z(signal_1562) );
  MUX2_X1 cell_608_Ins_1_U1 ( .A(plaintext_s1[11]), .B(ciphertext_s1[3]), .S(
        n280), .Z(signal_2835) );
  MUX2_X1 cell_609_Ins_0_U1 ( .A(plaintext_s0[12]), .B(ciphertext_s0[4]), .S(
        n286), .Z(signal_1561) );
  MUX2_X1 cell_609_Ins_1_U1 ( .A(plaintext_s1[12]), .B(ciphertext_s1[4]), .S(
        n286), .Z(signal_2838) );
  MUX2_X1 cell_610_Ins_0_U1 ( .A(plaintext_s0[13]), .B(ciphertext_s0[5]), .S(
        n301), .Z(signal_1560) );
  MUX2_X1 cell_610_Ins_1_U1 ( .A(plaintext_s1[13]), .B(ciphertext_s1[5]), .S(
        n301), .Z(signal_2841) );
  MUX2_X1 cell_611_Ins_0_U1 ( .A(plaintext_s0[14]), .B(ciphertext_s0[6]), .S(
        n304), .Z(signal_1559) );
  MUX2_X1 cell_611_Ins_1_U1 ( .A(plaintext_s1[14]), .B(ciphertext_s1[6]), .S(
        n304), .Z(signal_2844) );
  MUX2_X1 cell_612_Ins_0_U1 ( .A(plaintext_s0[15]), .B(ciphertext_s0[7]), .S(
        n297), .Z(signal_1558) );
  MUX2_X1 cell_612_Ins_1_U1 ( .A(plaintext_s1[15]), .B(ciphertext_s1[7]), .S(
        n297), .Z(signal_2847) );
  MUX2_X1 cell_632_Ins_0_U1 ( .A(signal_1485), .B(ciphertext_s0[24]), .S(n470), 
        .Z(signal_1453) );
  MUX2_X1 cell_632_Ins_1_U1 ( .A(signal_3231), .B(ciphertext_s1[24]), .S(n470), 
        .Z(signal_3262) );
  MUX2_X1 cell_633_Ins_0_U1 ( .A(signal_1484), .B(ciphertext_s0[25]), .S(n473), 
        .Z(signal_1452) );
  MUX2_X1 cell_633_Ins_1_U1 ( .A(signal_3255), .B(ciphertext_s1[25]), .S(n473), 
        .Z(signal_3263) );
  MUX2_X1 cell_634_Ins_0_U1 ( .A(signal_1483), .B(ciphertext_s0[26]), .S(n471), 
        .Z(signal_1451) );
  MUX2_X1 cell_634_Ins_1_U1 ( .A(signal_3229), .B(ciphertext_s1[26]), .S(n471), 
        .Z(signal_3240) );
  MUX2_X1 cell_635_Ins_0_U1 ( .A(signal_1482), .B(ciphertext_s0[27]), .S(n472), 
        .Z(signal_1450) );
  MUX2_X1 cell_635_Ins_1_U1 ( .A(signal_3254), .B(ciphertext_s1[27]), .S(n472), 
        .Z(signal_3264) );
  MUX2_X1 cell_636_Ins_0_U1 ( .A(signal_1481), .B(ciphertext_s0[28]), .S(
        signal_399), .Z(signal_1449) );
  MUX2_X1 cell_636_Ins_1_U1 ( .A(signal_3253), .B(ciphertext_s1[28]), .S(
        signal_399), .Z(signal_3265) );
  MUX2_X1 cell_637_Ins_0_U1 ( .A(signal_1480), .B(ciphertext_s0[29]), .S(
        signal_399), .Z(signal_1448) );
  MUX2_X1 cell_637_Ins_1_U1 ( .A(signal_3226), .B(ciphertext_s1[29]), .S(
        signal_399), .Z(signal_3241) );
  MUX2_X1 cell_638_Ins_0_U1 ( .A(signal_1479), .B(ciphertext_s0[30]), .S(
        signal_399), .Z(signal_1447) );
  MUX2_X1 cell_638_Ins_1_U1 ( .A(signal_3225), .B(ciphertext_s1[30]), .S(
        signal_399), .Z(signal_3242) );
  MUX2_X1 cell_639_Ins_0_U1 ( .A(signal_1478), .B(ciphertext_s0[31]), .S(n470), 
        .Z(signal_1446) );
  MUX2_X1 cell_639_Ins_1_U1 ( .A(signal_3224), .B(ciphertext_s1[31]), .S(n470), 
        .Z(signal_3243) );
  MUX2_X1 cell_640_Ins_0_U1 ( .A(signal_1477), .B(ciphertext_s0[56]), .S(n470), 
        .Z(signal_1445) );
  MUX2_X1 cell_640_Ins_1_U1 ( .A(signal_3223), .B(ciphertext_s1[56]), .S(n470), 
        .Z(signal_3266) );
  MUX2_X1 cell_641_Ins_0_U1 ( .A(signal_1476), .B(ciphertext_s0[57]), .S(n470), 
        .Z(signal_1444) );
  MUX2_X1 cell_641_Ins_1_U1 ( .A(signal_3252), .B(ciphertext_s1[57]), .S(n470), 
        .Z(signal_3267) );
  MUX2_X1 cell_642_Ins_0_U1 ( .A(signal_1475), .B(ciphertext_s0[58]), .S(n470), 
        .Z(signal_1443) );
  MUX2_X1 cell_642_Ins_1_U1 ( .A(signal_3221), .B(ciphertext_s1[58]), .S(n470), 
        .Z(signal_3268) );
  MUX2_X1 cell_643_Ins_0_U1 ( .A(signal_1474), .B(ciphertext_s0[59]), .S(n470), 
        .Z(signal_1442) );
  MUX2_X1 cell_643_Ins_1_U1 ( .A(signal_3251), .B(ciphertext_s1[59]), .S(n470), 
        .Z(signal_3269) );
  MUX2_X1 cell_644_Ins_0_U1 ( .A(signal_1473), .B(ciphertext_s0[60]), .S(n470), 
        .Z(signal_1441) );
  MUX2_X1 cell_644_Ins_1_U1 ( .A(signal_3250), .B(ciphertext_s1[60]), .S(n470), 
        .Z(signal_3270) );
  MUX2_X1 cell_645_Ins_0_U1 ( .A(signal_1472), .B(ciphertext_s0[61]), .S(n470), 
        .Z(signal_1440) );
  MUX2_X1 cell_645_Ins_1_U1 ( .A(signal_3218), .B(ciphertext_s1[61]), .S(n470), 
        .Z(signal_3271) );
  MUX2_X1 cell_646_Ins_0_U1 ( .A(signal_1471), .B(ciphertext_s0[62]), .S(n471), 
        .Z(signal_1439) );
  MUX2_X1 cell_646_Ins_1_U1 ( .A(signal_3217), .B(ciphertext_s1[62]), .S(n471), 
        .Z(signal_3272) );
  MUX2_X1 cell_647_Ins_0_U1 ( .A(signal_1470), .B(ciphertext_s0[63]), .S(n471), 
        .Z(signal_1438) );
  MUX2_X1 cell_647_Ins_1_U1 ( .A(signal_3216), .B(ciphertext_s1[63]), .S(n471), 
        .Z(signal_3273) );
  MUX2_X1 cell_648_Ins_0_U1 ( .A(signal_1469), .B(ciphertext_s0[88]), .S(n471), 
        .Z(signal_1437) );
  MUX2_X1 cell_648_Ins_1_U1 ( .A(signal_3215), .B(ciphertext_s1[88]), .S(n471), 
        .Z(signal_3274) );
  MUX2_X1 cell_649_Ins_0_U1 ( .A(signal_1468), .B(ciphertext_s0[89]), .S(n471), 
        .Z(signal_1436) );
  MUX2_X1 cell_649_Ins_1_U1 ( .A(signal_3249), .B(ciphertext_s1[89]), .S(n471), 
        .Z(signal_3275) );
  MUX2_X1 cell_650_Ins_0_U1 ( .A(signal_1467), .B(ciphertext_s0[90]), .S(n471), 
        .Z(signal_1435) );
  MUX2_X1 cell_650_Ins_1_U1 ( .A(signal_3213), .B(ciphertext_s1[90]), .S(n471), 
        .Z(signal_3276) );
  MUX2_X1 cell_651_Ins_0_U1 ( .A(signal_1466), .B(ciphertext_s0[91]), .S(n471), 
        .Z(signal_1434) );
  MUX2_X1 cell_651_Ins_1_U1 ( .A(signal_3248), .B(ciphertext_s1[91]), .S(n471), 
        .Z(signal_3277) );
  MUX2_X1 cell_652_Ins_0_U1 ( .A(signal_1465), .B(ciphertext_s0[92]), .S(n471), 
        .Z(signal_1433) );
  MUX2_X1 cell_652_Ins_1_U1 ( .A(signal_3247), .B(ciphertext_s1[92]), .S(n471), 
        .Z(signal_3278) );
  MUX2_X1 cell_653_Ins_0_U1 ( .A(signal_1464), .B(ciphertext_s0[93]), .S(n472), 
        .Z(signal_1432) );
  MUX2_X1 cell_653_Ins_1_U1 ( .A(signal_3210), .B(ciphertext_s1[93]), .S(n472), 
        .Z(signal_3279) );
  MUX2_X1 cell_654_Ins_0_U1 ( .A(signal_1463), .B(ciphertext_s0[94]), .S(n472), 
        .Z(signal_1431) );
  MUX2_X1 cell_654_Ins_1_U1 ( .A(signal_3209), .B(ciphertext_s1[94]), .S(n472), 
        .Z(signal_3280) );
  MUX2_X1 cell_655_Ins_0_U1 ( .A(signal_1462), .B(ciphertext_s0[95]), .S(n472), 
        .Z(signal_1430) );
  MUX2_X1 cell_655_Ins_1_U1 ( .A(signal_3208), .B(ciphertext_s1[95]), .S(n472), 
        .Z(signal_3281) );
  MUX2_X1 cell_656_Ins_0_U1 ( .A(signal_1461), .B(ciphertext_s0[120]), .S(n472), .Z(signal_1429) );
  MUX2_X1 cell_656_Ins_1_U1 ( .A(signal_3207), .B(ciphertext_s1[120]), .S(n472), .Z(signal_3282) );
  MUX2_X1 cell_657_Ins_0_U1 ( .A(signal_1460), .B(ciphertext_s0[121]), .S(n472), .Z(signal_1428) );
  MUX2_X1 cell_657_Ins_1_U1 ( .A(signal_3246), .B(ciphertext_s1[121]), .S(n472), .Z(signal_3283) );
  MUX2_X1 cell_658_Ins_0_U1 ( .A(signal_1459), .B(ciphertext_s0[122]), .S(n472), .Z(signal_1427) );
  MUX2_X1 cell_658_Ins_1_U1 ( .A(signal_3205), .B(ciphertext_s1[122]), .S(n472), .Z(signal_3284) );
  MUX2_X1 cell_659_Ins_0_U1 ( .A(signal_1458), .B(ciphertext_s0[123]), .S(n472), .Z(signal_1426) );
  MUX2_X1 cell_659_Ins_1_U1 ( .A(signal_3245), .B(ciphertext_s1[123]), .S(n472), .Z(signal_3285) );
  MUX2_X1 cell_660_Ins_0_U1 ( .A(signal_1457), .B(ciphertext_s0[124]), .S(n473), .Z(signal_1425) );
  MUX2_X1 cell_660_Ins_1_U1 ( .A(signal_3244), .B(ciphertext_s1[124]), .S(n473), .Z(signal_3286) );
  MUX2_X1 cell_661_Ins_0_U1 ( .A(signal_1456), .B(ciphertext_s0[125]), .S(n473), .Z(signal_1424) );
  MUX2_X1 cell_661_Ins_1_U1 ( .A(signal_3202), .B(ciphertext_s1[125]), .S(n473), .Z(signal_3287) );
  MUX2_X1 cell_662_Ins_0_U1 ( .A(signal_1455), .B(ciphertext_s0[126]), .S(n473), .Z(signal_1423) );
  MUX2_X1 cell_662_Ins_1_U1 ( .A(signal_3201), .B(ciphertext_s1[126]), .S(n473), .Z(signal_3288) );
  MUX2_X1 cell_663_Ins_0_U1 ( .A(signal_1454), .B(ciphertext_s0[127]), .S(n473), .Z(signal_1422) );
  MUX2_X1 cell_663_Ins_1_U1 ( .A(signal_3200), .B(ciphertext_s1[127]), .S(n473), .Z(signal_3289) );
  XOR2_X1 cell_664_Ins_0_U1 ( .A(signal_765), .B(signal_1486), .Z(signal_1686)
         );
  XOR2_X1 cell_664_Ins_1_U1 ( .A(signal_2412), .B(signal_2410), .Z(signal_2413) );
  XOR2_X1 cell_665_Ins_0_U1 ( .A(signal_764), .B(signal_1487), .Z(signal_1687)
         );
  XOR2_X1 cell_665_Ins_1_U1 ( .A(signal_2414), .B(signal_2407), .Z(signal_2415) );
  XOR2_X1 cell_666_Ins_0_U1 ( .A(signal_763), .B(signal_1488), .Z(signal_1688)
         );
  XOR2_X1 cell_666_Ins_1_U1 ( .A(signal_2416), .B(signal_2404), .Z(signal_2417) );
  XOR2_X1 cell_667_Ins_0_U1 ( .A(signal_762), .B(signal_1489), .Z(signal_1689)
         );
  XOR2_X1 cell_667_Ins_1_U1 ( .A(signal_2418), .B(signal_2401), .Z(signal_2419) );
  XOR2_X1 cell_668_Ins_0_U1 ( .A(signal_761), .B(signal_1490), .Z(signal_1690)
         );
  XOR2_X1 cell_668_Ins_1_U1 ( .A(signal_2420), .B(signal_2398), .Z(signal_2421) );
  XOR2_X1 cell_669_Ins_0_U1 ( .A(signal_760), .B(signal_1491), .Z(signal_1691)
         );
  XOR2_X1 cell_669_Ins_1_U1 ( .A(signal_2422), .B(signal_2395), .Z(signal_2423) );
  XOR2_X1 cell_670_Ins_0_U1 ( .A(signal_759), .B(signal_1492), .Z(signal_1692)
         );
  XOR2_X1 cell_670_Ins_1_U1 ( .A(signal_2424), .B(signal_2392), .Z(signal_2425) );
  XOR2_X1 cell_671_Ins_0_U1 ( .A(signal_758), .B(signal_1493), .Z(signal_1693)
         );
  XOR2_X1 cell_671_Ins_1_U1 ( .A(signal_2426), .B(signal_2389), .Z(signal_2427) );
  MUX2_X1 cell_714_Ins_0_U1 ( .A(signal_1493), .B(signal_767), .S(n330), .Z(
        signal_766) );
  MUX2_X1 cell_714_Ins_1_U1 ( .A(signal_2389), .B(signal_3986), .S(n330), .Z(
        signal_4122) );
  MUX2_X1 cell_715_Ins_0_U1 ( .A(signal_1933), .B(signal_1877), .S(n309), .Z(
        signal_767) );
  MUX2_X1 cell_715_Ins_1_U1 ( .A(signal_3907), .B(signal_2897), .S(n309), .Z(
        signal_3986) );
  MUX2_X1 cell_718_Ins_0_U1 ( .A(signal_1492), .B(signal_770), .S(n330), .Z(
        signal_769) );
  MUX2_X1 cell_718_Ins_1_U1 ( .A(signal_2392), .B(signal_3987), .S(n330), .Z(
        signal_4123) );
  MUX2_X1 cell_719_Ins_0_U1 ( .A(signal_1932), .B(signal_1876), .S(n309), .Z(
        signal_770) );
  MUX2_X1 cell_719_Ins_1_U1 ( .A(signal_3909), .B(signal_2900), .S(n309), .Z(
        signal_3987) );
  MUX2_X1 cell_722_Ins_0_U1 ( .A(signal_1491), .B(signal_773), .S(n337), .Z(
        signal_772) );
  MUX2_X1 cell_722_Ins_1_U1 ( .A(signal_2395), .B(signal_3988), .S(n337), .Z(
        signal_4124) );
  MUX2_X1 cell_723_Ins_0_U1 ( .A(signal_1931), .B(signal_1875), .S(n309), .Z(
        signal_773) );
  MUX2_X1 cell_723_Ins_1_U1 ( .A(signal_3911), .B(signal_2903), .S(n309), .Z(
        signal_3988) );
  MUX2_X1 cell_726_Ins_0_U1 ( .A(signal_1490), .B(signal_776), .S(n326), .Z(
        signal_775) );
  MUX2_X1 cell_726_Ins_1_U1 ( .A(signal_2398), .B(signal_3989), .S(n326), .Z(
        signal_4125) );
  MUX2_X1 cell_727_Ins_0_U1 ( .A(signal_1930), .B(signal_1874), .S(n309), .Z(
        signal_776) );
  MUX2_X1 cell_727_Ins_1_U1 ( .A(signal_3913), .B(signal_2906), .S(n309), .Z(
        signal_3989) );
  MUX2_X1 cell_730_Ins_0_U1 ( .A(signal_1489), .B(signal_779), .S(n337), .Z(
        signal_778) );
  MUX2_X1 cell_730_Ins_1_U1 ( .A(signal_2401), .B(signal_3990), .S(n337), .Z(
        signal_4126) );
  MUX2_X1 cell_731_Ins_0_U1 ( .A(signal_1929), .B(signal_1873), .S(n310), .Z(
        signal_779) );
  MUX2_X1 cell_731_Ins_1_U1 ( .A(signal_3915), .B(signal_2909), .S(n310), .Z(
        signal_3990) );
  MUX2_X1 cell_734_Ins_0_U1 ( .A(signal_1488), .B(signal_782), .S(n337), .Z(
        signal_781) );
  MUX2_X1 cell_734_Ins_1_U1 ( .A(signal_2404), .B(signal_3991), .S(n337), .Z(
        signal_4127) );
  MUX2_X1 cell_735_Ins_0_U1 ( .A(signal_1928), .B(signal_1872), .S(n310), .Z(
        signal_782) );
  MUX2_X1 cell_735_Ins_1_U1 ( .A(signal_3917), .B(signal_2912), .S(n310), .Z(
        signal_3991) );
  MUX2_X1 cell_738_Ins_0_U1 ( .A(signal_1487), .B(signal_785), .S(n337), .Z(
        signal_784) );
  MUX2_X1 cell_738_Ins_1_U1 ( .A(signal_2407), .B(signal_3992), .S(n337), .Z(
        signal_4128) );
  MUX2_X1 cell_739_Ins_0_U1 ( .A(signal_1927), .B(signal_1871), .S(n310), .Z(
        signal_785) );
  MUX2_X1 cell_739_Ins_1_U1 ( .A(signal_3919), .B(signal_2915), .S(n310), .Z(
        signal_3992) );
  MUX2_X1 cell_742_Ins_0_U1 ( .A(signal_1486), .B(signal_788), .S(n337), .Z(
        signal_787) );
  MUX2_X1 cell_742_Ins_1_U1 ( .A(signal_2410), .B(signal_3993), .S(n337), .Z(
        signal_4129) );
  MUX2_X1 cell_743_Ins_0_U1 ( .A(signal_1926), .B(signal_1870), .S(n310), .Z(
        signal_788) );
  MUX2_X1 cell_743_Ins_1_U1 ( .A(signal_3921), .B(signal_2918), .S(n310), .Z(
        signal_3993) );
  MUX2_X1 cell_746_Ins_0_U1 ( .A(signal_758), .B(signal_791), .S(n337), .Z(
        signal_790) );
  MUX2_X1 cell_746_Ins_1_U1 ( .A(signal_2426), .B(signal_3290), .S(n337), .Z(
        signal_3994) );
  MUX2_X1 cell_747_Ins_0_U1 ( .A(signal_1925), .B(signal_1861), .S(n310), .Z(
        signal_791) );
  MUX2_X1 cell_747_Ins_1_U1 ( .A(signal_2850), .B(signal_2921), .S(n310), .Z(
        signal_3290) );
  MUX2_X1 cell_750_Ins_0_U1 ( .A(signal_759), .B(signal_794), .S(n337), .Z(
        signal_793) );
  MUX2_X1 cell_750_Ins_1_U1 ( .A(signal_2424), .B(signal_3291), .S(n337), .Z(
        signal_3995) );
  MUX2_X1 cell_751_Ins_0_U1 ( .A(signal_1924), .B(signal_1860), .S(n310), .Z(
        signal_794) );
  MUX2_X1 cell_751_Ins_1_U1 ( .A(signal_2853), .B(signal_2924), .S(n310), .Z(
        signal_3291) );
  MUX2_X1 cell_754_Ins_0_U1 ( .A(signal_760), .B(signal_797), .S(n336), .Z(
        signal_796) );
  MUX2_X1 cell_754_Ins_1_U1 ( .A(signal_2422), .B(signal_3292), .S(n336), .Z(
        signal_3996) );
  MUX2_X1 cell_755_Ins_0_U1 ( .A(signal_1923), .B(signal_1859), .S(n310), .Z(
        signal_797) );
  MUX2_X1 cell_755_Ins_1_U1 ( .A(signal_2856), .B(signal_2927), .S(n310), .Z(
        signal_3292) );
  MUX2_X1 cell_758_Ins_0_U1 ( .A(signal_761), .B(signal_800), .S(n336), .Z(
        signal_799) );
  MUX2_X1 cell_758_Ins_1_U1 ( .A(signal_2420), .B(signal_3293), .S(n336), .Z(
        signal_3997) );
  MUX2_X1 cell_759_Ins_0_U1 ( .A(signal_1922), .B(signal_1858), .S(n311), .Z(
        signal_800) );
  MUX2_X1 cell_759_Ins_1_U1 ( .A(signal_2859), .B(signal_2930), .S(n311), .Z(
        signal_3293) );
  MUX2_X1 cell_762_Ins_0_U1 ( .A(signal_762), .B(signal_803), .S(n336), .Z(
        signal_802) );
  MUX2_X1 cell_762_Ins_1_U1 ( .A(signal_2418), .B(signal_3294), .S(n336), .Z(
        signal_3998) );
  MUX2_X1 cell_763_Ins_0_U1 ( .A(signal_1921), .B(signal_1857), .S(n311), .Z(
        signal_803) );
  MUX2_X1 cell_763_Ins_1_U1 ( .A(signal_2862), .B(signal_2933), .S(n311), .Z(
        signal_3294) );
  MUX2_X1 cell_766_Ins_0_U1 ( .A(signal_763), .B(signal_806), .S(n336), .Z(
        signal_805) );
  MUX2_X1 cell_766_Ins_1_U1 ( .A(signal_2416), .B(signal_3295), .S(n336), .Z(
        signal_3999) );
  MUX2_X1 cell_767_Ins_0_U1 ( .A(signal_1920), .B(signal_1856), .S(n311), .Z(
        signal_806) );
  MUX2_X1 cell_767_Ins_1_U1 ( .A(signal_2865), .B(signal_2936), .S(n311), .Z(
        signal_3295) );
  MUX2_X1 cell_770_Ins_0_U1 ( .A(signal_764), .B(signal_809), .S(n336), .Z(
        signal_808) );
  MUX2_X1 cell_770_Ins_1_U1 ( .A(signal_2414), .B(signal_3296), .S(n336), .Z(
        signal_4000) );
  MUX2_X1 cell_771_Ins_0_U1 ( .A(signal_1919), .B(signal_1855), .S(n311), .Z(
        signal_809) );
  MUX2_X1 cell_771_Ins_1_U1 ( .A(signal_2868), .B(signal_2939), .S(n311), .Z(
        signal_3296) );
  MUX2_X1 cell_774_Ins_0_U1 ( .A(signal_765), .B(signal_812), .S(n336), .Z(
        signal_811) );
  MUX2_X1 cell_774_Ins_1_U1 ( .A(signal_2412), .B(signal_3297), .S(n336), .Z(
        signal_4001) );
  MUX2_X1 cell_775_Ins_0_U1 ( .A(signal_1918), .B(signal_1854), .S(n311), .Z(
        signal_812) );
  MUX2_X1 cell_775_Ins_1_U1 ( .A(signal_2871), .B(signal_2942), .S(n311), .Z(
        signal_3297) );
  MUX2_X1 cell_778_Ins_0_U1 ( .A(signal_1909), .B(signal_815), .S(n335), .Z(
        signal_814) );
  MUX2_X1 cell_778_Ins_1_U1 ( .A(signal_2849), .B(signal_3298), .S(n335), .Z(
        signal_4002) );
  MUX2_X1 cell_779_Ins_0_U1 ( .A(signal_1917), .B(signal_1845), .S(n311), .Z(
        signal_815) );
  MUX2_X1 cell_779_Ins_1_U1 ( .A(signal_2874), .B(signal_2945), .S(n311), .Z(
        signal_3298) );
  MUX2_X1 cell_782_Ins_0_U1 ( .A(signal_1908), .B(signal_818), .S(n336), .Z(
        signal_817) );
  MUX2_X1 cell_782_Ins_1_U1 ( .A(signal_2852), .B(signal_3299), .S(n336), .Z(
        signal_4003) );
  MUX2_X1 cell_783_Ins_0_U1 ( .A(signal_1916), .B(signal_1844), .S(n311), .Z(
        signal_818) );
  MUX2_X1 cell_783_Ins_1_U1 ( .A(signal_2877), .B(signal_2948), .S(n311), .Z(
        signal_3299) );
  MUX2_X1 cell_786_Ins_0_U1 ( .A(signal_1907), .B(signal_821), .S(n335), .Z(
        signal_820) );
  MUX2_X1 cell_786_Ins_1_U1 ( .A(signal_2855), .B(signal_3300), .S(n335), .Z(
        signal_4004) );
  MUX2_X1 cell_787_Ins_0_U1 ( .A(signal_1915), .B(signal_1843), .S(n312), .Z(
        signal_821) );
  MUX2_X1 cell_787_Ins_1_U1 ( .A(signal_2880), .B(signal_2951), .S(n312), .Z(
        signal_3300) );
  MUX2_X1 cell_790_Ins_0_U1 ( .A(signal_1906), .B(signal_824), .S(n335), .Z(
        signal_823) );
  MUX2_X1 cell_790_Ins_1_U1 ( .A(signal_2858), .B(signal_3301), .S(n335), .Z(
        signal_4005) );
  MUX2_X1 cell_791_Ins_0_U1 ( .A(signal_1914), .B(signal_1842), .S(n312), .Z(
        signal_824) );
  MUX2_X1 cell_791_Ins_1_U1 ( .A(signal_2883), .B(signal_2954), .S(n312), .Z(
        signal_3301) );
  MUX2_X1 cell_794_Ins_0_U1 ( .A(signal_1905), .B(signal_827), .S(n335), .Z(
        signal_826) );
  MUX2_X1 cell_794_Ins_1_U1 ( .A(signal_2861), .B(signal_3302), .S(n335), .Z(
        signal_4006) );
  MUX2_X1 cell_795_Ins_0_U1 ( .A(signal_1913), .B(signal_1841), .S(n312), .Z(
        signal_827) );
  MUX2_X1 cell_795_Ins_1_U1 ( .A(signal_2886), .B(signal_2957), .S(n312), .Z(
        signal_3302) );
  MUX2_X1 cell_798_Ins_0_U1 ( .A(signal_1904), .B(signal_830), .S(n335), .Z(
        signal_829) );
  MUX2_X1 cell_798_Ins_1_U1 ( .A(signal_2864), .B(signal_3303), .S(n335), .Z(
        signal_4007) );
  MUX2_X1 cell_799_Ins_0_U1 ( .A(signal_1912), .B(signal_1840), .S(n312), .Z(
        signal_830) );
  MUX2_X1 cell_799_Ins_1_U1 ( .A(signal_2889), .B(signal_2960), .S(n312), .Z(
        signal_3303) );
  MUX2_X1 cell_802_Ins_0_U1 ( .A(signal_1903), .B(signal_833), .S(n335), .Z(
        signal_832) );
  MUX2_X1 cell_802_Ins_1_U1 ( .A(signal_2867), .B(signal_3304), .S(n335), .Z(
        signal_4008) );
  MUX2_X1 cell_803_Ins_0_U1 ( .A(signal_1911), .B(signal_1839), .S(n312), .Z(
        signal_833) );
  MUX2_X1 cell_803_Ins_1_U1 ( .A(signal_2892), .B(signal_2963), .S(n312), .Z(
        signal_3304) );
  MUX2_X1 cell_806_Ins_0_U1 ( .A(signal_1902), .B(signal_836), .S(n335), .Z(
        signal_835) );
  MUX2_X1 cell_806_Ins_1_U1 ( .A(signal_2870), .B(signal_3305), .S(n335), .Z(
        signal_4009) );
  MUX2_X1 cell_807_Ins_0_U1 ( .A(signal_1910), .B(signal_1838), .S(n312), .Z(
        signal_836) );
  MUX2_X1 cell_807_Ins_1_U1 ( .A(signal_2895), .B(signal_2966), .S(n312), .Z(
        signal_3305) );
  MUX2_X1 cell_810_Ins_0_U1 ( .A(signal_1893), .B(signal_839), .S(n334), .Z(
        signal_838) );
  MUX2_X1 cell_810_Ins_1_U1 ( .A(signal_2873), .B(signal_3306), .S(n334), .Z(
        signal_4010) );
  MUX2_X1 cell_811_Ins_0_U1 ( .A(signal_1901), .B(signal_1509), .S(n312), .Z(
        signal_839) );
  MUX2_X1 cell_811_Ins_1_U1 ( .A(signal_2898), .B(signal_2969), .S(n312), .Z(
        signal_3306) );
  MUX2_X1 cell_814_Ins_0_U1 ( .A(signal_1892), .B(signal_842), .S(n334), .Z(
        signal_841) );
  MUX2_X1 cell_814_Ins_1_U1 ( .A(signal_2876), .B(signal_3307), .S(n334), .Z(
        signal_4011) );
  MUX2_X1 cell_815_Ins_0_U1 ( .A(signal_1900), .B(signal_1508), .S(n313), .Z(
        signal_842) );
  MUX2_X1 cell_815_Ins_1_U1 ( .A(signal_2901), .B(signal_2972), .S(n313), .Z(
        signal_3307) );
  MUX2_X1 cell_818_Ins_0_U1 ( .A(signal_1891), .B(signal_845), .S(n334), .Z(
        signal_844) );
  MUX2_X1 cell_818_Ins_1_U1 ( .A(signal_2879), .B(signal_3308), .S(n334), .Z(
        signal_4012) );
  MUX2_X1 cell_819_Ins_0_U1 ( .A(signal_1899), .B(signal_1507), .S(n313), .Z(
        signal_845) );
  MUX2_X1 cell_819_Ins_1_U1 ( .A(signal_2904), .B(signal_2975), .S(n313), .Z(
        signal_3308) );
  MUX2_X1 cell_822_Ins_0_U1 ( .A(signal_1890), .B(signal_848), .S(n334), .Z(
        signal_847) );
  MUX2_X1 cell_822_Ins_1_U1 ( .A(signal_2882), .B(signal_3309), .S(n334), .Z(
        signal_4013) );
  MUX2_X1 cell_823_Ins_0_U1 ( .A(signal_1898), .B(signal_1506), .S(n313), .Z(
        signal_848) );
  MUX2_X1 cell_823_Ins_1_U1 ( .A(signal_2907), .B(signal_2978), .S(n313), .Z(
        signal_3309) );
  MUX2_X1 cell_826_Ins_0_U1 ( .A(signal_1889), .B(signal_851), .S(n334), .Z(
        signal_850) );
  MUX2_X1 cell_826_Ins_1_U1 ( .A(signal_2885), .B(signal_3310), .S(n334), .Z(
        signal_4014) );
  MUX2_X1 cell_827_Ins_0_U1 ( .A(signal_1897), .B(signal_1505), .S(n313), .Z(
        signal_851) );
  MUX2_X1 cell_827_Ins_1_U1 ( .A(signal_2910), .B(signal_2981), .S(n313), .Z(
        signal_3310) );
  MUX2_X1 cell_830_Ins_0_U1 ( .A(signal_1888), .B(signal_854), .S(n334), .Z(
        signal_853) );
  MUX2_X1 cell_830_Ins_1_U1 ( .A(signal_2888), .B(signal_3311), .S(n334), .Z(
        signal_4015) );
  MUX2_X1 cell_831_Ins_0_U1 ( .A(signal_1896), .B(signal_1504), .S(n313), .Z(
        signal_854) );
  MUX2_X1 cell_831_Ins_1_U1 ( .A(signal_2913), .B(signal_2984), .S(n313), .Z(
        signal_3311) );
  MUX2_X1 cell_834_Ins_0_U1 ( .A(signal_1887), .B(signal_857), .S(n334), .Z(
        signal_856) );
  MUX2_X1 cell_834_Ins_1_U1 ( .A(signal_2891), .B(signal_3312), .S(n334), .Z(
        signal_4016) );
  MUX2_X1 cell_835_Ins_0_U1 ( .A(signal_1895), .B(signal_1503), .S(n313), .Z(
        signal_857) );
  MUX2_X1 cell_835_Ins_1_U1 ( .A(signal_2916), .B(signal_2987), .S(n313), .Z(
        signal_3312) );
  MUX2_X1 cell_838_Ins_0_U1 ( .A(signal_1886), .B(signal_860), .S(n333), .Z(
        signal_859) );
  MUX2_X1 cell_838_Ins_1_U1 ( .A(signal_2894), .B(signal_3313), .S(n333), .Z(
        signal_4017) );
  MUX2_X1 cell_839_Ins_0_U1 ( .A(signal_1894), .B(signal_1502), .S(n313), .Z(
        signal_860) );
  MUX2_X1 cell_839_Ins_1_U1 ( .A(signal_2919), .B(signal_2990), .S(n313), .Z(
        signal_3313) );
  MUX2_X1 cell_842_Ins_0_U1 ( .A(signal_1877), .B(signal_863), .S(n333), .Z(
        signal_862) );
  MUX2_X1 cell_842_Ins_1_U1 ( .A(signal_2897), .B(signal_3314), .S(n333), .Z(
        signal_4018) );
  MUX2_X1 cell_843_Ins_0_U1 ( .A(signal_1885), .B(signal_1821), .S(n314), .Z(
        signal_863) );
  MUX2_X1 cell_843_Ins_1_U1 ( .A(signal_2922), .B(signal_2993), .S(n314), .Z(
        signal_3314) );
  MUX2_X1 cell_846_Ins_0_U1 ( .A(signal_1876), .B(signal_866), .S(n333), .Z(
        signal_865) );
  MUX2_X1 cell_846_Ins_1_U1 ( .A(signal_2900), .B(signal_3315), .S(n333), .Z(
        signal_4019) );
  MUX2_X1 cell_847_Ins_0_U1 ( .A(signal_1884), .B(signal_1820), .S(n314), .Z(
        signal_866) );
  MUX2_X1 cell_847_Ins_1_U1 ( .A(signal_2925), .B(signal_2996), .S(n314), .Z(
        signal_3315) );
  MUX2_X1 cell_850_Ins_0_U1 ( .A(signal_1875), .B(signal_869), .S(n333), .Z(
        signal_868) );
  MUX2_X1 cell_850_Ins_1_U1 ( .A(signal_2903), .B(signal_3316), .S(n333), .Z(
        signal_4020) );
  MUX2_X1 cell_851_Ins_0_U1 ( .A(signal_1883), .B(signal_1819), .S(n314), .Z(
        signal_869) );
  MUX2_X1 cell_851_Ins_1_U1 ( .A(signal_2928), .B(signal_2999), .S(n314), .Z(
        signal_3316) );
  MUX2_X1 cell_854_Ins_0_U1 ( .A(signal_1874), .B(signal_872), .S(n333), .Z(
        signal_871) );
  MUX2_X1 cell_854_Ins_1_U1 ( .A(signal_2906), .B(signal_3317), .S(n333), .Z(
        signal_4021) );
  MUX2_X1 cell_855_Ins_0_U1 ( .A(signal_1882), .B(signal_1818), .S(n314), .Z(
        signal_872) );
  MUX2_X1 cell_855_Ins_1_U1 ( .A(signal_2931), .B(signal_3002), .S(n314), .Z(
        signal_3317) );
  MUX2_X1 cell_858_Ins_0_U1 ( .A(signal_1873), .B(signal_875), .S(n333), .Z(
        signal_874) );
  MUX2_X1 cell_858_Ins_1_U1 ( .A(signal_2909), .B(signal_3318), .S(n333), .Z(
        signal_4022) );
  MUX2_X1 cell_859_Ins_0_U1 ( .A(signal_1881), .B(signal_1817), .S(n314), .Z(
        signal_875) );
  MUX2_X1 cell_859_Ins_1_U1 ( .A(signal_2934), .B(signal_3005), .S(n314), .Z(
        signal_3318) );
  MUX2_X1 cell_862_Ins_0_U1 ( .A(signal_1872), .B(signal_878), .S(n333), .Z(
        signal_877) );
  MUX2_X1 cell_862_Ins_1_U1 ( .A(signal_2912), .B(signal_3319), .S(n333), .Z(
        signal_4023) );
  MUX2_X1 cell_863_Ins_0_U1 ( .A(signal_1880), .B(signal_1816), .S(n314), .Z(
        signal_878) );
  MUX2_X1 cell_863_Ins_1_U1 ( .A(signal_2937), .B(signal_3008), .S(n314), .Z(
        signal_3319) );
  MUX2_X1 cell_866_Ins_0_U1 ( .A(signal_1871), .B(signal_881), .S(n332), .Z(
        signal_880) );
  MUX2_X1 cell_866_Ins_1_U1 ( .A(signal_2915), .B(signal_3320), .S(n332), .Z(
        signal_4024) );
  MUX2_X1 cell_867_Ins_0_U1 ( .A(signal_1879), .B(signal_1815), .S(n314), .Z(
        signal_881) );
  MUX2_X1 cell_867_Ins_1_U1 ( .A(signal_2940), .B(signal_3011), .S(n314), .Z(
        signal_3320) );
  MUX2_X1 cell_870_Ins_0_U1 ( .A(signal_1870), .B(signal_884), .S(n332), .Z(
        signal_883) );
  MUX2_X1 cell_870_Ins_1_U1 ( .A(signal_2918), .B(signal_3321), .S(n332), .Z(
        signal_4025) );
  MUX2_X1 cell_871_Ins_0_U1 ( .A(signal_1878), .B(signal_1814), .S(n315), .Z(
        signal_884) );
  MUX2_X1 cell_871_Ins_1_U1 ( .A(signal_2943), .B(signal_3014), .S(n315), .Z(
        signal_3321) );
  MUX2_X1 cell_874_Ins_0_U1 ( .A(signal_1861), .B(signal_887), .S(n332), .Z(
        signal_886) );
  MUX2_X1 cell_874_Ins_1_U1 ( .A(signal_2921), .B(signal_3322), .S(n332), .Z(
        signal_4026) );
  MUX2_X1 cell_875_Ins_0_U1 ( .A(signal_1869), .B(signal_1805), .S(n315), .Z(
        signal_887) );
  MUX2_X1 cell_875_Ins_1_U1 ( .A(signal_2946), .B(signal_3017), .S(n315), .Z(
        signal_3322) );
  MUX2_X1 cell_878_Ins_0_U1 ( .A(signal_1860), .B(signal_890), .S(n332), .Z(
        signal_889) );
  MUX2_X1 cell_878_Ins_1_U1 ( .A(signal_2924), .B(signal_3323), .S(n332), .Z(
        signal_4027) );
  MUX2_X1 cell_879_Ins_0_U1 ( .A(signal_1868), .B(signal_1804), .S(n315), .Z(
        signal_890) );
  MUX2_X1 cell_879_Ins_1_U1 ( .A(signal_2949), .B(signal_3020), .S(n315), .Z(
        signal_3323) );
  MUX2_X1 cell_882_Ins_0_U1 ( .A(signal_1859), .B(signal_893), .S(n332), .Z(
        signal_892) );
  MUX2_X1 cell_882_Ins_1_U1 ( .A(signal_2927), .B(signal_3324), .S(n332), .Z(
        signal_4028) );
  MUX2_X1 cell_883_Ins_0_U1 ( .A(signal_1867), .B(signal_1803), .S(n315), .Z(
        signal_893) );
  MUX2_X1 cell_883_Ins_1_U1 ( .A(signal_2952), .B(signal_3023), .S(n315), .Z(
        signal_3324) );
  MUX2_X1 cell_886_Ins_0_U1 ( .A(signal_1858), .B(signal_896), .S(n332), .Z(
        signal_895) );
  MUX2_X1 cell_886_Ins_1_U1 ( .A(signal_2930), .B(signal_3325), .S(n332), .Z(
        signal_4029) );
  MUX2_X1 cell_887_Ins_0_U1 ( .A(signal_1866), .B(signal_1802), .S(n315), .Z(
        signal_896) );
  MUX2_X1 cell_887_Ins_1_U1 ( .A(signal_2955), .B(signal_3026), .S(n315), .Z(
        signal_3325) );
  MUX2_X1 cell_890_Ins_0_U1 ( .A(signal_1857), .B(signal_899), .S(n332), .Z(
        signal_898) );
  MUX2_X1 cell_890_Ins_1_U1 ( .A(signal_2933), .B(signal_3326), .S(n332), .Z(
        signal_4030) );
  MUX2_X1 cell_891_Ins_0_U1 ( .A(signal_1865), .B(signal_1801), .S(n315), .Z(
        signal_899) );
  MUX2_X1 cell_891_Ins_1_U1 ( .A(signal_2958), .B(signal_3029), .S(n315), .Z(
        signal_3326) );
  MUX2_X1 cell_894_Ins_0_U1 ( .A(signal_1856), .B(signal_902), .S(n331), .Z(
        signal_901) );
  MUX2_X1 cell_894_Ins_1_U1 ( .A(signal_2936), .B(signal_3327), .S(n331), .Z(
        signal_4031) );
  MUX2_X1 cell_895_Ins_0_U1 ( .A(signal_1864), .B(signal_1800), .S(n315), .Z(
        signal_902) );
  MUX2_X1 cell_895_Ins_1_U1 ( .A(signal_2961), .B(signal_3032), .S(n315), .Z(
        signal_3327) );
  MUX2_X1 cell_898_Ins_0_U1 ( .A(signal_1855), .B(signal_905), .S(n331), .Z(
        signal_904) );
  MUX2_X1 cell_898_Ins_1_U1 ( .A(signal_2939), .B(signal_3328), .S(n331), .Z(
        signal_4032) );
  MUX2_X1 cell_899_Ins_0_U1 ( .A(signal_1863), .B(signal_1799), .S(n316), .Z(
        signal_905) );
  MUX2_X1 cell_899_Ins_1_U1 ( .A(signal_2964), .B(signal_3035), .S(n316), .Z(
        signal_3328) );
  MUX2_X1 cell_902_Ins_0_U1 ( .A(signal_1854), .B(signal_908), .S(n331), .Z(
        signal_907) );
  MUX2_X1 cell_902_Ins_1_U1 ( .A(signal_2942), .B(signal_3329), .S(n331), .Z(
        signal_4033) );
  MUX2_X1 cell_903_Ins_0_U1 ( .A(signal_1862), .B(signal_1798), .S(n316), .Z(
        signal_908) );
  MUX2_X1 cell_903_Ins_1_U1 ( .A(signal_2967), .B(signal_3038), .S(n316), .Z(
        signal_3329) );
  MUX2_X1 cell_906_Ins_0_U1 ( .A(signal_1845), .B(signal_911), .S(n331), .Z(
        signal_910) );
  MUX2_X1 cell_906_Ins_1_U1 ( .A(signal_2945), .B(signal_3330), .S(n331), .Z(
        signal_3639) );
  MUX2_X1 cell_907_Ins_0_U1 ( .A(signal_1853), .B(signal_1789), .S(n316), .Z(
        signal_911) );
  MUX2_X1 cell_907_Ins_1_U1 ( .A(signal_2970), .B(signal_3041), .S(n316), .Z(
        signal_3330) );
  MUX2_X1 cell_910_Ins_0_U1 ( .A(signal_1844), .B(signal_914), .S(n331), .Z(
        signal_913) );
  MUX2_X1 cell_910_Ins_1_U1 ( .A(signal_2948), .B(signal_3331), .S(n331), .Z(
        signal_3640) );
  MUX2_X1 cell_911_Ins_0_U1 ( .A(signal_1852), .B(signal_1788), .S(n316), .Z(
        signal_914) );
  MUX2_X1 cell_911_Ins_1_U1 ( .A(signal_2973), .B(signal_3044), .S(n316), .Z(
        signal_3331) );
  MUX2_X1 cell_914_Ins_0_U1 ( .A(signal_1843), .B(signal_917), .S(n331), .Z(
        signal_916) );
  MUX2_X1 cell_914_Ins_1_U1 ( .A(signal_2951), .B(signal_3332), .S(n331), .Z(
        signal_3641) );
  MUX2_X1 cell_915_Ins_0_U1 ( .A(signal_1851), .B(signal_1787), .S(n316), .Z(
        signal_917) );
  MUX2_X1 cell_915_Ins_1_U1 ( .A(signal_2976), .B(signal_3047), .S(n316), .Z(
        signal_3332) );
  MUX2_X1 cell_918_Ins_0_U1 ( .A(signal_1842), .B(signal_920), .S(n331), .Z(
        signal_919) );
  MUX2_X1 cell_918_Ins_1_U1 ( .A(signal_2954), .B(signal_3333), .S(n331), .Z(
        signal_3642) );
  MUX2_X1 cell_919_Ins_0_U1 ( .A(signal_1850), .B(signal_1786), .S(n316), .Z(
        signal_920) );
  MUX2_X1 cell_919_Ins_1_U1 ( .A(signal_2979), .B(signal_3050), .S(n316), .Z(
        signal_3333) );
  MUX2_X1 cell_922_Ins_0_U1 ( .A(signal_1841), .B(signal_923), .S(n337), .Z(
        signal_922) );
  MUX2_X1 cell_922_Ins_1_U1 ( .A(signal_2957), .B(signal_3334), .S(n337), .Z(
        signal_3643) );
  MUX2_X1 cell_923_Ins_0_U1 ( .A(signal_1849), .B(signal_1785), .S(n316), .Z(
        signal_923) );
  MUX2_X1 cell_923_Ins_1_U1 ( .A(signal_2982), .B(signal_3053), .S(n316), .Z(
        signal_3334) );
  MUX2_X1 cell_926_Ins_0_U1 ( .A(signal_1840), .B(signal_926), .S(n328), .Z(
        signal_925) );
  MUX2_X1 cell_926_Ins_1_U1 ( .A(signal_2960), .B(signal_3335), .S(n328), .Z(
        signal_3644) );
  MUX2_X1 cell_927_Ins_0_U1 ( .A(signal_1848), .B(signal_1784), .S(n317), .Z(
        signal_926) );
  MUX2_X1 cell_927_Ins_1_U1 ( .A(signal_2985), .B(signal_3056), .S(n317), .Z(
        signal_3335) );
  MUX2_X1 cell_930_Ins_0_U1 ( .A(signal_1839), .B(signal_929), .S(n336), .Z(
        signal_928) );
  MUX2_X1 cell_930_Ins_1_U1 ( .A(signal_2963), .B(signal_3336), .S(n336), .Z(
        signal_3645) );
  MUX2_X1 cell_931_Ins_0_U1 ( .A(signal_1847), .B(signal_1783), .S(n317), .Z(
        signal_929) );
  MUX2_X1 cell_931_Ins_1_U1 ( .A(signal_2988), .B(signal_3059), .S(n317), .Z(
        signal_3336) );
  MUX2_X1 cell_934_Ins_0_U1 ( .A(signal_1838), .B(signal_932), .S(n331), .Z(
        signal_931) );
  MUX2_X1 cell_934_Ins_1_U1 ( .A(signal_2966), .B(signal_3337), .S(n331), .Z(
        signal_3646) );
  MUX2_X1 cell_935_Ins_0_U1 ( .A(signal_1846), .B(signal_1782), .S(n317), .Z(
        signal_932) );
  MUX2_X1 cell_935_Ins_1_U1 ( .A(signal_2991), .B(signal_3062), .S(n317), .Z(
        signal_3337) );
  MUX2_X1 cell_938_Ins_0_U1 ( .A(signal_1509), .B(signal_935), .S(n327), .Z(
        signal_934) );
  MUX2_X1 cell_938_Ins_1_U1 ( .A(signal_2969), .B(signal_3338), .S(n327), .Z(
        signal_3647) );
  MUX2_X1 cell_939_Ins_0_U1 ( .A(signal_1837), .B(signal_1773), .S(n317), .Z(
        signal_935) );
  MUX2_X1 cell_939_Ins_1_U1 ( .A(signal_2994), .B(signal_3065), .S(n317), .Z(
        signal_3338) );
  MUX2_X1 cell_942_Ins_0_U1 ( .A(signal_1508), .B(signal_938), .S(n334), .Z(
        signal_937) );
  MUX2_X1 cell_942_Ins_1_U1 ( .A(signal_2972), .B(signal_3339), .S(n334), .Z(
        signal_3648) );
  MUX2_X1 cell_943_Ins_0_U1 ( .A(signal_1836), .B(signal_1772), .S(n317), .Z(
        signal_938) );
  MUX2_X1 cell_943_Ins_1_U1 ( .A(signal_2997), .B(signal_3068), .S(n317), .Z(
        signal_3339) );
  MUX2_X1 cell_946_Ins_0_U1 ( .A(signal_1507), .B(signal_941), .S(n333), .Z(
        signal_940) );
  MUX2_X1 cell_946_Ins_1_U1 ( .A(signal_2975), .B(signal_3340), .S(n333), .Z(
        signal_3649) );
  MUX2_X1 cell_947_Ins_0_U1 ( .A(signal_1835), .B(signal_1771), .S(n317), .Z(
        signal_941) );
  MUX2_X1 cell_947_Ins_1_U1 ( .A(signal_3000), .B(signal_3071), .S(n317), .Z(
        signal_3340) );
  MUX2_X1 cell_950_Ins_0_U1 ( .A(signal_1506), .B(signal_944), .S(n330), .Z(
        signal_943) );
  MUX2_X1 cell_950_Ins_1_U1 ( .A(signal_2978), .B(signal_3341), .S(n330), .Z(
        signal_3650) );
  MUX2_X1 cell_951_Ins_0_U1 ( .A(signal_1834), .B(signal_1770), .S(n317), .Z(
        signal_944) );
  MUX2_X1 cell_951_Ins_1_U1 ( .A(signal_3003), .B(signal_3074), .S(n317), .Z(
        signal_3341) );
  MUX2_X1 cell_954_Ins_0_U1 ( .A(signal_1505), .B(signal_947), .S(n330), .Z(
        signal_946) );
  MUX2_X1 cell_954_Ins_1_U1 ( .A(signal_2981), .B(signal_3342), .S(n330), .Z(
        signal_3651) );
  MUX2_X1 cell_955_Ins_0_U1 ( .A(signal_1833), .B(signal_1769), .S(n318), .Z(
        signal_947) );
  MUX2_X1 cell_955_Ins_1_U1 ( .A(signal_3006), .B(signal_3077), .S(n318), .Z(
        signal_3342) );
  MUX2_X1 cell_958_Ins_0_U1 ( .A(signal_1504), .B(signal_950), .S(n330), .Z(
        signal_949) );
  MUX2_X1 cell_958_Ins_1_U1 ( .A(signal_2984), .B(signal_3343), .S(n330), .Z(
        signal_3652) );
  MUX2_X1 cell_959_Ins_0_U1 ( .A(signal_1832), .B(signal_1768), .S(n318), .Z(
        signal_950) );
  MUX2_X1 cell_959_Ins_1_U1 ( .A(signal_3009), .B(signal_3080), .S(n318), .Z(
        signal_3343) );
  MUX2_X1 cell_962_Ins_0_U1 ( .A(signal_1503), .B(signal_953), .S(n330), .Z(
        signal_952) );
  MUX2_X1 cell_962_Ins_1_U1 ( .A(signal_2987), .B(signal_3344), .S(n330), .Z(
        signal_3653) );
  MUX2_X1 cell_963_Ins_0_U1 ( .A(signal_1831), .B(signal_1767), .S(n318), .Z(
        signal_953) );
  MUX2_X1 cell_963_Ins_1_U1 ( .A(signal_3012), .B(signal_3083), .S(n318), .Z(
        signal_3344) );
  MUX2_X1 cell_966_Ins_0_U1 ( .A(signal_1502), .B(signal_956), .S(n330), .Z(
        signal_955) );
  MUX2_X1 cell_966_Ins_1_U1 ( .A(signal_2990), .B(signal_3345), .S(n330), .Z(
        signal_3654) );
  MUX2_X1 cell_967_Ins_0_U1 ( .A(signal_1830), .B(signal_1766), .S(n318), .Z(
        signal_956) );
  MUX2_X1 cell_967_Ins_1_U1 ( .A(signal_3015), .B(signal_3086), .S(n318), .Z(
        signal_3345) );
  MUX2_X1 cell_970_Ins_0_U1 ( .A(signal_1821), .B(signal_959), .S(n330), .Z(
        signal_958) );
  MUX2_X1 cell_970_Ins_1_U1 ( .A(signal_2993), .B(signal_3346), .S(n330), .Z(
        signal_4034) );
  MUX2_X1 cell_971_Ins_0_U1 ( .A(signal_1829), .B(signal_1749), .S(n318), .Z(
        signal_959) );
  MUX2_X1 cell_971_Ins_1_U1 ( .A(signal_3018), .B(signal_3089), .S(n318), .Z(
        signal_3346) );
  MUX2_X1 cell_974_Ins_0_U1 ( .A(signal_1820), .B(signal_962), .S(n329), .Z(
        signal_961) );
  MUX2_X1 cell_974_Ins_1_U1 ( .A(signal_2996), .B(signal_3347), .S(n329), .Z(
        signal_4035) );
  MUX2_X1 cell_975_Ins_0_U1 ( .A(signal_1828), .B(signal_1748), .S(n318), .Z(
        signal_962) );
  MUX2_X1 cell_975_Ins_1_U1 ( .A(signal_3021), .B(signal_3092), .S(n318), .Z(
        signal_3347) );
  MUX2_X1 cell_978_Ins_0_U1 ( .A(signal_1819), .B(signal_965), .S(n329), .Z(
        signal_964) );
  MUX2_X1 cell_978_Ins_1_U1 ( .A(signal_2999), .B(signal_3348), .S(n329), .Z(
        signal_4036) );
  MUX2_X1 cell_979_Ins_0_U1 ( .A(signal_1827), .B(signal_1747), .S(n318), .Z(
        signal_965) );
  MUX2_X1 cell_979_Ins_1_U1 ( .A(signal_3024), .B(signal_3095), .S(n318), .Z(
        signal_3348) );
  MUX2_X1 cell_982_Ins_0_U1 ( .A(signal_1818), .B(signal_968), .S(n329), .Z(
        signal_967) );
  MUX2_X1 cell_982_Ins_1_U1 ( .A(signal_3002), .B(signal_3349), .S(n329), .Z(
        signal_4037) );
  MUX2_X1 cell_983_Ins_0_U1 ( .A(signal_1826), .B(signal_1746), .S(n319), .Z(
        signal_968) );
  MUX2_X1 cell_983_Ins_1_U1 ( .A(signal_3027), .B(signal_3098), .S(n319), .Z(
        signal_3349) );
  MUX2_X1 cell_986_Ins_0_U1 ( .A(signal_1817), .B(signal_971), .S(n329), .Z(
        signal_970) );
  MUX2_X1 cell_986_Ins_1_U1 ( .A(signal_3005), .B(signal_3350), .S(n329), .Z(
        signal_4038) );
  MUX2_X1 cell_987_Ins_0_U1 ( .A(signal_1825), .B(signal_1745), .S(n319), .Z(
        signal_971) );
  MUX2_X1 cell_987_Ins_1_U1 ( .A(signal_3030), .B(signal_3101), .S(n319), .Z(
        signal_3350) );
  MUX2_X1 cell_990_Ins_0_U1 ( .A(signal_1816), .B(signal_974), .S(n329), .Z(
        signal_973) );
  MUX2_X1 cell_990_Ins_1_U1 ( .A(signal_3008), .B(signal_3351), .S(n329), .Z(
        signal_4039) );
  MUX2_X1 cell_991_Ins_0_U1 ( .A(signal_1824), .B(signal_1744), .S(n319), .Z(
        signal_974) );
  MUX2_X1 cell_991_Ins_1_U1 ( .A(signal_3033), .B(signal_3104), .S(n319), .Z(
        signal_3351) );
  MUX2_X1 cell_994_Ins_0_U1 ( .A(signal_1815), .B(signal_977), .S(n329), .Z(
        signal_976) );
  MUX2_X1 cell_994_Ins_1_U1 ( .A(signal_3011), .B(signal_3352), .S(n329), .Z(
        signal_4040) );
  MUX2_X1 cell_995_Ins_0_U1 ( .A(signal_1823), .B(signal_1743), .S(n319), .Z(
        signal_977) );
  MUX2_X1 cell_995_Ins_1_U1 ( .A(signal_3036), .B(signal_3107), .S(n319), .Z(
        signal_3352) );
  MUX2_X1 cell_998_Ins_0_U1 ( .A(signal_1814), .B(signal_980), .S(n329), .Z(
        signal_979) );
  MUX2_X1 cell_998_Ins_1_U1 ( .A(signal_3014), .B(signal_3353), .S(n329), .Z(
        signal_4041) );
  MUX2_X1 cell_999_Ins_0_U1 ( .A(signal_1822), .B(signal_1742), .S(n319), .Z(
        signal_980) );
  MUX2_X1 cell_999_Ins_1_U1 ( .A(signal_3039), .B(signal_3110), .S(n319), .Z(
        signal_3353) );
  MUX2_X1 cell_1002_Ins_0_U1 ( .A(signal_1805), .B(signal_983), .S(n328), .Z(
        signal_982) );
  MUX2_X1 cell_1002_Ins_1_U1 ( .A(signal_3017), .B(signal_3354), .S(n328), .Z(
        signal_4042) );
  MUX2_X1 cell_1003_Ins_0_U1 ( .A(signal_1813), .B(signal_1733), .S(n319), .Z(
        signal_983) );
  MUX2_X1 cell_1003_Ins_1_U1 ( .A(signal_3042), .B(signal_3113), .S(n319), .Z(
        signal_3354) );
  MUX2_X1 cell_1006_Ins_0_U1 ( .A(signal_1804), .B(signal_986), .S(n328), .Z(
        signal_985) );
  MUX2_X1 cell_1006_Ins_1_U1 ( .A(signal_3020), .B(signal_3355), .S(n328), .Z(
        signal_4043) );
  MUX2_X1 cell_1007_Ins_0_U1 ( .A(signal_1812), .B(signal_1732), .S(n319), .Z(
        signal_986) );
  MUX2_X1 cell_1007_Ins_1_U1 ( .A(signal_3045), .B(signal_3116), .S(n319), .Z(
        signal_3355) );
  MUX2_X1 cell_1010_Ins_0_U1 ( .A(signal_1803), .B(signal_989), .S(n328), .Z(
        signal_988) );
  MUX2_X1 cell_1010_Ins_1_U1 ( .A(signal_3023), .B(signal_3356), .S(n328), .Z(
        signal_4044) );
  MUX2_X1 cell_1011_Ins_0_U1 ( .A(signal_1811), .B(signal_1731), .S(n320), .Z(
        signal_989) );
  MUX2_X1 cell_1011_Ins_1_U1 ( .A(signal_3048), .B(signal_3119), .S(n320), .Z(
        signal_3356) );
  MUX2_X1 cell_1014_Ins_0_U1 ( .A(signal_1802), .B(signal_992), .S(n328), .Z(
        signal_991) );
  MUX2_X1 cell_1014_Ins_1_U1 ( .A(signal_3026), .B(signal_3357), .S(n328), .Z(
        signal_4045) );
  MUX2_X1 cell_1015_Ins_0_U1 ( .A(signal_1810), .B(signal_1730), .S(n320), .Z(
        signal_992) );
  MUX2_X1 cell_1015_Ins_1_U1 ( .A(signal_3051), .B(signal_3122), .S(n320), .Z(
        signal_3357) );
  MUX2_X1 cell_1018_Ins_0_U1 ( .A(signal_1801), .B(signal_995), .S(n328), .Z(
        signal_994) );
  MUX2_X1 cell_1018_Ins_1_U1 ( .A(signal_3029), .B(signal_3358), .S(n328), .Z(
        signal_4046) );
  MUX2_X1 cell_1019_Ins_0_U1 ( .A(signal_1809), .B(signal_1729), .S(n320), .Z(
        signal_995) );
  MUX2_X1 cell_1019_Ins_1_U1 ( .A(signal_3054), .B(signal_3125), .S(n320), .Z(
        signal_3358) );
  MUX2_X1 cell_1022_Ins_0_U1 ( .A(signal_1800), .B(signal_998), .S(n328), .Z(
        signal_997) );
  MUX2_X1 cell_1022_Ins_1_U1 ( .A(signal_3032), .B(signal_3359), .S(n328), .Z(
        signal_4047) );
  MUX2_X1 cell_1023_Ins_0_U1 ( .A(signal_1808), .B(signal_1728), .S(n320), .Z(
        signal_998) );
  MUX2_X1 cell_1023_Ins_1_U1 ( .A(signal_3057), .B(signal_3128), .S(n320), .Z(
        signal_3359) );
  MUX2_X1 cell_1026_Ins_0_U1 ( .A(signal_1799), .B(signal_1001), .S(n328), .Z(
        signal_1000) );
  MUX2_X1 cell_1026_Ins_1_U1 ( .A(signal_3035), .B(signal_3360), .S(n328), .Z(
        signal_4048) );
  MUX2_X1 cell_1027_Ins_0_U1 ( .A(signal_1807), .B(signal_1727), .S(n320), .Z(
        signal_1001) );
  MUX2_X1 cell_1027_Ins_1_U1 ( .A(signal_3060), .B(signal_3131), .S(n320), .Z(
        signal_3360) );
  MUX2_X1 cell_1030_Ins_0_U1 ( .A(signal_1798), .B(signal_1004), .S(n327), .Z(
        signal_1003) );
  MUX2_X1 cell_1030_Ins_1_U1 ( .A(signal_3038), .B(signal_3361), .S(n327), .Z(
        signal_4049) );
  MUX2_X1 cell_1031_Ins_0_U1 ( .A(signal_1806), .B(signal_1726), .S(n320), .Z(
        signal_1004) );
  MUX2_X1 cell_1031_Ins_1_U1 ( .A(signal_3063), .B(signal_3134), .S(n320), .Z(
        signal_3361) );
  MUX2_X1 cell_1034_Ins_0_U1 ( .A(signal_1789), .B(signal_1007), .S(n327), .Z(
        signal_1006) );
  MUX2_X1 cell_1034_Ins_1_U1 ( .A(signal_3041), .B(signal_3362), .S(n327), .Z(
        signal_4050) );
  MUX2_X1 cell_1035_Ins_0_U1 ( .A(signal_1797), .B(signal_1717), .S(n320), .Z(
        signal_1007) );
  MUX2_X1 cell_1035_Ins_1_U1 ( .A(signal_3066), .B(signal_3137), .S(n320), .Z(
        signal_3362) );
  MUX2_X1 cell_1038_Ins_0_U1 ( .A(signal_1788), .B(signal_1010), .S(n327), .Z(
        signal_1009) );
  MUX2_X1 cell_1038_Ins_1_U1 ( .A(signal_3044), .B(signal_3363), .S(n327), .Z(
        signal_4051) );
  MUX2_X1 cell_1039_Ins_0_U1 ( .A(signal_1796), .B(signal_1716), .S(n321), .Z(
        signal_1010) );
  MUX2_X1 cell_1039_Ins_1_U1 ( .A(signal_3069), .B(signal_3140), .S(n321), .Z(
        signal_3363) );
  MUX2_X1 cell_1042_Ins_0_U1 ( .A(signal_1787), .B(signal_1013), .S(n327), .Z(
        signal_1012) );
  MUX2_X1 cell_1042_Ins_1_U1 ( .A(signal_3047), .B(signal_3364), .S(n327), .Z(
        signal_4052) );
  MUX2_X1 cell_1043_Ins_0_U1 ( .A(signal_1795), .B(signal_1715), .S(n321), .Z(
        signal_1013) );
  MUX2_X1 cell_1043_Ins_1_U1 ( .A(signal_3072), .B(signal_3143), .S(n321), .Z(
        signal_3364) );
  MUX2_X1 cell_1046_Ins_0_U1 ( .A(signal_1786), .B(signal_1016), .S(n327), .Z(
        signal_1015) );
  MUX2_X1 cell_1046_Ins_1_U1 ( .A(signal_3050), .B(signal_3365), .S(n327), .Z(
        signal_4053) );
  MUX2_X1 cell_1047_Ins_0_U1 ( .A(signal_1794), .B(signal_1714), .S(n321), .Z(
        signal_1016) );
  MUX2_X1 cell_1047_Ins_1_U1 ( .A(signal_3075), .B(signal_3146), .S(n321), .Z(
        signal_3365) );
  MUX2_X1 cell_1050_Ins_0_U1 ( .A(signal_1785), .B(signal_1019), .S(n327), .Z(
        signal_1018) );
  MUX2_X1 cell_1050_Ins_1_U1 ( .A(signal_3053), .B(signal_3366), .S(n327), .Z(
        signal_4054) );
  MUX2_X1 cell_1051_Ins_0_U1 ( .A(signal_1793), .B(signal_1713), .S(n321), .Z(
        signal_1019) );
  MUX2_X1 cell_1051_Ins_1_U1 ( .A(signal_3078), .B(signal_3149), .S(n321), .Z(
        signal_3366) );
  MUX2_X1 cell_1054_Ins_0_U1 ( .A(signal_1784), .B(signal_1022), .S(n327), .Z(
        signal_1021) );
  MUX2_X1 cell_1054_Ins_1_U1 ( .A(signal_3056), .B(signal_3367), .S(n327), .Z(
        signal_4055) );
  MUX2_X1 cell_1055_Ins_0_U1 ( .A(signal_1792), .B(signal_1712), .S(n321), .Z(
        signal_1022) );
  MUX2_X1 cell_1055_Ins_1_U1 ( .A(signal_3081), .B(signal_3152), .S(n321), .Z(
        signal_3367) );
  MUX2_X1 cell_1058_Ins_0_U1 ( .A(signal_1783), .B(signal_1025), .S(n334), .Z(
        signal_1024) );
  MUX2_X1 cell_1058_Ins_1_U1 ( .A(signal_3059), .B(signal_3368), .S(n334), .Z(
        signal_4056) );
  MUX2_X1 cell_1059_Ins_0_U1 ( .A(signal_1791), .B(signal_1711), .S(n321), .Z(
        signal_1025) );
  MUX2_X1 cell_1059_Ins_1_U1 ( .A(signal_3084), .B(signal_3155), .S(n321), .Z(
        signal_3368) );
  MUX2_X1 cell_1062_Ins_0_U1 ( .A(signal_1782), .B(signal_1028), .S(n324), .Z(
        signal_1027) );
  MUX2_X1 cell_1062_Ins_1_U1 ( .A(signal_3062), .B(signal_3369), .S(n324), .Z(
        signal_4057) );
  MUX2_X1 cell_1063_Ins_0_U1 ( .A(signal_1790), .B(signal_1710), .S(n321), .Z(
        signal_1028) );
  MUX2_X1 cell_1063_Ins_1_U1 ( .A(signal_3087), .B(signal_3158), .S(n321), .Z(
        signal_3369) );
  MUX2_X1 cell_1066_Ins_0_U1 ( .A(signal_1773), .B(signal_1031), .S(n331), .Z(
        signal_1030) );
  MUX2_X1 cell_1066_Ins_1_U1 ( .A(signal_3065), .B(signal_3370), .S(n331), .Z(
        signal_4058) );
  MUX2_X1 cell_1067_Ins_0_U1 ( .A(signal_1781), .B(signal_1701), .S(n322), .Z(
        signal_1031) );
  MUX2_X1 cell_1067_Ins_1_U1 ( .A(signal_3090), .B(signal_3161), .S(n322), .Z(
        signal_3370) );
  MUX2_X1 cell_1070_Ins_0_U1 ( .A(signal_1772), .B(signal_1034), .S(n327), .Z(
        signal_1033) );
  MUX2_X1 cell_1070_Ins_1_U1 ( .A(signal_3068), .B(signal_3371), .S(n327), .Z(
        signal_4059) );
  MUX2_X1 cell_1071_Ins_0_U1 ( .A(signal_1780), .B(signal_1700), .S(n322), .Z(
        signal_1034) );
  MUX2_X1 cell_1071_Ins_1_U1 ( .A(signal_3093), .B(signal_3164), .S(n322), .Z(
        signal_3371) );
  MUX2_X1 cell_1074_Ins_0_U1 ( .A(signal_1771), .B(signal_1037), .S(n334), .Z(
        signal_1036) );
  MUX2_X1 cell_1074_Ins_1_U1 ( .A(signal_3071), .B(signal_3372), .S(n334), .Z(
        signal_4060) );
  MUX2_X1 cell_1075_Ins_0_U1 ( .A(signal_1779), .B(signal_1699), .S(n322), .Z(
        signal_1037) );
  MUX2_X1 cell_1075_Ins_1_U1 ( .A(signal_3096), .B(signal_3167), .S(n322), .Z(
        signal_3372) );
  MUX2_X1 cell_1078_Ins_0_U1 ( .A(signal_1770), .B(signal_1040), .S(n329), .Z(
        signal_1039) );
  MUX2_X1 cell_1078_Ins_1_U1 ( .A(signal_3074), .B(signal_3373), .S(n329), .Z(
        signal_4061) );
  MUX2_X1 cell_1079_Ins_0_U1 ( .A(signal_1778), .B(signal_1698), .S(n322), .Z(
        signal_1040) );
  MUX2_X1 cell_1079_Ins_1_U1 ( .A(signal_3099), .B(signal_3170), .S(n322), .Z(
        signal_3373) );
  MUX2_X1 cell_1082_Ins_0_U1 ( .A(signal_1769), .B(signal_1043), .S(n335), .Z(
        signal_1042) );
  MUX2_X1 cell_1082_Ins_1_U1 ( .A(signal_3077), .B(signal_3374), .S(n335), .Z(
        signal_4062) );
  MUX2_X1 cell_1083_Ins_0_U1 ( .A(signal_1777), .B(signal_1697), .S(n322), .Z(
        signal_1043) );
  MUX2_X1 cell_1083_Ins_1_U1 ( .A(signal_3102), .B(signal_3173), .S(n322), .Z(
        signal_3374) );
  MUX2_X1 cell_1086_Ins_0_U1 ( .A(signal_1768), .B(signal_1046), .S(n326), .Z(
        signal_1045) );
  MUX2_X1 cell_1086_Ins_1_U1 ( .A(signal_3080), .B(signal_3375), .S(n326), .Z(
        signal_4063) );
  MUX2_X1 cell_1087_Ins_0_U1 ( .A(signal_1776), .B(signal_1696), .S(n322), .Z(
        signal_1046) );
  MUX2_X1 cell_1087_Ins_1_U1 ( .A(signal_3105), .B(signal_3176), .S(n322), .Z(
        signal_3375) );
  MUX2_X1 cell_1090_Ins_0_U1 ( .A(signal_1767), .B(signal_1049), .S(n326), .Z(
        signal_1048) );
  MUX2_X1 cell_1090_Ins_1_U1 ( .A(signal_3083), .B(signal_3376), .S(n326), .Z(
        signal_4064) );
  MUX2_X1 cell_1091_Ins_0_U1 ( .A(signal_1775), .B(signal_1695), .S(n322), .Z(
        signal_1049) );
  MUX2_X1 cell_1091_Ins_1_U1 ( .A(signal_3108), .B(signal_3179), .S(n322), .Z(
        signal_3376) );
  MUX2_X1 cell_1094_Ins_0_U1 ( .A(signal_1766), .B(signal_1052), .S(n326), .Z(
        signal_1051) );
  MUX2_X1 cell_1094_Ins_1_U1 ( .A(signal_3086), .B(signal_3377), .S(n326), .Z(
        signal_4065) );
  MUX2_X1 cell_1095_Ins_0_U1 ( .A(signal_1774), .B(signal_1694), .S(n323), .Z(
        signal_1052) );
  MUX2_X1 cell_1095_Ins_1_U1 ( .A(signal_3111), .B(signal_3182), .S(n323), .Z(
        signal_3377) );
  MUX2_X1 cell_1130_Ins_0_U1 ( .A(signal_1733), .B(signal_1079), .S(n326), .Z(
        signal_1078) );
  MUX2_X1 cell_1130_Ins_1_U1 ( .A(signal_3113), .B(signal_3378), .S(n326), .Z(
        signal_4066) );
  MUX2_X1 cell_1131_Ins_0_U1 ( .A(signal_1741), .B(signal_758), .S(n323), .Z(
        signal_1079) );
  MUX2_X1 cell_1131_Ins_1_U1 ( .A(signal_3138), .B(signal_2426), .S(n323), .Z(
        signal_3378) );
  MUX2_X1 cell_1134_Ins_0_U1 ( .A(signal_1732), .B(signal_1082), .S(n326), .Z(
        signal_1081) );
  MUX2_X1 cell_1134_Ins_1_U1 ( .A(signal_3116), .B(signal_3379), .S(n326), .Z(
        signal_4067) );
  MUX2_X1 cell_1135_Ins_0_U1 ( .A(signal_1740), .B(signal_759), .S(n323), .Z(
        signal_1082) );
  MUX2_X1 cell_1135_Ins_1_U1 ( .A(signal_3141), .B(signal_2424), .S(n323), .Z(
        signal_3379) );
  MUX2_X1 cell_1138_Ins_0_U1 ( .A(signal_1731), .B(signal_1085), .S(n326), .Z(
        signal_1084) );
  MUX2_X1 cell_1138_Ins_1_U1 ( .A(signal_3119), .B(signal_3380), .S(n326), .Z(
        signal_4068) );
  MUX2_X1 cell_1139_Ins_0_U1 ( .A(signal_1739), .B(signal_760), .S(n323), .Z(
        signal_1085) );
  MUX2_X1 cell_1139_Ins_1_U1 ( .A(signal_3144), .B(signal_2422), .S(n323), .Z(
        signal_3380) );
  MUX2_X1 cell_1142_Ins_0_U1 ( .A(signal_1730), .B(signal_1088), .S(n326), .Z(
        signal_1087) );
  MUX2_X1 cell_1142_Ins_1_U1 ( .A(signal_3122), .B(signal_3381), .S(n326), .Z(
        signal_4069) );
  MUX2_X1 cell_1143_Ins_0_U1 ( .A(signal_1738), .B(signal_761), .S(n323), .Z(
        signal_1088) );
  MUX2_X1 cell_1143_Ins_1_U1 ( .A(signal_3147), .B(signal_2420), .S(n323), .Z(
        signal_3381) );
  MUX2_X1 cell_1146_Ins_0_U1 ( .A(signal_1729), .B(signal_1091), .S(n325), .Z(
        signal_1090) );
  MUX2_X1 cell_1146_Ins_1_U1 ( .A(signal_3125), .B(signal_3382), .S(n325), .Z(
        signal_4070) );
  MUX2_X1 cell_1147_Ins_0_U1 ( .A(signal_1737), .B(signal_762), .S(n323), .Z(
        signal_1091) );
  MUX2_X1 cell_1147_Ins_1_U1 ( .A(signal_3150), .B(signal_2418), .S(n323), .Z(
        signal_3382) );
  MUX2_X1 cell_1150_Ins_0_U1 ( .A(signal_1728), .B(signal_1094), .S(n330), .Z(
        signal_1093) );
  MUX2_X1 cell_1150_Ins_1_U1 ( .A(signal_3128), .B(signal_3383), .S(n330), .Z(
        signal_4071) );
  MUX2_X1 cell_1151_Ins_0_U1 ( .A(signal_1736), .B(signal_763), .S(n323), .Z(
        signal_1094) );
  MUX2_X1 cell_1151_Ins_1_U1 ( .A(signal_3153), .B(signal_2416), .S(n323), .Z(
        signal_3383) );
  MUX2_X1 cell_1154_Ins_0_U1 ( .A(signal_1727), .B(signal_1097), .S(n325), .Z(
        signal_1096) );
  MUX2_X1 cell_1154_Ins_1_U1 ( .A(signal_3131), .B(signal_3384), .S(n325), .Z(
        signal_4072) );
  MUX2_X1 cell_1155_Ins_0_U1 ( .A(signal_1735), .B(signal_764), .S(n310), .Z(
        signal_1097) );
  MUX2_X1 cell_1155_Ins_1_U1 ( .A(signal_3156), .B(signal_2414), .S(n310), .Z(
        signal_3384) );
  MUX2_X1 cell_1158_Ins_0_U1 ( .A(signal_1726), .B(signal_1100), .S(n325), .Z(
        signal_1099) );
  MUX2_X1 cell_1158_Ins_1_U1 ( .A(signal_3134), .B(signal_3385), .S(n325), .Z(
        signal_4073) );
  MUX2_X1 cell_1159_Ins_0_U1 ( .A(signal_1734), .B(signal_765), .S(n315), .Z(
        signal_1100) );
  MUX2_X1 cell_1159_Ins_1_U1 ( .A(signal_3159), .B(signal_2412), .S(n315), .Z(
        signal_3385) );
  MUX2_X1 cell_1162_Ins_0_U1 ( .A(signal_1717), .B(signal_1103), .S(n325), .Z(
        signal_1102) );
  MUX2_X1 cell_1162_Ins_1_U1 ( .A(signal_3137), .B(signal_3386), .S(n325), .Z(
        signal_4074) );
  MUX2_X1 cell_1163_Ins_0_U1 ( .A(signal_1725), .B(signal_1909), .S(n313), .Z(
        signal_1103) );
  MUX2_X1 cell_1163_Ins_1_U1 ( .A(signal_3162), .B(signal_2849), .S(n313), .Z(
        signal_3386) );
  MUX2_X1 cell_1166_Ins_0_U1 ( .A(signal_1716), .B(signal_1106), .S(n325), .Z(
        signal_1105) );
  MUX2_X1 cell_1166_Ins_1_U1 ( .A(signal_3140), .B(signal_3387), .S(n325), .Z(
        signal_4075) );
  MUX2_X1 cell_1167_Ins_0_U1 ( .A(signal_1724), .B(signal_1908), .S(n322), .Z(
        signal_1106) );
  MUX2_X1 cell_1167_Ins_1_U1 ( .A(signal_3165), .B(signal_2852), .S(n322), .Z(
        signal_3387) );
  MUX2_X1 cell_1170_Ins_0_U1 ( .A(signal_1715), .B(signal_1109), .S(n325), .Z(
        signal_1108) );
  MUX2_X1 cell_1170_Ins_1_U1 ( .A(signal_3143), .B(signal_3388), .S(n325), .Z(
        signal_4076) );
  MUX2_X1 cell_1171_Ins_0_U1 ( .A(signal_1723), .B(signal_1907), .S(n320), .Z(
        signal_1109) );
  MUX2_X1 cell_1171_Ins_1_U1 ( .A(signal_3168), .B(signal_2855), .S(n320), .Z(
        signal_3388) );
  MUX2_X1 cell_1174_Ins_0_U1 ( .A(signal_1714), .B(signal_1112), .S(n325), .Z(
        signal_1111) );
  MUX2_X1 cell_1174_Ins_1_U1 ( .A(signal_3146), .B(signal_3389), .S(n325), .Z(
        signal_4077) );
  MUX2_X1 cell_1175_Ins_0_U1 ( .A(signal_1722), .B(signal_1906), .S(n312), .Z(
        signal_1112) );
  MUX2_X1 cell_1175_Ins_1_U1 ( .A(signal_3171), .B(signal_2858), .S(n312), .Z(
        signal_3389) );
  MUX2_X1 cell_1178_Ins_0_U1 ( .A(signal_1713), .B(signal_1115), .S(n324), .Z(
        signal_1114) );
  MUX2_X1 cell_1178_Ins_1_U1 ( .A(signal_3149), .B(signal_3390), .S(n324), .Z(
        signal_4078) );
  MUX2_X1 cell_1179_Ins_0_U1 ( .A(signal_1721), .B(signal_1905), .S(n311), .Z(
        signal_1115) );
  MUX2_X1 cell_1179_Ins_1_U1 ( .A(signal_3174), .B(signal_2861), .S(n311), .Z(
        signal_3390) );
  MUX2_X1 cell_1182_Ins_0_U1 ( .A(signal_1712), .B(signal_1118), .S(n324), .Z(
        signal_1117) );
  MUX2_X1 cell_1182_Ins_1_U1 ( .A(signal_3152), .B(signal_3391), .S(n324), .Z(
        signal_4079) );
  MUX2_X1 cell_1183_Ins_0_U1 ( .A(signal_1720), .B(signal_1904), .S(n313), .Z(
        signal_1118) );
  MUX2_X1 cell_1183_Ins_1_U1 ( .A(signal_3177), .B(signal_2864), .S(n313), .Z(
        signal_3391) );
  MUX2_X1 cell_1186_Ins_0_U1 ( .A(signal_1711), .B(signal_1121), .S(n324), .Z(
        signal_1120) );
  MUX2_X1 cell_1186_Ins_1_U1 ( .A(signal_3155), .B(signal_3392), .S(n324), .Z(
        signal_4080) );
  MUX2_X1 cell_1187_Ins_0_U1 ( .A(signal_1719), .B(signal_1903), .S(n322), .Z(
        signal_1121) );
  MUX2_X1 cell_1187_Ins_1_U1 ( .A(signal_3180), .B(signal_2867), .S(n322), .Z(
        signal_3392) );
  MUX2_X1 cell_1190_Ins_0_U1 ( .A(signal_1710), .B(signal_1124), .S(n324), .Z(
        signal_1123) );
  MUX2_X1 cell_1190_Ins_1_U1 ( .A(signal_3158), .B(signal_3393), .S(n324), .Z(
        signal_4081) );
  MUX2_X1 cell_1191_Ins_0_U1 ( .A(signal_1718), .B(signal_1902), .S(n320), .Z(
        signal_1124) );
  MUX2_X1 cell_1191_Ins_1_U1 ( .A(signal_3183), .B(signal_2870), .S(n320), .Z(
        signal_3393) );
  MUX2_X1 cell_1194_Ins_0_U1 ( .A(signal_1701), .B(signal_1127), .S(n324), .Z(
        signal_1126) );
  MUX2_X1 cell_1194_Ins_1_U1 ( .A(signal_3161), .B(signal_3394), .S(n324), .Z(
        signal_4082) );
  MUX2_X1 cell_1195_Ins_0_U1 ( .A(signal_1709), .B(signal_1893), .S(n312), .Z(
        signal_1127) );
  MUX2_X1 cell_1195_Ins_1_U1 ( .A(signal_3185), .B(signal_2873), .S(n312), .Z(
        signal_3394) );
  MUX2_X1 cell_1198_Ins_0_U1 ( .A(signal_1700), .B(signal_1130), .S(n324), .Z(
        signal_1129) );
  MUX2_X1 cell_1198_Ins_1_U1 ( .A(signal_3164), .B(signal_3395), .S(n324), .Z(
        signal_4083) );
  MUX2_X1 cell_1199_Ins_0_U1 ( .A(signal_1708), .B(signal_1892), .S(n311), .Z(
        signal_1130) );
  MUX2_X1 cell_1199_Ins_1_U1 ( .A(signal_3187), .B(signal_2876), .S(n311), .Z(
        signal_3395) );
  MUX2_X1 cell_1202_Ins_0_U1 ( .A(signal_1699), .B(signal_1133), .S(n324), .Z(
        signal_1132) );
  MUX2_X1 cell_1202_Ins_1_U1 ( .A(signal_3167), .B(signal_3396), .S(n324), .Z(
        signal_4084) );
  MUX2_X1 cell_1203_Ins_0_U1 ( .A(signal_1707), .B(signal_1891), .S(n318), .Z(
        signal_1133) );
  MUX2_X1 cell_1203_Ins_1_U1 ( .A(signal_3189), .B(signal_2879), .S(n318), .Z(
        signal_3396) );
  MUX2_X1 cell_1206_Ins_0_U1 ( .A(signal_1698), .B(signal_1136), .S(n326), .Z(
        signal_1135) );
  MUX2_X1 cell_1206_Ins_1_U1 ( .A(signal_3170), .B(signal_3397), .S(n326), .Z(
        signal_4085) );
  MUX2_X1 cell_1207_Ins_0_U1 ( .A(signal_1706), .B(signal_1890), .S(n314), .Z(
        signal_1136) );
  MUX2_X1 cell_1207_Ins_1_U1 ( .A(signal_3191), .B(signal_2882), .S(n314), .Z(
        signal_3397) );
  MUX2_X1 cell_1210_Ins_0_U1 ( .A(signal_1697), .B(signal_1139), .S(n324), .Z(
        signal_1138) );
  MUX2_X1 cell_1210_Ins_1_U1 ( .A(signal_3173), .B(signal_3398), .S(n324), .Z(
        signal_4086) );
  MUX2_X1 cell_1211_Ins_0_U1 ( .A(signal_1705), .B(signal_1889), .S(n314), .Z(
        signal_1139) );
  MUX2_X1 cell_1211_Ins_1_U1 ( .A(signal_3193), .B(signal_2885), .S(n314), .Z(
        signal_3398) );
  MUX2_X1 cell_1214_Ins_0_U1 ( .A(signal_1696), .B(signal_1142), .S(n335), .Z(
        signal_1141) );
  MUX2_X1 cell_1214_Ins_1_U1 ( .A(signal_3176), .B(signal_3399), .S(n335), .Z(
        signal_4087) );
  MUX2_X1 cell_1215_Ins_0_U1 ( .A(signal_1704), .B(signal_1888), .S(n242), .Z(
        signal_1142) );
  MUX2_X1 cell_1215_Ins_1_U1 ( .A(signal_3195), .B(signal_2888), .S(n242), .Z(
        signal_3399) );
  MUX2_X1 cell_1218_Ins_0_U1 ( .A(signal_1695), .B(signal_1145), .S(n333), .Z(
        signal_1144) );
  MUX2_X1 cell_1218_Ins_1_U1 ( .A(signal_3179), .B(signal_3400), .S(n333), .Z(
        signal_4088) );
  MUX2_X1 cell_1219_Ins_0_U1 ( .A(signal_1703), .B(signal_1887), .S(n242), .Z(
        signal_1145) );
  MUX2_X1 cell_1219_Ins_1_U1 ( .A(signal_3197), .B(signal_2891), .S(n242), .Z(
        signal_3400) );
  MUX2_X1 cell_1222_Ins_0_U1 ( .A(signal_1694), .B(signal_1148), .S(n337), .Z(
        signal_1147) );
  MUX2_X1 cell_1222_Ins_1_U1 ( .A(signal_3182), .B(signal_3401), .S(n337), .Z(
        signal_4089) );
  MUX2_X1 cell_1223_Ins_0_U1 ( .A(signal_1702), .B(signal_1886), .S(n242), .Z(
        signal_1148) );
  MUX2_X1 cell_1223_Ins_1_U1 ( .A(signal_3199), .B(signal_2894), .S(n242), .Z(
        signal_3401) );
  MUX2_X1 cell_1226_Ins_0_U1 ( .A(signal_758), .B(signal_1693), .S(signal_400), 
        .Z(signal_1685) );
  MUX2_X1 cell_1226_Ins_1_U1 ( .A(signal_2426), .B(signal_2427), .S(signal_400), .Z(signal_3655) );
  MUX2_X1 cell_1227_Ins_0_U1 ( .A(signal_759), .B(signal_1692), .S(signal_400), 
        .Z(signal_1684) );
  MUX2_X1 cell_1227_Ins_1_U1 ( .A(signal_2424), .B(signal_2425), .S(signal_400), .Z(signal_3656) );
  MUX2_X1 cell_1228_Ins_0_U1 ( .A(signal_760), .B(signal_1691), .S(signal_400), 
        .Z(signal_1683) );
  MUX2_X1 cell_1228_Ins_1_U1 ( .A(signal_2422), .B(signal_2423), .S(signal_400), .Z(signal_3657) );
  MUX2_X1 cell_1229_Ins_0_U1 ( .A(signal_761), .B(signal_1690), .S(signal_400), 
        .Z(signal_1682) );
  MUX2_X1 cell_1229_Ins_1_U1 ( .A(signal_2420), .B(signal_2421), .S(signal_400), .Z(signal_3658) );
  MUX2_X1 cell_1230_Ins_0_U1 ( .A(signal_762), .B(signal_1689), .S(signal_400), 
        .Z(signal_1681) );
  MUX2_X1 cell_1230_Ins_1_U1 ( .A(signal_2418), .B(signal_2419), .S(signal_400), .Z(signal_3659) );
  MUX2_X1 cell_1231_Ins_0_U1 ( .A(signal_763), .B(signal_1688), .S(signal_400), 
        .Z(signal_1680) );
  MUX2_X1 cell_1231_Ins_1_U1 ( .A(signal_2416), .B(signal_2417), .S(signal_400), .Z(signal_3660) );
  MUX2_X1 cell_1232_Ins_0_U1 ( .A(signal_764), .B(signal_1687), .S(signal_400), 
        .Z(signal_1679) );
  MUX2_X1 cell_1232_Ins_1_U1 ( .A(signal_2414), .B(signal_2415), .S(signal_400), .Z(signal_3661) );
  MUX2_X1 cell_1233_Ins_0_U1 ( .A(signal_765), .B(signal_1686), .S(signal_400), 
        .Z(signal_1678) );
  MUX2_X1 cell_1233_Ins_1_U1 ( .A(signal_2412), .B(signal_2413), .S(signal_400), .Z(signal_3662) );
  MUX2_X1 cell_1234_Ins_0_U1 ( .A(key_s0[120]), .B(signal_1685), .S(n281), .Z(
        signal_1933) );
  MUX2_X1 cell_1234_Ins_1_U1 ( .A(key_s1[120]), .B(signal_3655), .S(n281), .Z(
        signal_3907) );
  MUX2_X1 cell_1235_Ins_0_U1 ( .A(key_s0[121]), .B(signal_1684), .S(n282), .Z(
        signal_1932) );
  MUX2_X1 cell_1235_Ins_1_U1 ( .A(key_s1[121]), .B(signal_3656), .S(n282), .Z(
        signal_3909) );
  MUX2_X1 cell_1236_Ins_0_U1 ( .A(key_s0[122]), .B(signal_1683), .S(n284), .Z(
        signal_1931) );
  MUX2_X1 cell_1236_Ins_1_U1 ( .A(key_s1[122]), .B(signal_3657), .S(n284), .Z(
        signal_3911) );
  MUX2_X1 cell_1237_Ins_0_U1 ( .A(key_s0[123]), .B(signal_1682), .S(n283), .Z(
        signal_1930) );
  MUX2_X1 cell_1237_Ins_1_U1 ( .A(key_s1[123]), .B(signal_3658), .S(n283), .Z(
        signal_3913) );
  MUX2_X1 cell_1238_Ins_0_U1 ( .A(key_s0[124]), .B(signal_1681), .S(n285), .Z(
        signal_1929) );
  MUX2_X1 cell_1238_Ins_1_U1 ( .A(key_s1[124]), .B(signal_3659), .S(n285), .Z(
        signal_3915) );
  MUX2_X1 cell_1239_Ins_0_U1 ( .A(key_s0[125]), .B(signal_1680), .S(n286), .Z(
        signal_1928) );
  MUX2_X1 cell_1239_Ins_1_U1 ( .A(key_s1[125]), .B(signal_3660), .S(n286), .Z(
        signal_3917) );
  MUX2_X1 cell_1240_Ins_0_U1 ( .A(key_s0[126]), .B(signal_1679), .S(n288), .Z(
        signal_1927) );
  MUX2_X1 cell_1240_Ins_1_U1 ( .A(key_s1[126]), .B(signal_3661), .S(n288), .Z(
        signal_3919) );
  MUX2_X1 cell_1241_Ins_0_U1 ( .A(key_s0[127]), .B(signal_1678), .S(n280), .Z(
        signal_1926) );
  MUX2_X1 cell_1241_Ins_1_U1 ( .A(key_s1[127]), .B(signal_3662), .S(n280), .Z(
        signal_3921) );
  MUX2_X1 cell_1242_Ins_0_U1 ( .A(key_s0[112]), .B(signal_1909), .S(n280), .Z(
        signal_1925) );
  MUX2_X1 cell_1242_Ins_1_U1 ( .A(key_s1[112]), .B(signal_2849), .S(n280), .Z(
        signal_2850) );
  MUX2_X1 cell_1243_Ins_0_U1 ( .A(key_s0[113]), .B(signal_1908), .S(n280), .Z(
        signal_1924) );
  MUX2_X1 cell_1243_Ins_1_U1 ( .A(key_s1[113]), .B(signal_2852), .S(n280), .Z(
        signal_2853) );
  MUX2_X1 cell_1244_Ins_0_U1 ( .A(key_s0[114]), .B(signal_1907), .S(n280), .Z(
        signal_1923) );
  MUX2_X1 cell_1244_Ins_1_U1 ( .A(key_s1[114]), .B(signal_2855), .S(n280), .Z(
        signal_2856) );
  MUX2_X1 cell_1245_Ins_0_U1 ( .A(key_s0[115]), .B(signal_1906), .S(n280), .Z(
        signal_1922) );
  MUX2_X1 cell_1245_Ins_1_U1 ( .A(key_s1[115]), .B(signal_2858), .S(n280), .Z(
        signal_2859) );
  MUX2_X1 cell_1246_Ins_0_U1 ( .A(key_s0[116]), .B(signal_1905), .S(n280), .Z(
        signal_1921) );
  MUX2_X1 cell_1246_Ins_1_U1 ( .A(key_s1[116]), .B(signal_2861), .S(n280), .Z(
        signal_2862) );
  MUX2_X1 cell_1247_Ins_0_U1 ( .A(key_s0[117]), .B(signal_1904), .S(n281), .Z(
        signal_1920) );
  MUX2_X1 cell_1247_Ins_1_U1 ( .A(key_s1[117]), .B(signal_2864), .S(n281), .Z(
        signal_2865) );
  MUX2_X1 cell_1248_Ins_0_U1 ( .A(key_s0[118]), .B(signal_1903), .S(n281), .Z(
        signal_1919) );
  MUX2_X1 cell_1248_Ins_1_U1 ( .A(key_s1[118]), .B(signal_2867), .S(n281), .Z(
        signal_2868) );
  MUX2_X1 cell_1249_Ins_0_U1 ( .A(key_s0[119]), .B(signal_1902), .S(n281), .Z(
        signal_1918) );
  MUX2_X1 cell_1249_Ins_1_U1 ( .A(key_s1[119]), .B(signal_2870), .S(n281), .Z(
        signal_2871) );
  MUX2_X1 cell_1250_Ins_0_U1 ( .A(key_s0[104]), .B(signal_1893), .S(n281), .Z(
        signal_1917) );
  MUX2_X1 cell_1250_Ins_1_U1 ( .A(key_s1[104]), .B(signal_2873), .S(n281), .Z(
        signal_2874) );
  MUX2_X1 cell_1251_Ins_0_U1 ( .A(key_s0[105]), .B(signal_1892), .S(n281), .Z(
        signal_1916) );
  MUX2_X1 cell_1251_Ins_1_U1 ( .A(key_s1[105]), .B(signal_2876), .S(n281), .Z(
        signal_2877) );
  MUX2_X1 cell_1252_Ins_0_U1 ( .A(key_s0[106]), .B(signal_1891), .S(n281), .Z(
        signal_1915) );
  MUX2_X1 cell_1252_Ins_1_U1 ( .A(key_s1[106]), .B(signal_2879), .S(n281), .Z(
        signal_2880) );
  MUX2_X1 cell_1253_Ins_0_U1 ( .A(key_s0[107]), .B(signal_1890), .S(n281), .Z(
        signal_1914) );
  MUX2_X1 cell_1253_Ins_1_U1 ( .A(key_s1[107]), .B(signal_2882), .S(n281), .Z(
        signal_2883) );
  MUX2_X1 cell_1254_Ins_0_U1 ( .A(key_s0[108]), .B(signal_1889), .S(n282), .Z(
        signal_1913) );
  MUX2_X1 cell_1254_Ins_1_U1 ( .A(key_s1[108]), .B(signal_2885), .S(n282), .Z(
        signal_2886) );
  MUX2_X1 cell_1255_Ins_0_U1 ( .A(key_s0[109]), .B(signal_1888), .S(n282), .Z(
        signal_1912) );
  MUX2_X1 cell_1255_Ins_1_U1 ( .A(key_s1[109]), .B(signal_2888), .S(n282), .Z(
        signal_2889) );
  MUX2_X1 cell_1256_Ins_0_U1 ( .A(key_s0[110]), .B(signal_1887), .S(n282), .Z(
        signal_1911) );
  MUX2_X1 cell_1256_Ins_1_U1 ( .A(key_s1[110]), .B(signal_2891), .S(n282), .Z(
        signal_2892) );
  MUX2_X1 cell_1257_Ins_0_U1 ( .A(key_s0[111]), .B(signal_1886), .S(n282), .Z(
        signal_1910) );
  MUX2_X1 cell_1257_Ins_1_U1 ( .A(key_s1[111]), .B(signal_2894), .S(n282), .Z(
        signal_2895) );
  MUX2_X1 cell_1258_Ins_0_U1 ( .A(key_s0[96]), .B(signal_1877), .S(n282), .Z(
        signal_1901) );
  MUX2_X1 cell_1258_Ins_1_U1 ( .A(key_s1[96]), .B(signal_2897), .S(n282), .Z(
        signal_2898) );
  MUX2_X1 cell_1259_Ins_0_U1 ( .A(key_s0[97]), .B(signal_1876), .S(n282), .Z(
        signal_1900) );
  MUX2_X1 cell_1259_Ins_1_U1 ( .A(key_s1[97]), .B(signal_2900), .S(n282), .Z(
        signal_2901) );
  MUX2_X1 cell_1260_Ins_0_U1 ( .A(key_s0[98]), .B(signal_1875), .S(n282), .Z(
        signal_1899) );
  MUX2_X1 cell_1260_Ins_1_U1 ( .A(key_s1[98]), .B(signal_2903), .S(n282), .Z(
        signal_2904) );
  MUX2_X1 cell_1261_Ins_0_U1 ( .A(key_s0[99]), .B(signal_1874), .S(n283), .Z(
        signal_1898) );
  MUX2_X1 cell_1261_Ins_1_U1 ( .A(key_s1[99]), .B(signal_2906), .S(n283), .Z(
        signal_2907) );
  MUX2_X1 cell_1262_Ins_0_U1 ( .A(key_s0[100]), .B(signal_1873), .S(n283), .Z(
        signal_1897) );
  MUX2_X1 cell_1262_Ins_1_U1 ( .A(key_s1[100]), .B(signal_2909), .S(n283), .Z(
        signal_2910) );
  MUX2_X1 cell_1263_Ins_0_U1 ( .A(key_s0[101]), .B(signal_1872), .S(n283), .Z(
        signal_1896) );
  MUX2_X1 cell_1263_Ins_1_U1 ( .A(key_s1[101]), .B(signal_2912), .S(n283), .Z(
        signal_2913) );
  MUX2_X1 cell_1264_Ins_0_U1 ( .A(key_s0[102]), .B(signal_1871), .S(n283), .Z(
        signal_1895) );
  MUX2_X1 cell_1264_Ins_1_U1 ( .A(key_s1[102]), .B(signal_2915), .S(n283), .Z(
        signal_2916) );
  MUX2_X1 cell_1265_Ins_0_U1 ( .A(key_s0[103]), .B(signal_1870), .S(n283), .Z(
        signal_1894) );
  MUX2_X1 cell_1265_Ins_1_U1 ( .A(key_s1[103]), .B(signal_2918), .S(n283), .Z(
        signal_2919) );
  MUX2_X1 cell_1266_Ins_0_U1 ( .A(key_s0[88]), .B(signal_1861), .S(n283), .Z(
        signal_1885) );
  MUX2_X1 cell_1266_Ins_1_U1 ( .A(key_s1[88]), .B(signal_2921), .S(n283), .Z(
        signal_2922) );
  MUX2_X1 cell_1267_Ins_0_U1 ( .A(key_s0[89]), .B(signal_1860), .S(n283), .Z(
        signal_1884) );
  MUX2_X1 cell_1267_Ins_1_U1 ( .A(key_s1[89]), .B(signal_2924), .S(n283), .Z(
        signal_2925) );
  MUX2_X1 cell_1268_Ins_0_U1 ( .A(key_s0[90]), .B(signal_1859), .S(n284), .Z(
        signal_1883) );
  MUX2_X1 cell_1268_Ins_1_U1 ( .A(key_s1[90]), .B(signal_2927), .S(n284), .Z(
        signal_2928) );
  MUX2_X1 cell_1269_Ins_0_U1 ( .A(key_s0[91]), .B(signal_1858), .S(n284), .Z(
        signal_1882) );
  MUX2_X1 cell_1269_Ins_1_U1 ( .A(key_s1[91]), .B(signal_2930), .S(n284), .Z(
        signal_2931) );
  MUX2_X1 cell_1270_Ins_0_U1 ( .A(key_s0[92]), .B(signal_1857), .S(n284), .Z(
        signal_1881) );
  MUX2_X1 cell_1270_Ins_1_U1 ( .A(key_s1[92]), .B(signal_2933), .S(n284), .Z(
        signal_2934) );
  MUX2_X1 cell_1271_Ins_0_U1 ( .A(key_s0[93]), .B(signal_1856), .S(n284), .Z(
        signal_1880) );
  MUX2_X1 cell_1271_Ins_1_U1 ( .A(key_s1[93]), .B(signal_2936), .S(n284), .Z(
        signal_2937) );
  MUX2_X1 cell_1272_Ins_0_U1 ( .A(key_s0[94]), .B(signal_1855), .S(n284), .Z(
        signal_1879) );
  MUX2_X1 cell_1272_Ins_1_U1 ( .A(key_s1[94]), .B(signal_2939), .S(n284), .Z(
        signal_2940) );
  MUX2_X1 cell_1273_Ins_0_U1 ( .A(key_s0[95]), .B(signal_1854), .S(n284), .Z(
        signal_1878) );
  MUX2_X1 cell_1273_Ins_1_U1 ( .A(key_s1[95]), .B(signal_2942), .S(n284), .Z(
        signal_2943) );
  MUX2_X1 cell_1274_Ins_0_U1 ( .A(key_s0[80]), .B(signal_1845), .S(n284), .Z(
        signal_1869) );
  MUX2_X1 cell_1274_Ins_1_U1 ( .A(key_s1[80]), .B(signal_2945), .S(n284), .Z(
        signal_2946) );
  MUX2_X1 cell_1275_Ins_0_U1 ( .A(key_s0[81]), .B(signal_1844), .S(n285), .Z(
        signal_1868) );
  MUX2_X1 cell_1275_Ins_1_U1 ( .A(key_s1[81]), .B(signal_2948), .S(n285), .Z(
        signal_2949) );
  MUX2_X1 cell_1276_Ins_0_U1 ( .A(key_s0[82]), .B(signal_1843), .S(n285), .Z(
        signal_1867) );
  MUX2_X1 cell_1276_Ins_1_U1 ( .A(key_s1[82]), .B(signal_2951), .S(n285), .Z(
        signal_2952) );
  MUX2_X1 cell_1277_Ins_0_U1 ( .A(key_s0[83]), .B(signal_1842), .S(n285), .Z(
        signal_1866) );
  MUX2_X1 cell_1277_Ins_1_U1 ( .A(key_s1[83]), .B(signal_2954), .S(n285), .Z(
        signal_2955) );
  MUX2_X1 cell_1278_Ins_0_U1 ( .A(key_s0[84]), .B(signal_1841), .S(n285), .Z(
        signal_1865) );
  MUX2_X1 cell_1278_Ins_1_U1 ( .A(key_s1[84]), .B(signal_2957), .S(n285), .Z(
        signal_2958) );
  MUX2_X1 cell_1279_Ins_0_U1 ( .A(key_s0[85]), .B(signal_1840), .S(n285), .Z(
        signal_1864) );
  MUX2_X1 cell_1279_Ins_1_U1 ( .A(key_s1[85]), .B(signal_2960), .S(n285), .Z(
        signal_2961) );
  MUX2_X1 cell_1280_Ins_0_U1 ( .A(key_s0[86]), .B(signal_1839), .S(n285), .Z(
        signal_1863) );
  MUX2_X1 cell_1280_Ins_1_U1 ( .A(key_s1[86]), .B(signal_2963), .S(n285), .Z(
        signal_2964) );
  MUX2_X1 cell_1281_Ins_0_U1 ( .A(key_s0[87]), .B(signal_1838), .S(n285), .Z(
        signal_1862) );
  MUX2_X1 cell_1281_Ins_1_U1 ( .A(key_s1[87]), .B(signal_2966), .S(n285), .Z(
        signal_2967) );
  MUX2_X1 cell_1282_Ins_0_U1 ( .A(key_s0[72]), .B(signal_1509), .S(n286), .Z(
        signal_1853) );
  MUX2_X1 cell_1282_Ins_1_U1 ( .A(key_s1[72]), .B(signal_2969), .S(n286), .Z(
        signal_2970) );
  MUX2_X1 cell_1283_Ins_0_U1 ( .A(key_s0[73]), .B(signal_1508), .S(n286), .Z(
        signal_1852) );
  MUX2_X1 cell_1283_Ins_1_U1 ( .A(key_s1[73]), .B(signal_2972), .S(n286), .Z(
        signal_2973) );
  MUX2_X1 cell_1284_Ins_0_U1 ( .A(key_s0[74]), .B(signal_1507), .S(n286), .Z(
        signal_1851) );
  MUX2_X1 cell_1284_Ins_1_U1 ( .A(key_s1[74]), .B(signal_2975), .S(n286), .Z(
        signal_2976) );
  MUX2_X1 cell_1285_Ins_0_U1 ( .A(key_s0[75]), .B(signal_1506), .S(n286), .Z(
        signal_1850) );
  MUX2_X1 cell_1285_Ins_1_U1 ( .A(key_s1[75]), .B(signal_2978), .S(n286), .Z(
        signal_2979) );
  MUX2_X1 cell_1286_Ins_0_U1 ( .A(key_s0[76]), .B(signal_1505), .S(n286), .Z(
        signal_1849) );
  MUX2_X1 cell_1286_Ins_1_U1 ( .A(key_s1[76]), .B(signal_2981), .S(n286), .Z(
        signal_2982) );
  MUX2_X1 cell_1287_Ins_0_U1 ( .A(key_s0[77]), .B(signal_1504), .S(n286), .Z(
        signal_1848) );
  MUX2_X1 cell_1287_Ins_1_U1 ( .A(key_s1[77]), .B(signal_2984), .S(n286), .Z(
        signal_2985) );
  MUX2_X1 cell_1288_Ins_0_U1 ( .A(key_s0[78]), .B(signal_1503), .S(n286), .Z(
        signal_1847) );
  MUX2_X1 cell_1288_Ins_1_U1 ( .A(key_s1[78]), .B(signal_2987), .S(n286), .Z(
        signal_2988) );
  MUX2_X1 cell_1289_Ins_0_U1 ( .A(key_s0[79]), .B(signal_1502), .S(n287), .Z(
        signal_1846) );
  MUX2_X1 cell_1289_Ins_1_U1 ( .A(key_s1[79]), .B(signal_2990), .S(n287), .Z(
        signal_2991) );
  MUX2_X1 cell_1290_Ins_0_U1 ( .A(key_s0[64]), .B(signal_1821), .S(n287), .Z(
        signal_1837) );
  MUX2_X1 cell_1290_Ins_1_U1 ( .A(key_s1[64]), .B(signal_2993), .S(n287), .Z(
        signal_2994) );
  MUX2_X1 cell_1291_Ins_0_U1 ( .A(key_s0[65]), .B(signal_1820), .S(n287), .Z(
        signal_1836) );
  MUX2_X1 cell_1291_Ins_1_U1 ( .A(key_s1[65]), .B(signal_2996), .S(n287), .Z(
        signal_2997) );
  MUX2_X1 cell_1292_Ins_0_U1 ( .A(key_s0[66]), .B(signal_1819), .S(n287), .Z(
        signal_1835) );
  MUX2_X1 cell_1292_Ins_1_U1 ( .A(key_s1[66]), .B(signal_2999), .S(n287), .Z(
        signal_3000) );
  MUX2_X1 cell_1293_Ins_0_U1 ( .A(key_s0[67]), .B(signal_1818), .S(n287), .Z(
        signal_1834) );
  MUX2_X1 cell_1293_Ins_1_U1 ( .A(key_s1[67]), .B(signal_3002), .S(n287), .Z(
        signal_3003) );
  MUX2_X1 cell_1294_Ins_0_U1 ( .A(key_s0[68]), .B(signal_1817), .S(n287), .Z(
        signal_1833) );
  MUX2_X1 cell_1294_Ins_1_U1 ( .A(key_s1[68]), .B(signal_3005), .S(n287), .Z(
        signal_3006) );
  MUX2_X1 cell_1295_Ins_0_U1 ( .A(key_s0[69]), .B(signal_1816), .S(n287), .Z(
        signal_1832) );
  MUX2_X1 cell_1295_Ins_1_U1 ( .A(key_s1[69]), .B(signal_3008), .S(n287), .Z(
        signal_3009) );
  MUX2_X1 cell_1296_Ins_0_U1 ( .A(key_s0[70]), .B(signal_1815), .S(n288), .Z(
        signal_1831) );
  MUX2_X1 cell_1296_Ins_1_U1 ( .A(key_s1[70]), .B(signal_3011), .S(n288), .Z(
        signal_3012) );
  MUX2_X1 cell_1297_Ins_0_U1 ( .A(key_s0[71]), .B(signal_1814), .S(n288), .Z(
        signal_1830) );
  MUX2_X1 cell_1297_Ins_1_U1 ( .A(key_s1[71]), .B(signal_3014), .S(n288), .Z(
        signal_3015) );
  MUX2_X1 cell_1298_Ins_0_U1 ( .A(key_s0[56]), .B(signal_1805), .S(n288), .Z(
        signal_1829) );
  MUX2_X1 cell_1298_Ins_1_U1 ( .A(key_s1[56]), .B(signal_3017), .S(n288), .Z(
        signal_3018) );
  MUX2_X1 cell_1299_Ins_0_U1 ( .A(key_s0[57]), .B(signal_1804), .S(n288), .Z(
        signal_1828) );
  MUX2_X1 cell_1299_Ins_1_U1 ( .A(key_s1[57]), .B(signal_3020), .S(n288), .Z(
        signal_3021) );
  MUX2_X1 cell_1300_Ins_0_U1 ( .A(key_s0[58]), .B(signal_1803), .S(n288), .Z(
        signal_1827) );
  MUX2_X1 cell_1300_Ins_1_U1 ( .A(key_s1[58]), .B(signal_3023), .S(n288), .Z(
        signal_3024) );
  MUX2_X1 cell_1301_Ins_0_U1 ( .A(key_s0[59]), .B(signal_1802), .S(n288), .Z(
        signal_1826) );
  MUX2_X1 cell_1301_Ins_1_U1 ( .A(key_s1[59]), .B(signal_3026), .S(n288), .Z(
        signal_3027) );
  MUX2_X1 cell_1302_Ins_0_U1 ( .A(key_s0[60]), .B(signal_1801), .S(n289), .Z(
        signal_1825) );
  MUX2_X1 cell_1302_Ins_1_U1 ( .A(key_s1[60]), .B(signal_3029), .S(n289), .Z(
        signal_3030) );
  MUX2_X1 cell_1303_Ins_0_U1 ( .A(key_s0[61]), .B(signal_1800), .S(n289), .Z(
        signal_1824) );
  MUX2_X1 cell_1303_Ins_1_U1 ( .A(key_s1[61]), .B(signal_3032), .S(n289), .Z(
        signal_3033) );
  MUX2_X1 cell_1304_Ins_0_U1 ( .A(key_s0[62]), .B(signal_1799), .S(n289), .Z(
        signal_1823) );
  MUX2_X1 cell_1304_Ins_1_U1 ( .A(key_s1[62]), .B(signal_3035), .S(n289), .Z(
        signal_3036) );
  MUX2_X1 cell_1305_Ins_0_U1 ( .A(key_s0[63]), .B(signal_1798), .S(n289), .Z(
        signal_1822) );
  MUX2_X1 cell_1305_Ins_1_U1 ( .A(key_s1[63]), .B(signal_3038), .S(n289), .Z(
        signal_3039) );
  MUX2_X1 cell_1306_Ins_0_U1 ( .A(key_s0[48]), .B(signal_1789), .S(n289), .Z(
        signal_1813) );
  MUX2_X1 cell_1306_Ins_1_U1 ( .A(key_s1[48]), .B(signal_3041), .S(n289), .Z(
        signal_3042) );
  MUX2_X1 cell_1307_Ins_0_U1 ( .A(key_s0[49]), .B(signal_1788), .S(n289), .Z(
        signal_1812) );
  MUX2_X1 cell_1307_Ins_1_U1 ( .A(key_s1[49]), .B(signal_3044), .S(n289), .Z(
        signal_3045) );
  MUX2_X1 cell_1308_Ins_0_U1 ( .A(key_s0[50]), .B(signal_1787), .S(n299), .Z(
        signal_1811) );
  MUX2_X1 cell_1308_Ins_1_U1 ( .A(key_s1[50]), .B(signal_3047), .S(n299), .Z(
        signal_3048) );
  MUX2_X1 cell_1309_Ins_0_U1 ( .A(key_s0[51]), .B(signal_1786), .S(n289), .Z(
        signal_1810) );
  MUX2_X1 cell_1309_Ins_1_U1 ( .A(key_s1[51]), .B(signal_3050), .S(n289), .Z(
        signal_3051) );
  MUX2_X1 cell_1310_Ins_0_U1 ( .A(key_s0[52]), .B(signal_1785), .S(n290), .Z(
        signal_1809) );
  MUX2_X1 cell_1310_Ins_1_U1 ( .A(key_s1[52]), .B(signal_3053), .S(n290), .Z(
        signal_3054) );
  MUX2_X1 cell_1311_Ins_0_U1 ( .A(key_s0[53]), .B(signal_1784), .S(n290), .Z(
        signal_1808) );
  MUX2_X1 cell_1311_Ins_1_U1 ( .A(key_s1[53]), .B(signal_3056), .S(n290), .Z(
        signal_3057) );
  MUX2_X1 cell_1312_Ins_0_U1 ( .A(key_s0[54]), .B(signal_1783), .S(n290), .Z(
        signal_1807) );
  MUX2_X1 cell_1312_Ins_1_U1 ( .A(key_s1[54]), .B(signal_3059), .S(n290), .Z(
        signal_3060) );
  MUX2_X1 cell_1313_Ins_0_U1 ( .A(key_s0[55]), .B(signal_1782), .S(n290), .Z(
        signal_1806) );
  MUX2_X1 cell_1313_Ins_1_U1 ( .A(key_s1[55]), .B(signal_3062), .S(n290), .Z(
        signal_3063) );
  MUX2_X1 cell_1314_Ins_0_U1 ( .A(key_s0[40]), .B(signal_1773), .S(n290), .Z(
        signal_1797) );
  MUX2_X1 cell_1314_Ins_1_U1 ( .A(key_s1[40]), .B(signal_3065), .S(n290), .Z(
        signal_3066) );
  MUX2_X1 cell_1315_Ins_0_U1 ( .A(key_s0[41]), .B(signal_1772), .S(n290), .Z(
        signal_1796) );
  MUX2_X1 cell_1315_Ins_1_U1 ( .A(key_s1[41]), .B(signal_3068), .S(n290), .Z(
        signal_3069) );
  MUX2_X1 cell_1316_Ins_0_U1 ( .A(key_s0[42]), .B(signal_1771), .S(n290), .Z(
        signal_1795) );
  MUX2_X1 cell_1316_Ins_1_U1 ( .A(key_s1[42]), .B(signal_3071), .S(n290), .Z(
        signal_3072) );
  MUX2_X1 cell_1317_Ins_0_U1 ( .A(key_s0[43]), .B(signal_1770), .S(n291), .Z(
        signal_1794) );
  MUX2_X1 cell_1317_Ins_1_U1 ( .A(key_s1[43]), .B(signal_3074), .S(n291), .Z(
        signal_3075) );
  MUX2_X1 cell_1318_Ins_0_U1 ( .A(key_s0[44]), .B(signal_1769), .S(n291), .Z(
        signal_1793) );
  MUX2_X1 cell_1318_Ins_1_U1 ( .A(key_s1[44]), .B(signal_3077), .S(n291), .Z(
        signal_3078) );
  MUX2_X1 cell_1319_Ins_0_U1 ( .A(key_s0[45]), .B(signal_1768), .S(n291), .Z(
        signal_1792) );
  MUX2_X1 cell_1319_Ins_1_U1 ( .A(key_s1[45]), .B(signal_3080), .S(n291), .Z(
        signal_3081) );
  MUX2_X1 cell_1320_Ins_0_U1 ( .A(key_s0[46]), .B(signal_1767), .S(n291), .Z(
        signal_1791) );
  MUX2_X1 cell_1320_Ins_1_U1 ( .A(key_s1[46]), .B(signal_3083), .S(n291), .Z(
        signal_3084) );
  MUX2_X1 cell_1321_Ins_0_U1 ( .A(key_s0[47]), .B(signal_1766), .S(n291), .Z(
        signal_1790) );
  MUX2_X1 cell_1321_Ins_1_U1 ( .A(key_s1[47]), .B(signal_3086), .S(n291), .Z(
        signal_3087) );
  MUX2_X1 cell_1322_Ins_0_U1 ( .A(key_s0[32]), .B(signal_1749), .S(n291), .Z(
        signal_1781) );
  MUX2_X1 cell_1322_Ins_1_U1 ( .A(key_s1[32]), .B(signal_3089), .S(n291), .Z(
        signal_3090) );
  MUX2_X1 cell_1323_Ins_0_U1 ( .A(key_s0[33]), .B(signal_1748), .S(n291), .Z(
        signal_1780) );
  MUX2_X1 cell_1323_Ins_1_U1 ( .A(key_s1[33]), .B(signal_3092), .S(n291), .Z(
        signal_3093) );
  MUX2_X1 cell_1324_Ins_0_U1 ( .A(key_s0[34]), .B(signal_1747), .S(n302), .Z(
        signal_1779) );
  MUX2_X1 cell_1324_Ins_1_U1 ( .A(key_s1[34]), .B(signal_3095), .S(n302), .Z(
        signal_3096) );
  MUX2_X1 cell_1325_Ins_0_U1 ( .A(key_s0[35]), .B(signal_1746), .S(n306), .Z(
        signal_1778) );
  MUX2_X1 cell_1325_Ins_1_U1 ( .A(key_s1[35]), .B(signal_3098), .S(n306), .Z(
        signal_3099) );
  MUX2_X1 cell_1326_Ins_0_U1 ( .A(key_s0[36]), .B(signal_1745), .S(n299), .Z(
        signal_1777) );
  MUX2_X1 cell_1326_Ins_1_U1 ( .A(key_s1[36]), .B(signal_3101), .S(n299), .Z(
        signal_3102) );
  MUX2_X1 cell_1327_Ins_0_U1 ( .A(key_s0[37]), .B(signal_1744), .S(n292), .Z(
        signal_1776) );
  MUX2_X1 cell_1327_Ins_1_U1 ( .A(key_s1[37]), .B(signal_3104), .S(n292), .Z(
        signal_3105) );
  MUX2_X1 cell_1328_Ins_0_U1 ( .A(key_s0[38]), .B(signal_1743), .S(n304), .Z(
        signal_1775) );
  MUX2_X1 cell_1328_Ins_1_U1 ( .A(key_s1[38]), .B(signal_3107), .S(n304), .Z(
        signal_3108) );
  MUX2_X1 cell_1329_Ins_0_U1 ( .A(key_s0[39]), .B(signal_1742), .S(n289), .Z(
        signal_1774) );
  MUX2_X1 cell_1329_Ins_1_U1 ( .A(key_s1[39]), .B(signal_3110), .S(n289), .Z(
        signal_3111) );
  MUX2_X1 cell_1330_Ins_0_U1 ( .A(key_s0[24]), .B(signal_1733), .S(n301), .Z(
        signal_1765) );
  MUX2_X1 cell_1330_Ins_1_U1 ( .A(key_s1[24]), .B(signal_3113), .S(n301), .Z(
        signal_3114) );
  MUX2_X1 cell_1331_Ins_0_U1 ( .A(key_s0[25]), .B(signal_1732), .S(n292), .Z(
        signal_1764) );
  MUX2_X1 cell_1331_Ins_1_U1 ( .A(key_s1[25]), .B(signal_3116), .S(n292), .Z(
        signal_3117) );
  MUX2_X1 cell_1332_Ins_0_U1 ( .A(key_s0[26]), .B(signal_1731), .S(n292), .Z(
        signal_1763) );
  MUX2_X1 cell_1332_Ins_1_U1 ( .A(key_s1[26]), .B(signal_3119), .S(n292), .Z(
        signal_3120) );
  MUX2_X1 cell_1333_Ins_0_U1 ( .A(key_s0[27]), .B(signal_1730), .S(n292), .Z(
        signal_1762) );
  MUX2_X1 cell_1333_Ins_1_U1 ( .A(key_s1[27]), .B(signal_3122), .S(n292), .Z(
        signal_3123) );
  MUX2_X1 cell_1334_Ins_0_U1 ( .A(key_s0[28]), .B(signal_1729), .S(n292), .Z(
        signal_1761) );
  MUX2_X1 cell_1334_Ins_1_U1 ( .A(key_s1[28]), .B(signal_3125), .S(n292), .Z(
        signal_3126) );
  MUX2_X1 cell_1335_Ins_0_U1 ( .A(key_s0[29]), .B(signal_1728), .S(n292), .Z(
        signal_1760) );
  MUX2_X1 cell_1335_Ins_1_U1 ( .A(key_s1[29]), .B(signal_3128), .S(n292), .Z(
        signal_3129) );
  MUX2_X1 cell_1336_Ins_0_U1 ( .A(key_s0[30]), .B(signal_1727), .S(n292), .Z(
        signal_1759) );
  MUX2_X1 cell_1336_Ins_1_U1 ( .A(key_s1[30]), .B(signal_3131), .S(n292), .Z(
        signal_3132) );
  MUX2_X1 cell_1337_Ins_0_U1 ( .A(key_s0[31]), .B(signal_1726), .S(n292), .Z(
        signal_1758) );
  MUX2_X1 cell_1337_Ins_1_U1 ( .A(key_s1[31]), .B(signal_3134), .S(n292), .Z(
        signal_3135) );
  MUX2_X1 cell_1338_Ins_0_U1 ( .A(key_s0[16]), .B(signal_1717), .S(n293), .Z(
        signal_1741) );
  MUX2_X1 cell_1338_Ins_1_U1 ( .A(key_s1[16]), .B(signal_3137), .S(n293), .Z(
        signal_3138) );
  MUX2_X1 cell_1339_Ins_0_U1 ( .A(key_s0[17]), .B(signal_1716), .S(n293), .Z(
        signal_1740) );
  MUX2_X1 cell_1339_Ins_1_U1 ( .A(key_s1[17]), .B(signal_3140), .S(n293), .Z(
        signal_3141) );
  MUX2_X1 cell_1340_Ins_0_U1 ( .A(key_s0[18]), .B(signal_1715), .S(n293), .Z(
        signal_1739) );
  MUX2_X1 cell_1340_Ins_1_U1 ( .A(key_s1[18]), .B(signal_3143), .S(n293), .Z(
        signal_3144) );
  MUX2_X1 cell_1341_Ins_0_U1 ( .A(key_s0[19]), .B(signal_1714), .S(n293), .Z(
        signal_1738) );
  MUX2_X1 cell_1341_Ins_1_U1 ( .A(key_s1[19]), .B(signal_3146), .S(n293), .Z(
        signal_3147) );
  MUX2_X1 cell_1342_Ins_0_U1 ( .A(key_s0[20]), .B(signal_1713), .S(n293), .Z(
        signal_1737) );
  MUX2_X1 cell_1342_Ins_1_U1 ( .A(key_s1[20]), .B(signal_3149), .S(n293), .Z(
        signal_3150) );
  MUX2_X1 cell_1343_Ins_0_U1 ( .A(key_s0[21]), .B(signal_1712), .S(n293), .Z(
        signal_1736) );
  MUX2_X1 cell_1343_Ins_1_U1 ( .A(key_s1[21]), .B(signal_3152), .S(n293), .Z(
        signal_3153) );
  MUX2_X1 cell_1344_Ins_0_U1 ( .A(key_s0[22]), .B(signal_1711), .S(n293), .Z(
        signal_1735) );
  MUX2_X1 cell_1344_Ins_1_U1 ( .A(key_s1[22]), .B(signal_3155), .S(n293), .Z(
        signal_3156) );
  MUX2_X1 cell_1345_Ins_0_U1 ( .A(key_s0[23]), .B(signal_1710), .S(n294), .Z(
        signal_1734) );
  MUX2_X1 cell_1345_Ins_1_U1 ( .A(key_s1[23]), .B(signal_3158), .S(n294), .Z(
        signal_3159) );
  MUX2_X1 cell_1346_Ins_0_U1 ( .A(key_s0[8]), .B(signal_1701), .S(n294), .Z(
        signal_1725) );
  MUX2_X1 cell_1346_Ins_1_U1 ( .A(key_s1[8]), .B(signal_3161), .S(n294), .Z(
        signal_3162) );
  MUX2_X1 cell_1347_Ins_0_U1 ( .A(key_s0[9]), .B(signal_1700), .S(n294), .Z(
        signal_1724) );
  MUX2_X1 cell_1347_Ins_1_U1 ( .A(key_s1[9]), .B(signal_3164), .S(n294), .Z(
        signal_3165) );
  MUX2_X1 cell_1348_Ins_0_U1 ( .A(key_s0[10]), .B(signal_1699), .S(n294), .Z(
        signal_1723) );
  MUX2_X1 cell_1348_Ins_1_U1 ( .A(key_s1[10]), .B(signal_3167), .S(n294), .Z(
        signal_3168) );
  MUX2_X1 cell_1349_Ins_0_U1 ( .A(key_s0[11]), .B(signal_1698), .S(n294), .Z(
        signal_1722) );
  MUX2_X1 cell_1349_Ins_1_U1 ( .A(key_s1[11]), .B(signal_3170), .S(n294), .Z(
        signal_3171) );
  MUX2_X1 cell_1350_Ins_0_U1 ( .A(key_s0[12]), .B(signal_1697), .S(n294), .Z(
        signal_1721) );
  MUX2_X1 cell_1350_Ins_1_U1 ( .A(key_s1[12]), .B(signal_3173), .S(n294), .Z(
        signal_3174) );
  MUX2_X1 cell_1351_Ins_0_U1 ( .A(key_s0[13]), .B(signal_1696), .S(n294), .Z(
        signal_1720) );
  MUX2_X1 cell_1351_Ins_1_U1 ( .A(key_s1[13]), .B(signal_3176), .S(n294), .Z(
        signal_3177) );
  MUX2_X1 cell_1352_Ins_0_U1 ( .A(key_s0[14]), .B(signal_1695), .S(n300), .Z(
        signal_1719) );
  MUX2_X1 cell_1352_Ins_1_U1 ( .A(key_s1[14]), .B(signal_3179), .S(n300), .Z(
        signal_3180) );
  MUX2_X1 cell_1353_Ins_0_U1 ( .A(key_s0[15]), .B(signal_1694), .S(n292), .Z(
        signal_1718) );
  MUX2_X1 cell_1353_Ins_1_U1 ( .A(key_s1[15]), .B(signal_3182), .S(n292), .Z(
        signal_3183) );
  MUX2_X1 cell_1354_Ins_0_U1 ( .A(key_s0[0]), .B(signal_1493), .S(n289), .Z(
        signal_1709) );
  MUX2_X1 cell_1354_Ins_1_U1 ( .A(key_s1[0]), .B(signal_2389), .S(n289), .Z(
        signal_3185) );
  MUX2_X1 cell_1355_Ins_0_U1 ( .A(key_s0[1]), .B(signal_1492), .S(n292), .Z(
        signal_1708) );
  MUX2_X1 cell_1355_Ins_1_U1 ( .A(key_s1[1]), .B(signal_2392), .S(n292), .Z(
        signal_3187) );
  MUX2_X1 cell_1356_Ins_0_U1 ( .A(key_s0[2]), .B(signal_1491), .S(n298), .Z(
        signal_1707) );
  MUX2_X1 cell_1356_Ins_1_U1 ( .A(key_s1[2]), .B(signal_2395), .S(n298), .Z(
        signal_3189) );
  MUX2_X1 cell_1357_Ins_0_U1 ( .A(key_s0[3]), .B(signal_1490), .S(n35), .Z(
        signal_1706) );
  MUX2_X1 cell_1357_Ins_1_U1 ( .A(key_s1[3]), .B(signal_2398), .S(n35), .Z(
        signal_3191) );
  MUX2_X1 cell_1358_Ins_0_U1 ( .A(key_s0[4]), .B(signal_1489), .S(n35), .Z(
        signal_1705) );
  MUX2_X1 cell_1358_Ins_1_U1 ( .A(key_s1[4]), .B(signal_2401), .S(n35), .Z(
        signal_3193) );
  MUX2_X1 cell_1359_Ins_0_U1 ( .A(key_s0[5]), .B(signal_1488), .S(n35), .Z(
        signal_1704) );
  MUX2_X1 cell_1359_Ins_1_U1 ( .A(key_s1[5]), .B(signal_2404), .S(n35), .Z(
        signal_3195) );
  MUX2_X1 cell_1360_Ins_0_U1 ( .A(key_s0[6]), .B(signal_1487), .S(n35), .Z(
        signal_1703) );
  MUX2_X1 cell_1360_Ins_1_U1 ( .A(key_s1[6]), .B(signal_2407), .S(n35), .Z(
        signal_3197) );
  MUX2_X1 cell_1361_Ins_0_U1 ( .A(key_s0[7]), .B(signal_1486), .S(n35), .Z(
        signal_1702) );
  MUX2_X1 cell_1361_Ins_1_U1 ( .A(key_s1[7]), .B(signal_2410), .S(n35), .Z(
        signal_3199) );
  XNOR2_X1 cell_1362_Ins0_U1 ( .A(signal_1150), .B(signal_1151), .ZN(
        signal_1454) );
  XOR2_X1 cell_1362_Ins_1_U1 ( .A(signal_2528), .B(signal_2430), .Z(
        signal_3200) );
  XNOR2_X1 cell_1363_Ins0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[31]), 
        .ZN(signal_1151) );
  XOR2_X1 cell_1363_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[31]), 
        .Z(signal_2430) );
  XOR2_X1 cell_1364_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(signal_1934), .Z(
        signal_1150) );
  XOR2_X1 cell_1364_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(signal_2457), .Z(
        signal_2528) );
  XNOR2_X1 cell_1365_Ins0_U1 ( .A(signal_1152), .B(signal_1153), .ZN(
        signal_1455) );
  XOR2_X1 cell_1365_Ins_1_U1 ( .A(signal_2529), .B(signal_2433), .Z(
        signal_3201) );
  XNOR2_X1 cell_1366_Ins0_U1 ( .A(ciphertext_s0[62]), .B(ciphertext_s0[30]), 
        .ZN(signal_1153) );
  XOR2_X1 cell_1366_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(ciphertext_s1[30]), 
        .Z(signal_2433) );
  XOR2_X1 cell_1367_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(signal_1935), .Z(
        signal_1152) );
  XOR2_X1 cell_1367_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(signal_2459), .Z(
        signal_2529) );
  XNOR2_X1 cell_1368_Ins0_U1 ( .A(signal_1154), .B(signal_1155), .ZN(
        signal_1456) );
  XOR2_X1 cell_1368_Ins_1_U1 ( .A(signal_2530), .B(signal_2436), .Z(
        signal_3202) );
  XNOR2_X1 cell_1369_Ins0_U1 ( .A(ciphertext_s0[61]), .B(ciphertext_s0[29]), 
        .ZN(signal_1155) );
  XOR2_X1 cell_1369_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(ciphertext_s1[29]), 
        .Z(signal_2436) );
  XOR2_X1 cell_1370_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(signal_1936), .Z(
        signal_1154) );
  XOR2_X1 cell_1370_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(signal_2461), .Z(
        signal_2530) );
  XNOR2_X1 cell_1371_Ins0_U1 ( .A(signal_1156), .B(signal_1157), .ZN(
        signal_1457) );
  XOR2_X1 cell_1371_Ins_1_U1 ( .A(signal_3203), .B(signal_2439), .Z(
        signal_3244) );
  XNOR2_X1 cell_1372_Ins0_U1 ( .A(ciphertext_s0[60]), .B(ciphertext_s0[28]), 
        .ZN(signal_1157) );
  XOR2_X1 cell_1372_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(ciphertext_s1[28]), 
        .Z(signal_2439) );
  XOR2_X1 cell_1373_Ins_0_U1 ( .A(signal_1942), .B(signal_1937), .Z(
        signal_1156) );
  XOR2_X1 cell_1373_Ins_1_U1 ( .A(signal_2452), .B(signal_2533), .Z(
        signal_3203) );
  XNOR2_X1 cell_1374_Ins0_U1 ( .A(signal_1158), .B(signal_1159), .ZN(
        signal_1458) );
  XOR2_X1 cell_1374_Ins_1_U1 ( .A(signal_3204), .B(signal_2442), .Z(
        signal_3245) );
  XNOR2_X1 cell_1375_Ins0_U1 ( .A(ciphertext_s0[59]), .B(ciphertext_s0[27]), 
        .ZN(signal_1159) );
  XOR2_X1 cell_1375_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(ciphertext_s1[27]), 
        .Z(signal_2442) );
  XOR2_X1 cell_1376_Ins_0_U1 ( .A(signal_1943), .B(signal_1938), .Z(
        signal_1158) );
  XOR2_X1 cell_1376_Ins_1_U1 ( .A(signal_2453), .B(signal_2534), .Z(
        signal_3204) );
  XNOR2_X1 cell_1377_Ins0_U1 ( .A(signal_1160), .B(signal_1161), .ZN(
        signal_1459) );
  XOR2_X1 cell_1377_Ins_1_U1 ( .A(signal_2531), .B(signal_2445), .Z(
        signal_3205) );
  XNOR2_X1 cell_1378_Ins0_U1 ( .A(ciphertext_s0[58]), .B(ciphertext_s0[26]), 
        .ZN(signal_1161) );
  XOR2_X1 cell_1378_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(ciphertext_s1[26]), 
        .Z(signal_2445) );
  XOR2_X1 cell_1379_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(signal_1939), .Z(
        signal_1160) );
  XOR2_X1 cell_1379_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(signal_2464), .Z(
        signal_2531) );
  XNOR2_X1 cell_1380_Ins0_U1 ( .A(signal_1162), .B(signal_1163), .ZN(
        signal_1460) );
  XOR2_X1 cell_1380_Ins_1_U1 ( .A(signal_3206), .B(signal_2448), .Z(
        signal_3246) );
  XNOR2_X1 cell_1381_Ins0_U1 ( .A(ciphertext_s0[25]), .B(ciphertext_s0[57]), 
        .ZN(signal_1163) );
  XOR2_X1 cell_1381_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(ciphertext_s1[57]), 
        .Z(signal_2448) );
  XOR2_X1 cell_1382_Ins_0_U1 ( .A(signal_1945), .B(signal_1940), .Z(
        signal_1162) );
  XOR2_X1 cell_1382_Ins_1_U1 ( .A(signal_2454), .B(signal_2535), .Z(
        signal_3206) );
  XNOR2_X1 cell_1383_Ins0_U1 ( .A(signal_1164), .B(signal_1165), .ZN(
        signal_1461) );
  XOR2_X1 cell_1383_Ins_1_U1 ( .A(signal_2532), .B(signal_2451), .Z(
        signal_3207) );
  XNOR2_X1 cell_1384_Ins0_U1 ( .A(ciphertext_s0[24]), .B(ciphertext_s0[56]), 
        .ZN(signal_1165) );
  XOR2_X1 cell_1384_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(ciphertext_s1[56]), 
        .Z(signal_2451) );
  XOR2_X1 cell_1385_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(signal_1941), .Z(
        signal_1164) );
  XOR2_X1 cell_1385_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(signal_2466), .Z(
        signal_2532) );
  XOR2_X1 cell_1386_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[123]), 
        .Z(signal_1942) );
  XOR2_X1 cell_1386_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[123]), 
        .Z(signal_2452) );
  XOR2_X1 cell_1387_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[122]), 
        .Z(signal_1943) );
  XOR2_X1 cell_1387_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[122]), 
        .Z(signal_2453) );
  XOR2_X1 cell_1388_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[120]), 
        .Z(signal_1945) );
  XOR2_X1 cell_1388_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[120]), 
        .Z(signal_2454) );
  XOR2_X1 cell_1389_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[94]), 
        .Z(signal_1934) );
  XOR2_X1 cell_1389_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[94]), 
        .Z(signal_2457) );
  XOR2_X1 cell_1390_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(ciphertext_s0[93]), 
        .Z(signal_1935) );
  XOR2_X1 cell_1390_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(ciphertext_s1[93]), 
        .Z(signal_2459) );
  XOR2_X1 cell_1391_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(ciphertext_s0[92]), 
        .Z(signal_1936) );
  XOR2_X1 cell_1391_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(ciphertext_s1[92]), 
        .Z(signal_2461) );
  XOR2_X1 cell_1392_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(signal_1946), .Z(
        signal_1937) );
  XOR2_X1 cell_1392_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(signal_2468), .Z(
        signal_2533) );
  XOR2_X1 cell_1393_Ins_0_U1 ( .A(ciphertext_s0[91]), .B(signal_1947), .Z(
        signal_1938) );
  XOR2_X1 cell_1393_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(signal_2469), .Z(
        signal_2534) );
  XOR2_X1 cell_1394_Ins_0_U1 ( .A(ciphertext_s0[90]), .B(ciphertext_s0[89]), 
        .Z(signal_1939) );
  XOR2_X1 cell_1394_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(ciphertext_s1[89]), 
        .Z(signal_2464) );
  XOR2_X1 cell_1395_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(signal_1949), .Z(
        signal_1940) );
  XOR2_X1 cell_1395_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(signal_2470), .Z(
        signal_2535) );
  XOR2_X1 cell_1396_Ins_0_U1 ( .A(ciphertext_s0[88]), .B(ciphertext_s0[95]), 
        .Z(signal_1941) );
  XOR2_X1 cell_1396_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(ciphertext_s1[95]), 
        .Z(signal_2466) );
  XOR2_X1 cell_1397_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[91]), 
        .Z(signal_1946) );
  XOR2_X1 cell_1397_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[91]), 
        .Z(signal_2468) );
  XOR2_X1 cell_1398_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[90]), 
        .Z(signal_1947) );
  XOR2_X1 cell_1398_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[90]), 
        .Z(signal_2469) );
  XOR2_X1 cell_1399_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[88]), 
        .Z(signal_1949) );
  XOR2_X1 cell_1399_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[88]), 
        .Z(signal_2470) );
  XNOR2_X1 cell_1400_Ins0_U1 ( .A(signal_1166), .B(signal_1167), .ZN(
        signal_1462) );
  XOR2_X1 cell_1400_Ins_1_U1 ( .A(signal_2536), .B(signal_2471), .Z(
        signal_3208) );
  XNOR2_X1 cell_1401_Ins0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[127]), 
        .ZN(signal_1167) );
  XOR2_X1 cell_1401_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[127]), 
        .Z(signal_2471) );
  XOR2_X1 cell_1402_Ins_0_U1 ( .A(ciphertext_s0[94]), .B(signal_1950), .Z(
        signal_1166) );
  XOR2_X1 cell_1402_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(signal_2482), .Z(
        signal_2536) );
  XNOR2_X1 cell_1403_Ins0_U1 ( .A(signal_1168), .B(signal_1169), .ZN(
        signal_1463) );
  XOR2_X1 cell_1403_Ins_1_U1 ( .A(signal_2537), .B(signal_2472), .Z(
        signal_3209) );
  XNOR2_X1 cell_1404_Ins0_U1 ( .A(ciphertext_s0[30]), .B(ciphertext_s0[126]), 
        .ZN(signal_1169) );
  XOR2_X1 cell_1404_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(ciphertext_s1[126]), 
        .Z(signal_2472) );
  XOR2_X1 cell_1405_Ins_0_U1 ( .A(ciphertext_s0[93]), .B(signal_1951), .Z(
        signal_1168) );
  XOR2_X1 cell_1405_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(signal_2483), .Z(
        signal_2537) );
  XNOR2_X1 cell_1406_Ins0_U1 ( .A(signal_1170), .B(signal_1171), .ZN(
        signal_1464) );
  XOR2_X1 cell_1406_Ins_1_U1 ( .A(signal_2538), .B(signal_2473), .Z(
        signal_3210) );
  XNOR2_X1 cell_1407_Ins0_U1 ( .A(ciphertext_s0[29]), .B(ciphertext_s0[125]), 
        .ZN(signal_1171) );
  XOR2_X1 cell_1407_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(ciphertext_s1[125]), 
        .Z(signal_2473) );
  XOR2_X1 cell_1408_Ins_0_U1 ( .A(ciphertext_s0[92]), .B(signal_1952), .Z(
        signal_1170) );
  XOR2_X1 cell_1408_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(signal_2484), .Z(
        signal_2538) );
  XNOR2_X1 cell_1409_Ins0_U1 ( .A(signal_1172), .B(signal_1173), .ZN(
        signal_1465) );
  XOR2_X1 cell_1409_Ins_1_U1 ( .A(signal_3211), .B(signal_2474), .Z(
        signal_3247) );
  XNOR2_X1 cell_1410_Ins0_U1 ( .A(ciphertext_s0[28]), .B(ciphertext_s0[124]), 
        .ZN(signal_1173) );
  XOR2_X1 cell_1410_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(ciphertext_s1[124]), 
        .Z(signal_2474) );
  XOR2_X1 cell_1411_Ins_0_U1 ( .A(signal_1184), .B(signal_1953), .Z(
        signal_1172) );
  XOR2_X1 cell_1411_Ins_1_U1 ( .A(signal_2479), .B(signal_2541), .Z(
        signal_3211) );
  XNOR2_X1 cell_1412_Ins0_U1 ( .A(signal_1174), .B(signal_1175), .ZN(
        signal_1466) );
  XOR2_X1 cell_1412_Ins_1_U1 ( .A(signal_3212), .B(signal_2475), .Z(
        signal_3248) );
  XNOR2_X1 cell_1413_Ins0_U1 ( .A(ciphertext_s0[27]), .B(ciphertext_s0[123]), 
        .ZN(signal_1175) );
  XOR2_X1 cell_1413_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(ciphertext_s1[123]), 
        .Z(signal_2475) );
  XOR2_X1 cell_1414_Ins_0_U1 ( .A(signal_1183), .B(signal_1954), .Z(
        signal_1174) );
  XOR2_X1 cell_1414_Ins_1_U1 ( .A(signal_2480), .B(signal_2542), .Z(
        signal_3212) );
  XNOR2_X1 cell_1415_Ins0_U1 ( .A(signal_1176), .B(signal_1177), .ZN(
        signal_1467) );
  XOR2_X1 cell_1415_Ins_1_U1 ( .A(signal_2539), .B(signal_2476), .Z(
        signal_3213) );
  XNOR2_X1 cell_1416_Ins0_U1 ( .A(ciphertext_s0[26]), .B(ciphertext_s0[122]), 
        .ZN(signal_1177) );
  XOR2_X1 cell_1416_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(ciphertext_s1[122]), 
        .Z(signal_2476) );
  XOR2_X1 cell_1417_Ins_0_U1 ( .A(ciphertext_s0[89]), .B(signal_1955), .Z(
        signal_1176) );
  XOR2_X1 cell_1417_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(signal_2485), .Z(
        signal_2539) );
  XNOR2_X1 cell_1418_Ins0_U1 ( .A(signal_1178), .B(signal_1179), .ZN(
        signal_1468) );
  XOR2_X1 cell_1418_Ins_1_U1 ( .A(signal_3214), .B(signal_2477), .Z(
        signal_3249) );
  XNOR2_X1 cell_1419_Ins0_U1 ( .A(ciphertext_s0[121]), .B(ciphertext_s0[25]), 
        .ZN(signal_1179) );
  XOR2_X1 cell_1419_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(ciphertext_s1[25]), 
        .Z(signal_2477) );
  XOR2_X1 cell_1420_Ins_0_U1 ( .A(signal_1182), .B(signal_1956), .Z(
        signal_1178) );
  XOR2_X1 cell_1420_Ins_1_U1 ( .A(signal_2481), .B(signal_2543), .Z(
        signal_3214) );
  XNOR2_X1 cell_1421_Ins0_U1 ( .A(signal_1180), .B(signal_1181), .ZN(
        signal_1469) );
  XOR2_X1 cell_1421_Ins_1_U1 ( .A(signal_2540), .B(signal_2478), .Z(
        signal_3215) );
  XNOR2_X1 cell_1422_Ins0_U1 ( .A(ciphertext_s0[120]), .B(ciphertext_s0[24]), 
        .ZN(signal_1181) );
  XOR2_X1 cell_1422_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(ciphertext_s1[24]), 
        .Z(signal_2478) );
  XOR2_X1 cell_1423_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(signal_1957), .Z(
        signal_1180) );
  XOR2_X1 cell_1423_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(signal_2486), .Z(
        signal_2540) );
  XOR2_X1 cell_1424_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[91]), 
        .Z(signal_1184) );
  XOR2_X1 cell_1424_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[91]), 
        .Z(signal_2479) );
  XOR2_X1 cell_1425_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[90]), 
        .Z(signal_1183) );
  XOR2_X1 cell_1425_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[90]), 
        .Z(signal_2480) );
  XOR2_X1 cell_1426_Ins_0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[88]), 
        .Z(signal_1182) );
  XOR2_X1 cell_1426_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[88]), 
        .Z(signal_2481) );
  XOR2_X1 cell_1427_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[62]), 
        .Z(signal_1950) );
  XOR2_X1 cell_1427_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[62]), 
        .Z(signal_2482) );
  XOR2_X1 cell_1428_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(ciphertext_s0[61]), 
        .Z(signal_1951) );
  XOR2_X1 cell_1428_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(ciphertext_s1[61]), 
        .Z(signal_2483) );
  XOR2_X1 cell_1429_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(ciphertext_s0[60]), 
        .Z(signal_1952) );
  XOR2_X1 cell_1429_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(ciphertext_s1[60]), 
        .Z(signal_2484) );
  XOR2_X1 cell_1430_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(signal_1958), .Z(
        signal_1953) );
  XOR2_X1 cell_1430_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(signal_2487), .Z(
        signal_2541) );
  XOR2_X1 cell_1431_Ins_0_U1 ( .A(ciphertext_s0[59]), .B(signal_1959), .Z(
        signal_1954) );
  XOR2_X1 cell_1431_Ins_1_U1 ( .A(ciphertext_s1[59]), .B(signal_2488), .Z(
        signal_2542) );
  XOR2_X1 cell_1432_Ins_0_U1 ( .A(ciphertext_s0[58]), .B(ciphertext_s0[57]), 
        .Z(signal_1955) );
  XOR2_X1 cell_1432_Ins_1_U1 ( .A(ciphertext_s1[58]), .B(ciphertext_s1[57]), 
        .Z(signal_2485) );
  XOR2_X1 cell_1433_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(signal_1961), .Z(
        signal_1956) );
  XOR2_X1 cell_1433_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(signal_2489), .Z(
        signal_2543) );
  XOR2_X1 cell_1434_Ins_0_U1 ( .A(ciphertext_s0[56]), .B(ciphertext_s0[63]), 
        .Z(signal_1957) );
  XOR2_X1 cell_1434_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(ciphertext_s1[63]), 
        .Z(signal_2486) );
  XOR2_X1 cell_1435_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[59]), 
        .Z(signal_1958) );
  XOR2_X1 cell_1435_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[59]), 
        .Z(signal_2487) );
  XOR2_X1 cell_1436_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[58]), 
        .Z(signal_1959) );
  XOR2_X1 cell_1436_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[58]), 
        .Z(signal_2488) );
  XOR2_X1 cell_1437_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[56]), 
        .Z(signal_1961) );
  XOR2_X1 cell_1437_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[56]), 
        .Z(signal_2489) );
  XNOR2_X1 cell_1438_Ins0_U1 ( .A(signal_1185), .B(signal_1186), .ZN(
        signal_1470) );
  XOR2_X1 cell_1438_Ins_1_U1 ( .A(signal_2544), .B(signal_2490), .Z(
        signal_3216) );
  XNOR2_X1 cell_1439_Ins0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[95]), 
        .ZN(signal_1186) );
  XOR2_X1 cell_1439_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[95]), 
        .Z(signal_2490) );
  XOR2_X1 cell_1440_Ins_0_U1 ( .A(ciphertext_s0[62]), .B(signal_1962), .Z(
        signal_1185) );
  XOR2_X1 cell_1440_Ins_1_U1 ( .A(ciphertext_s1[62]), .B(signal_2501), .Z(
        signal_2544) );
  XNOR2_X1 cell_1441_Ins0_U1 ( .A(signal_1187), .B(signal_1188), .ZN(
        signal_1471) );
  XOR2_X1 cell_1441_Ins_1_U1 ( .A(signal_2545), .B(signal_2491), .Z(
        signal_3217) );
  XNOR2_X1 cell_1442_Ins0_U1 ( .A(ciphertext_s0[126]), .B(ciphertext_s0[94]), 
        .ZN(signal_1188) );
  XOR2_X1 cell_1442_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(ciphertext_s1[94]), 
        .Z(signal_2491) );
  XOR2_X1 cell_1443_Ins_0_U1 ( .A(ciphertext_s0[61]), .B(signal_1963), .Z(
        signal_1187) );
  XOR2_X1 cell_1443_Ins_1_U1 ( .A(ciphertext_s1[61]), .B(signal_2502), .Z(
        signal_2545) );
  XNOR2_X1 cell_1444_Ins0_U1 ( .A(signal_1189), .B(signal_1190), .ZN(
        signal_1472) );
  XOR2_X1 cell_1444_Ins_1_U1 ( .A(signal_2546), .B(signal_2492), .Z(
        signal_3218) );
  XNOR2_X1 cell_1445_Ins0_U1 ( .A(ciphertext_s0[125]), .B(ciphertext_s0[93]), 
        .ZN(signal_1190) );
  XOR2_X1 cell_1445_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(ciphertext_s1[93]), 
        .Z(signal_2492) );
  XOR2_X1 cell_1446_Ins_0_U1 ( .A(ciphertext_s0[60]), .B(signal_1964), .Z(
        signal_1189) );
  XOR2_X1 cell_1446_Ins_1_U1 ( .A(ciphertext_s1[60]), .B(signal_2503), .Z(
        signal_2546) );
  XNOR2_X1 cell_1447_Ins0_U1 ( .A(signal_1191), .B(signal_1192), .ZN(
        signal_1473) );
  XOR2_X1 cell_1447_Ins_1_U1 ( .A(signal_3219), .B(signal_2493), .Z(
        signal_3250) );
  XNOR2_X1 cell_1448_Ins0_U1 ( .A(ciphertext_s0[124]), .B(ciphertext_s0[92]), 
        .ZN(signal_1192) );
  XOR2_X1 cell_1448_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(ciphertext_s1[92]), 
        .Z(signal_2493) );
  XOR2_X1 cell_1449_Ins_0_U1 ( .A(signal_1203), .B(signal_1965), .Z(
        signal_1191) );
  XOR2_X1 cell_1449_Ins_1_U1 ( .A(signal_2498), .B(signal_2549), .Z(
        signal_3219) );
  XNOR2_X1 cell_1450_Ins0_U1 ( .A(signal_1193), .B(signal_1194), .ZN(
        signal_1474) );
  XOR2_X1 cell_1450_Ins_1_U1 ( .A(signal_3220), .B(signal_2494), .Z(
        signal_3251) );
  XNOR2_X1 cell_1451_Ins0_U1 ( .A(ciphertext_s0[123]), .B(ciphertext_s0[91]), 
        .ZN(signal_1194) );
  XOR2_X1 cell_1451_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(ciphertext_s1[91]), 
        .Z(signal_2494) );
  XOR2_X1 cell_1452_Ins_0_U1 ( .A(signal_1202), .B(signal_1966), .Z(
        signal_1193) );
  XOR2_X1 cell_1452_Ins_1_U1 ( .A(signal_2499), .B(signal_2550), .Z(
        signal_3220) );
  XNOR2_X1 cell_1453_Ins0_U1 ( .A(signal_1195), .B(signal_1196), .ZN(
        signal_1475) );
  XOR2_X1 cell_1453_Ins_1_U1 ( .A(signal_2547), .B(signal_2495), .Z(
        signal_3221) );
  XNOR2_X1 cell_1454_Ins0_U1 ( .A(ciphertext_s0[122]), .B(ciphertext_s0[90]), 
        .ZN(signal_1196) );
  XOR2_X1 cell_1454_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(ciphertext_s1[90]), 
        .Z(signal_2495) );
  XOR2_X1 cell_1455_Ins_0_U1 ( .A(ciphertext_s0[57]), .B(signal_1967), .Z(
        signal_1195) );
  XOR2_X1 cell_1455_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(signal_2504), .Z(
        signal_2547) );
  XNOR2_X1 cell_1456_Ins0_U1 ( .A(signal_1197), .B(signal_1198), .ZN(
        signal_1476) );
  XOR2_X1 cell_1456_Ins_1_U1 ( .A(signal_3222), .B(signal_2496), .Z(
        signal_3252) );
  XNOR2_X1 cell_1457_Ins0_U1 ( .A(ciphertext_s0[89]), .B(ciphertext_s0[121]), 
        .ZN(signal_1198) );
  XOR2_X1 cell_1457_Ins_1_U1 ( .A(ciphertext_s1[89]), .B(ciphertext_s1[121]), 
        .Z(signal_2496) );
  XOR2_X1 cell_1458_Ins_0_U1 ( .A(signal_1201), .B(signal_1968), .Z(
        signal_1197) );
  XOR2_X1 cell_1458_Ins_1_U1 ( .A(signal_2500), .B(signal_2551), .Z(
        signal_3222) );
  XNOR2_X1 cell_1459_Ins0_U1 ( .A(signal_1199), .B(signal_1200), .ZN(
        signal_1477) );
  XOR2_X1 cell_1459_Ins_1_U1 ( .A(signal_2548), .B(signal_2497), .Z(
        signal_3223) );
  XNOR2_X1 cell_1460_Ins0_U1 ( .A(ciphertext_s0[88]), .B(ciphertext_s0[120]), 
        .ZN(signal_1200) );
  XOR2_X1 cell_1460_Ins_1_U1 ( .A(ciphertext_s1[88]), .B(ciphertext_s1[120]), 
        .Z(signal_2497) );
  XOR2_X1 cell_1461_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(signal_1969), .Z(
        signal_1199) );
  XOR2_X1 cell_1461_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(signal_2505), .Z(
        signal_2548) );
  XOR2_X1 cell_1462_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[59]), 
        .Z(signal_1203) );
  XOR2_X1 cell_1462_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[59]), 
        .Z(signal_2498) );
  XOR2_X1 cell_1463_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[58]), 
        .Z(signal_1202) );
  XOR2_X1 cell_1463_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[58]), 
        .Z(signal_2499) );
  XOR2_X1 cell_1464_Ins_0_U1 ( .A(ciphertext_s0[63]), .B(ciphertext_s0[56]), 
        .Z(signal_1201) );
  XOR2_X1 cell_1464_Ins_1_U1 ( .A(ciphertext_s1[63]), .B(ciphertext_s1[56]), 
        .Z(signal_2500) );
  XOR2_X1 cell_1465_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[30]), 
        .Z(signal_1962) );
  XOR2_X1 cell_1465_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[30]), 
        .Z(signal_2501) );
  XOR2_X1 cell_1466_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(ciphertext_s0[29]), 
        .Z(signal_1963) );
  XOR2_X1 cell_1466_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(ciphertext_s1[29]), 
        .Z(signal_2502) );
  XOR2_X1 cell_1467_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(ciphertext_s0[28]), 
        .Z(signal_1964) );
  XOR2_X1 cell_1467_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(ciphertext_s1[28]), 
        .Z(signal_2503) );
  XOR2_X1 cell_1468_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(signal_1970), .Z(
        signal_1965) );
  XOR2_X1 cell_1468_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(signal_2506), .Z(
        signal_2549) );
  XOR2_X1 cell_1469_Ins_0_U1 ( .A(ciphertext_s0[27]), .B(signal_1971), .Z(
        signal_1966) );
  XOR2_X1 cell_1469_Ins_1_U1 ( .A(ciphertext_s1[27]), .B(signal_2507), .Z(
        signal_2550) );
  XOR2_X1 cell_1470_Ins_0_U1 ( .A(ciphertext_s0[26]), .B(ciphertext_s0[25]), 
        .Z(signal_1967) );
  XOR2_X1 cell_1470_Ins_1_U1 ( .A(ciphertext_s1[26]), .B(ciphertext_s1[25]), 
        .Z(signal_2504) );
  XOR2_X1 cell_1471_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(signal_1973), .Z(
        signal_1968) );
  XOR2_X1 cell_1471_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(signal_2508), .Z(
        signal_2551) );
  XOR2_X1 cell_1472_Ins_0_U1 ( .A(ciphertext_s0[24]), .B(ciphertext_s0[31]), 
        .Z(signal_1969) );
  XOR2_X1 cell_1472_Ins_1_U1 ( .A(ciphertext_s1[24]), .B(ciphertext_s1[31]), 
        .Z(signal_2505) );
  XOR2_X1 cell_1473_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[27]), 
        .Z(signal_1970) );
  XOR2_X1 cell_1473_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[27]), 
        .Z(signal_2506) );
  XOR2_X1 cell_1474_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[26]), 
        .Z(signal_1971) );
  XOR2_X1 cell_1474_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[26]), 
        .Z(signal_2507) );
  XOR2_X1 cell_1475_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[24]), 
        .Z(signal_1973) );
  XOR2_X1 cell_1475_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[24]), 
        .Z(signal_2508) );
  XNOR2_X1 cell_1476_Ins0_U1 ( .A(signal_1204), .B(signal_1205), .ZN(
        signal_1478) );
  XOR2_X1 cell_1476_Ins_1_U1 ( .A(signal_2552), .B(signal_2509), .Z(
        signal_3224) );
  XNOR2_X1 cell_1477_Ins0_U1 ( .A(ciphertext_s0[95]), .B(ciphertext_s0[63]), 
        .ZN(signal_1205) );
  XOR2_X1 cell_1477_Ins_1_U1 ( .A(ciphertext_s1[95]), .B(ciphertext_s1[63]), 
        .Z(signal_2509) );
  XOR2_X1 cell_1478_Ins_0_U1 ( .A(ciphertext_s0[30]), .B(signal_1974), .Z(
        signal_1204) );
  XOR2_X1 cell_1478_Ins_1_U1 ( .A(ciphertext_s1[30]), .B(signal_2520), .Z(
        signal_2552) );
  XNOR2_X1 cell_1479_Ins0_U1 ( .A(signal_1206), .B(signal_1207), .ZN(
        signal_1479) );
  XOR2_X1 cell_1479_Ins_1_U1 ( .A(signal_2553), .B(signal_2510), .Z(
        signal_3225) );
  XNOR2_X1 cell_1480_Ins0_U1 ( .A(ciphertext_s0[94]), .B(ciphertext_s0[62]), 
        .ZN(signal_1207) );
  XOR2_X1 cell_1480_Ins_1_U1 ( .A(ciphertext_s1[94]), .B(ciphertext_s1[62]), 
        .Z(signal_2510) );
  XOR2_X1 cell_1481_Ins_0_U1 ( .A(ciphertext_s0[29]), .B(signal_1975), .Z(
        signal_1206) );
  XOR2_X1 cell_1481_Ins_1_U1 ( .A(ciphertext_s1[29]), .B(signal_2521), .Z(
        signal_2553) );
  XNOR2_X1 cell_1482_Ins0_U1 ( .A(signal_1208), .B(signal_1209), .ZN(
        signal_1480) );
  XOR2_X1 cell_1482_Ins_1_U1 ( .A(signal_2554), .B(signal_2511), .Z(
        signal_3226) );
  XNOR2_X1 cell_1483_Ins0_U1 ( .A(ciphertext_s0[93]), .B(ciphertext_s0[61]), 
        .ZN(signal_1209) );
  XOR2_X1 cell_1483_Ins_1_U1 ( .A(ciphertext_s1[93]), .B(ciphertext_s1[61]), 
        .Z(signal_2511) );
  XOR2_X1 cell_1484_Ins_0_U1 ( .A(ciphertext_s0[28]), .B(signal_1976), .Z(
        signal_1208) );
  XOR2_X1 cell_1484_Ins_1_U1 ( .A(ciphertext_s1[28]), .B(signal_2522), .Z(
        signal_2554) );
  XNOR2_X1 cell_1485_Ins0_U1 ( .A(signal_1210), .B(signal_1211), .ZN(
        signal_1481) );
  XOR2_X1 cell_1485_Ins_1_U1 ( .A(signal_3227), .B(signal_2512), .Z(
        signal_3253) );
  XNOR2_X1 cell_1486_Ins0_U1 ( .A(ciphertext_s0[92]), .B(ciphertext_s0[60]), 
        .ZN(signal_1211) );
  XOR2_X1 cell_1486_Ins_1_U1 ( .A(ciphertext_s1[92]), .B(ciphertext_s1[60]), 
        .Z(signal_2512) );
  XOR2_X1 cell_1487_Ins_0_U1 ( .A(signal_1222), .B(signal_1977), .Z(
        signal_1210) );
  XOR2_X1 cell_1487_Ins_1_U1 ( .A(signal_2517), .B(signal_2557), .Z(
        signal_3227) );
  XNOR2_X1 cell_1488_Ins0_U1 ( .A(signal_1212), .B(signal_1213), .ZN(
        signal_1482) );
  XOR2_X1 cell_1488_Ins_1_U1 ( .A(signal_3228), .B(signal_2513), .Z(
        signal_3254) );
  XNOR2_X1 cell_1489_Ins0_U1 ( .A(ciphertext_s0[91]), .B(ciphertext_s0[59]), 
        .ZN(signal_1213) );
  XOR2_X1 cell_1489_Ins_1_U1 ( .A(ciphertext_s1[91]), .B(ciphertext_s1[59]), 
        .Z(signal_2513) );
  XOR2_X1 cell_1490_Ins_0_U1 ( .A(signal_1221), .B(signal_1978), .Z(
        signal_1212) );
  XOR2_X1 cell_1490_Ins_1_U1 ( .A(signal_2518), .B(signal_2558), .Z(
        signal_3228) );
  XNOR2_X1 cell_1491_Ins0_U1 ( .A(signal_1214), .B(signal_1215), .ZN(
        signal_1483) );
  XOR2_X1 cell_1491_Ins_1_U1 ( .A(signal_2555), .B(signal_2514), .Z(
        signal_3229) );
  XNOR2_X1 cell_1492_Ins0_U1 ( .A(ciphertext_s0[90]), .B(ciphertext_s0[58]), 
        .ZN(signal_1215) );
  XOR2_X1 cell_1492_Ins_1_U1 ( .A(ciphertext_s1[90]), .B(ciphertext_s1[58]), 
        .Z(signal_2514) );
  XOR2_X1 cell_1493_Ins_0_U1 ( .A(ciphertext_s0[25]), .B(signal_1979), .Z(
        signal_1214) );
  XOR2_X1 cell_1493_Ins_1_U1 ( .A(ciphertext_s1[25]), .B(signal_2523), .Z(
        signal_2555) );
  XNOR2_X1 cell_1494_Ins0_U1 ( .A(signal_1216), .B(signal_1217), .ZN(
        signal_1484) );
  XOR2_X1 cell_1494_Ins_1_U1 ( .A(signal_3230), .B(signal_2515), .Z(
        signal_3255) );
  XNOR2_X1 cell_1495_Ins0_U1 ( .A(ciphertext_s0[57]), .B(ciphertext_s0[89]), 
        .ZN(signal_1217) );
  XOR2_X1 cell_1495_Ins_1_U1 ( .A(ciphertext_s1[57]), .B(ciphertext_s1[89]), 
        .Z(signal_2515) );
  XOR2_X1 cell_1496_Ins_0_U1 ( .A(signal_1220), .B(signal_1980), .Z(
        signal_1216) );
  XOR2_X1 cell_1496_Ins_1_U1 ( .A(signal_2519), .B(signal_2559), .Z(
        signal_3230) );
  XNOR2_X1 cell_1497_Ins0_U1 ( .A(signal_1218), .B(signal_1219), .ZN(
        signal_1485) );
  XOR2_X1 cell_1497_Ins_1_U1 ( .A(signal_2556), .B(signal_2516), .Z(
        signal_3231) );
  XNOR2_X1 cell_1498_Ins0_U1 ( .A(ciphertext_s0[56]), .B(ciphertext_s0[88]), 
        .ZN(signal_1219) );
  XOR2_X1 cell_1498_Ins_1_U1 ( .A(ciphertext_s1[56]), .B(ciphertext_s1[88]), 
        .Z(signal_2516) );
  XOR2_X1 cell_1499_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(signal_1981), .Z(
        signal_1218) );
  XOR2_X1 cell_1499_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(signal_2524), .Z(
        signal_2556) );
  XOR2_X1 cell_1500_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[27]), 
        .Z(signal_1222) );
  XOR2_X1 cell_1500_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[27]), 
        .Z(signal_2517) );
  XOR2_X1 cell_1501_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[26]), 
        .Z(signal_1221) );
  XOR2_X1 cell_1501_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[26]), 
        .Z(signal_2518) );
  XOR2_X1 cell_1502_Ins_0_U1 ( .A(ciphertext_s0[31]), .B(ciphertext_s0[24]), 
        .Z(signal_1220) );
  XOR2_X1 cell_1502_Ins_1_U1 ( .A(ciphertext_s1[31]), .B(ciphertext_s1[24]), 
        .Z(signal_2519) );
  XOR2_X1 cell_1503_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[126]), 
        .Z(signal_1974) );
  XOR2_X1 cell_1503_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[126]), 
        .Z(signal_2520) );
  XOR2_X1 cell_1504_Ins_0_U1 ( .A(ciphertext_s0[126]), .B(ciphertext_s0[125]), 
        .Z(signal_1975) );
  XOR2_X1 cell_1504_Ins_1_U1 ( .A(ciphertext_s1[126]), .B(ciphertext_s1[125]), 
        .Z(signal_2521) );
  XOR2_X1 cell_1505_Ins_0_U1 ( .A(ciphertext_s0[125]), .B(ciphertext_s0[124]), 
        .Z(signal_1976) );
  XOR2_X1 cell_1505_Ins_1_U1 ( .A(ciphertext_s1[125]), .B(ciphertext_s1[124]), 
        .Z(signal_2522) );
  XOR2_X1 cell_1506_Ins_0_U1 ( .A(ciphertext_s0[124]), .B(signal_1225), .Z(
        signal_1977) );
  XOR2_X1 cell_1506_Ins_1_U1 ( .A(ciphertext_s1[124]), .B(signal_2525), .Z(
        signal_2557) );
  XOR2_X1 cell_1507_Ins_0_U1 ( .A(ciphertext_s0[123]), .B(signal_1224), .Z(
        signal_1978) );
  XOR2_X1 cell_1507_Ins_1_U1 ( .A(ciphertext_s1[123]), .B(signal_2526), .Z(
        signal_2558) );
  XOR2_X1 cell_1508_Ins_0_U1 ( .A(ciphertext_s0[122]), .B(ciphertext_s0[121]), 
        .Z(signal_1979) );
  XOR2_X1 cell_1508_Ins_1_U1 ( .A(ciphertext_s1[122]), .B(ciphertext_s1[121]), 
        .Z(signal_2523) );
  XOR2_X1 cell_1509_Ins_0_U1 ( .A(ciphertext_s0[121]), .B(signal_1223), .Z(
        signal_1980) );
  XOR2_X1 cell_1509_Ins_1_U1 ( .A(ciphertext_s1[121]), .B(signal_2527), .Z(
        signal_2559) );
  XOR2_X1 cell_1510_Ins_0_U1 ( .A(ciphertext_s0[120]), .B(ciphertext_s0[127]), 
        .Z(signal_1981) );
  XOR2_X1 cell_1510_Ins_1_U1 ( .A(ciphertext_s1[120]), .B(ciphertext_s1[127]), 
        .Z(signal_2524) );
  XOR2_X1 cell_1511_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[123]), 
        .Z(signal_1225) );
  XOR2_X1 cell_1511_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[123]), 
        .Z(signal_2525) );
  XOR2_X1 cell_1512_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[122]), 
        .Z(signal_1224) );
  XOR2_X1 cell_1512_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[122]), 
        .Z(signal_2526) );
  XOR2_X1 cell_1513_Ins_0_U1 ( .A(ciphertext_s0[127]), .B(ciphertext_s0[120]), 
        .Z(signal_1223) );
  XOR2_X1 cell_1513_Ins_1_U1 ( .A(ciphertext_s1[127]), .B(ciphertext_s1[120]), 
        .Z(signal_2527) );
  MUX2_X1 cell_1576_Ins_0_U1 ( .A(signal_1413), .B(signal_1509), .S(n242), .Z(
        signal_1517) );
  MUX2_X1 cell_1576_Ins_1_U1 ( .A(signal_2390), .B(signal_2969), .S(n242), .Z(
        signal_3232) );
  MUX2_X1 cell_1577_Ins_0_U1 ( .A(signal_1412), .B(signal_1508), .S(n242), .Z(
        signal_1516) );
  MUX2_X1 cell_1577_Ins_1_U1 ( .A(signal_2393), .B(signal_2972), .S(n242), .Z(
        signal_3233) );
  MUX2_X1 cell_1578_Ins_0_U1 ( .A(signal_1411), .B(signal_1507), .S(n242), .Z(
        signal_1515) );
  MUX2_X1 cell_1578_Ins_1_U1 ( .A(signal_2396), .B(signal_2975), .S(n242), .Z(
        signal_3234) );
  MUX2_X1 cell_1579_Ins_0_U1 ( .A(signal_1410), .B(signal_1506), .S(n242), .Z(
        signal_1514) );
  MUX2_X1 cell_1579_Ins_1_U1 ( .A(signal_2399), .B(signal_2978), .S(n242), .Z(
        signal_3235) );
  MUX2_X1 cell_1580_Ins_0_U1 ( .A(signal_1409), .B(signal_1505), .S(n319), .Z(
        signal_1513) );
  MUX2_X1 cell_1580_Ins_1_U1 ( .A(signal_2402), .B(signal_2981), .S(n319), .Z(
        signal_3236) );
  MUX2_X1 cell_1581_Ins_0_U1 ( .A(signal_1408), .B(signal_1504), .S(n308), .Z(
        signal_1512) );
  MUX2_X1 cell_1581_Ins_1_U1 ( .A(signal_2405), .B(signal_2984), .S(n308), .Z(
        signal_3237) );
  MUX2_X1 cell_1582_Ins_0_U1 ( .A(signal_1407), .B(signal_1503), .S(n317), .Z(
        signal_1511) );
  MUX2_X1 cell_1582_Ins_1_U1 ( .A(signal_2408), .B(signal_2987), .S(n317), .Z(
        signal_3238) );
  MUX2_X1 cell_1583_Ins_0_U1 ( .A(signal_1406), .B(signal_1502), .S(n307), .Z(
        signal_1510) );
  MUX2_X1 cell_1583_Ins_1_U1 ( .A(signal_2411), .B(signal_2990), .S(n307), .Z(
        signal_3239) );
  NOR2_X1 cell_2128_U21 ( .A1(start), .A2(cell_2128_n26), .ZN(cell_2128_n9) );
  NOR2_X1 cell_2128_U20 ( .A1(start), .A2(cell_2128_n25), .ZN(cell_2128_n8) );
  NOR2_X1 cell_2128_U19 ( .A1(start), .A2(cell_2128_n24), .ZN(cell_2128_n7) );
  NOR2_X1 cell_2128_U18 ( .A1(start), .A2(cell_2128_n23), .ZN(cell_2128_n6) );
  NOR2_X1 cell_2128_U17 ( .A1(start), .A2(cell_2128_n22), .ZN(cell_2128_n5) );
  NOR2_X1 cell_2128_U16 ( .A1(start), .A2(cell_2128_n21), .ZN(cell_2128_n4) );
  NOR2_X1 cell_2128_U15 ( .A1(start), .A2(cell_2128_n20), .ZN(cell_2128_n3) );
  NOR2_X1 cell_2128_U14 ( .A1(start), .A2(cell_2128_n19), .ZN(cell_2128_n2) );
  NOR2_X1 cell_2128_U13 ( .A1(start), .A2(cell_2128_n33), .ZN(cell_2128_n16)
         );
  NOR2_X1 cell_2128_U12 ( .A1(start), .A2(cell_2128_n32), .ZN(cell_2128_n15)
         );
  NOR2_X1 cell_2128_U11 ( .A1(start), .A2(cell_2128_n31), .ZN(cell_2128_n14)
         );
  NOR2_X1 cell_2128_U10 ( .A1(start), .A2(cell_2128_n30), .ZN(cell_2128_n13)
         );
  NOR2_X1 cell_2128_U9 ( .A1(start), .A2(cell_2128_n29), .ZN(cell_2128_n12) );
  NOR2_X1 cell_2128_U8 ( .A1(start), .A2(cell_2128_n28), .ZN(cell_2128_n11) );
  NOR2_X1 cell_2128_U7 ( .A1(start), .A2(cell_2128_n27), .ZN(cell_2128_n10) );
  NOR2_X1 cell_2128_U6 ( .A1(start), .A2(cell_2128_n18), .ZN(cell_2128_n1) );
  NAND2_X1 cell_2128_U5 ( .A1(cell_2128_n34), .A2(cell_2128_n17), .ZN(
        cell_2128_N19) );
  INV_X1 cell_2128_U4 ( .A(start), .ZN(cell_2128_n17) );
  AND2_X1 cell_2128_U3 ( .A1(cell_2128_LatchedEnable), .A2(clk), .ZN(
        signal_4640) );
  DFF_X1 cell_2128_ShiftRegister_reg_2_ ( .D(cell_2128_n1), .CK(clk), .Q(), 
        .QN(cell_2128_n19) );
  DFF_X1 cell_2128_ShiftRegister_reg_3_ ( .D(cell_2128_n2), .CK(clk), .Q(), 
        .QN(cell_2128_n20) );
  DFF_X1 cell_2128_ShiftRegister_reg_4_ ( .D(cell_2128_n3), .CK(clk), .Q(), 
        .QN(cell_2128_n21) );
  DFF_X1 cell_2128_ShiftRegister_reg_5_ ( .D(cell_2128_n4), .CK(clk), .Q(), 
        .QN(cell_2128_n22) );
  DFF_X1 cell_2128_ShiftRegister_reg_6_ ( .D(cell_2128_n5), .CK(clk), .Q(), 
        .QN(cell_2128_n23) );
  DFF_X1 cell_2128_ShiftRegister_reg_7_ ( .D(cell_2128_n6), .CK(clk), .Q(), 
        .QN(cell_2128_n24) );
  DFF_X1 cell_2128_ShiftRegister_reg_8_ ( .D(cell_2128_n7), .CK(clk), .Q(), 
        .QN(cell_2128_n25) );
  DFF_X1 cell_2128_ShiftRegister_reg_9_ ( .D(cell_2128_n8), .CK(clk), .Q(), 
        .QN(cell_2128_n26) );
  DFF_X1 cell_2128_ShiftRegister_reg_10_ ( .D(cell_2128_n9), .CK(clk), .Q(), 
        .QN(cell_2128_n27) );
  DFF_X1 cell_2128_ShiftRegister_reg_11_ ( .D(cell_2128_n10), .CK(clk), .Q(), 
        .QN(cell_2128_n28) );
  DFF_X1 cell_2128_ShiftRegister_reg_12_ ( .D(cell_2128_n11), .CK(clk), .Q(), 
        .QN(cell_2128_n29) );
  DFF_X1 cell_2128_ShiftRegister_reg_13_ ( .D(cell_2128_n12), .CK(clk), .Q(), 
        .QN(cell_2128_n30) );
  DFF_X1 cell_2128_ShiftRegister_reg_14_ ( .D(cell_2128_n13), .CK(clk), .Q(), 
        .QN(cell_2128_n31) );
  DFF_X1 cell_2128_ShiftRegister_reg_15_ ( .D(cell_2128_n14), .CK(clk), .Q(), 
        .QN(cell_2128_n32) );
  DFF_X1 cell_2128_ShiftRegister_reg_16_ ( .D(cell_2128_n15), .CK(clk), .Q(), 
        .QN(cell_2128_n33) );
  DFF_X1 cell_2128_ShiftRegister_reg_17_ ( .D(cell_2128_n16), .CK(clk), .Q(
        cell_2128_ShiftRegister_17_), .QN(cell_2128_n34) );
  DLL_X1 cell_2128_LatchedEnable_reg ( .D(cell_2128_N19), .GN(clk), .Q(
        cell_2128_LatchedEnable) );
  DLL_X1 cell_2128_Synch_reg ( .D(cell_2128_ShiftRegister_17_), .GN(clk), .Q(
        Synch) );
  DFF_X1 cell_2128_ShiftRegister_reg_1_ ( .D(cell_2128_N19), .CK(clk), .Q(), 
        .QN(cell_2128_n18) );
  XOR2_X1 cell_1714_U4 ( .A(1'b0), .B(1'b0), .Z(cell_1714_and_in[1]) );
  XOR2_X1 cell_1714_U3 ( .A(1'b1), .B(1'b0), .Z(cell_1714_and_in[0]) );
  XOR2_X1 cell_1714_U2 ( .A(1'b0), .B(cell_1714_and_out[1]), .Z(signal_3256)
         );
  XOR2_X1 cell_1714_U1 ( .A(1'b1), .B(cell_1714_and_out[0]), .Z(signal_1982)
         );
  XOR2_X1 cell_1714_a_HPC2_and_U14 ( .A(Fresh[0]), .B(cell_1714_and_in[0]), 
        .Z(cell_1714_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1714_a_HPC2_and_U13 ( .A(Fresh[0]), .B(cell_1714_and_in[1]), 
        .Z(cell_1714_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1714_a_HPC2_and_U12 ( .A1(cell_1714_a_HPC2_and_a_reg[1]), .A2(
        cell_1714_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1714_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1714_a_HPC2_and_U11 ( .A1(cell_1714_a_HPC2_and_a_reg[0]), .A2(
        cell_1714_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1714_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1714_a_HPC2_and_U10 ( .A1(signal_3232), .A2(
        cell_1714_a_HPC2_and_n9), .ZN(cell_1714_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1714_a_HPC2_and_U9 ( .A1(signal_1517), .A2(
        cell_1714_a_HPC2_and_n9), .ZN(cell_1714_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1714_a_HPC2_and_U8 ( .A(Fresh[0]), .ZN(cell_1714_a_HPC2_and_n9)
         );
  AND2_X1 cell_1714_a_HPC2_and_U7 ( .A1(cell_1714_and_in[1]), .A2(signal_3232), 
        .ZN(cell_1714_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1714_a_HPC2_and_U6 ( .A1(cell_1714_and_in[0]), .A2(signal_1517), 
        .ZN(cell_1714_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1714_a_HPC2_and_U5 ( .A(cell_1714_a_HPC2_and_n8), .B(
        cell_1714_a_HPC2_and_z_1__1_), .ZN(cell_1714_and_out[1]) );
  XNOR2_X1 cell_1714_a_HPC2_and_U4 ( .A(
        cell_1714_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1714_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1714_a_HPC2_and_n8) );
  XNOR2_X1 cell_1714_a_HPC2_and_U3 ( .A(cell_1714_a_HPC2_and_n7), .B(
        cell_1714_a_HPC2_and_z_0__0_), .ZN(cell_1714_and_out[0]) );
  XNOR2_X1 cell_1714_a_HPC2_and_U2 ( .A(
        cell_1714_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1714_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1714_a_HPC2_and_n7) );
  DFF_X1 cell_1714_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1714_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1714_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1517), 
        .CK(clk), .Q(cell_1714_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1714_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1714_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3232), 
        .CK(clk), .Q(cell_1714_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1714_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1714_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1714_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1715_U4 ( .A(1'b0), .B(cell_1715_and_out[1]), .Z(signal_3257)
         );
  XOR2_X1 cell_1715_U3 ( .A(1'b1), .B(cell_1715_and_out[0]), .Z(signal_1983)
         );
  XOR2_X1 cell_1715_U2 ( .A(1'b0), .B(1'b0), .Z(cell_1715_and_in[1]) );
  XOR2_X1 cell_1715_U1 ( .A(1'b1), .B(1'b0), .Z(cell_1715_and_in[0]) );
  XOR2_X1 cell_1715_a_HPC2_and_U14 ( .A(Fresh[1]), .B(cell_1715_and_in[0]), 
        .Z(cell_1715_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1715_a_HPC2_and_U13 ( .A(Fresh[1]), .B(cell_1715_and_in[1]), 
        .Z(cell_1715_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1715_a_HPC2_and_U12 ( .A1(cell_1715_a_HPC2_and_a_reg[1]), .A2(
        cell_1715_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1715_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1715_a_HPC2_and_U11 ( .A1(cell_1715_a_HPC2_and_a_reg[0]), .A2(
        cell_1715_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1715_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1715_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1715_a_HPC2_and_n9), 
        .ZN(cell_1715_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1715_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1715_a_HPC2_and_n9), 
        .ZN(cell_1715_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1715_a_HPC2_and_U8 ( .A(Fresh[1]), .ZN(cell_1715_a_HPC2_and_n9)
         );
  AND2_X1 cell_1715_a_HPC2_and_U7 ( .A1(cell_1715_and_in[1]), .A2(n393), .ZN(
        cell_1715_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1715_a_HPC2_and_U6 ( .A1(cell_1715_and_in[0]), .A2(n392), .ZN(
        cell_1715_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1715_a_HPC2_and_U5 ( .A(cell_1715_a_HPC2_and_n8), .B(
        cell_1715_a_HPC2_and_z_1__1_), .ZN(cell_1715_and_out[1]) );
  XNOR2_X1 cell_1715_a_HPC2_and_U4 ( .A(
        cell_1715_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1715_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1715_a_HPC2_and_n8) );
  XNOR2_X1 cell_1715_a_HPC2_and_U3 ( .A(cell_1715_a_HPC2_and_n7), .B(
        cell_1715_a_HPC2_and_z_0__0_), .ZN(cell_1715_and_out[0]) );
  XNOR2_X1 cell_1715_a_HPC2_and_U2 ( .A(
        cell_1715_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1715_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1715_a_HPC2_and_n7) );
  DFF_X1 cell_1715_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1715_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1715_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1715_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1715_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1715_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1715_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1715_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1715_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1715_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1716_U4 ( .A(1'b0), .B(1'b0), .Z(cell_1716_and_in[1]) );
  XOR2_X1 cell_1716_U3 ( .A(1'b0), .B(1'b1), .Z(cell_1716_and_in[0]) );
  XOR2_X1 cell_1716_U2 ( .A(1'b0), .B(cell_1716_and_out[1]), .Z(signal_3258)
         );
  XOR2_X1 cell_1716_U1 ( .A(1'b0), .B(cell_1716_and_out[0]), .Z(signal_1984)
         );
  XOR2_X1 cell_1716_a_HPC2_and_U14 ( .A(Fresh[2]), .B(cell_1716_and_in[0]), 
        .Z(cell_1716_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1716_a_HPC2_and_U13 ( .A(Fresh[2]), .B(cell_1716_and_in[1]), 
        .Z(cell_1716_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1716_a_HPC2_and_U12 ( .A1(cell_1716_a_HPC2_and_a_reg[1]), .A2(
        cell_1716_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1716_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1716_a_HPC2_and_U11 ( .A1(cell_1716_a_HPC2_and_a_reg[0]), .A2(
        cell_1716_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1716_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1716_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1716_a_HPC2_and_n9), 
        .ZN(cell_1716_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1716_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1716_a_HPC2_and_n9), 
        .ZN(cell_1716_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1716_a_HPC2_and_U8 ( .A(Fresh[2]), .ZN(cell_1716_a_HPC2_and_n9)
         );
  AND2_X1 cell_1716_a_HPC2_and_U7 ( .A1(cell_1716_and_in[1]), .A2(n393), .ZN(
        cell_1716_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1716_a_HPC2_and_U6 ( .A1(cell_1716_and_in[0]), .A2(n392), .ZN(
        cell_1716_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1716_a_HPC2_and_U5 ( .A(cell_1716_a_HPC2_and_n8), .B(
        cell_1716_a_HPC2_and_z_1__1_), .ZN(cell_1716_and_out[1]) );
  XNOR2_X1 cell_1716_a_HPC2_and_U4 ( .A(
        cell_1716_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1716_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1716_a_HPC2_and_n8) );
  XNOR2_X1 cell_1716_a_HPC2_and_U3 ( .A(cell_1716_a_HPC2_and_n7), .B(
        cell_1716_a_HPC2_and_z_0__0_), .ZN(cell_1716_and_out[0]) );
  XNOR2_X1 cell_1716_a_HPC2_and_U2 ( .A(
        cell_1716_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1716_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1716_a_HPC2_and_n7) );
  DFF_X1 cell_1716_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1716_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1716_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1716_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1716_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1716_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1716_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1716_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1716_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1716_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1717_U4 ( .A(1'b0), .B(cell_1717_and_out[1]), .Z(signal_3259)
         );
  XOR2_X1 cell_1717_U3 ( .A(1'b0), .B(cell_1717_and_out[0]), .Z(signal_1985)
         );
  XOR2_X1 cell_1717_U2 ( .A(1'b0), .B(1'b0), .Z(cell_1717_and_in[1]) );
  XOR2_X1 cell_1717_U1 ( .A(1'b0), .B(1'b1), .Z(cell_1717_and_in[0]) );
  XOR2_X1 cell_1717_a_HPC2_and_U14 ( .A(Fresh[3]), .B(cell_1717_and_in[0]), 
        .Z(cell_1717_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1717_a_HPC2_and_U13 ( .A(Fresh[3]), .B(cell_1717_and_in[1]), 
        .Z(cell_1717_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1717_a_HPC2_and_U12 ( .A1(cell_1717_a_HPC2_and_a_reg[1]), .A2(
        cell_1717_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1717_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1717_a_HPC2_and_U11 ( .A1(cell_1717_a_HPC2_and_a_reg[0]), .A2(
        cell_1717_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1717_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1717_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1717_a_HPC2_and_n9), 
        .ZN(cell_1717_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1717_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1717_a_HPC2_and_n9), 
        .ZN(cell_1717_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1717_a_HPC2_and_U8 ( .A(Fresh[3]), .ZN(cell_1717_a_HPC2_and_n9)
         );
  AND2_X1 cell_1717_a_HPC2_and_U7 ( .A1(cell_1717_and_in[1]), .A2(n426), .ZN(
        cell_1717_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1717_a_HPC2_and_U6 ( .A1(cell_1717_and_in[0]), .A2(n409), .ZN(
        cell_1717_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1717_a_HPC2_and_U5 ( .A(cell_1717_a_HPC2_and_n8), .B(
        cell_1717_a_HPC2_and_z_1__1_), .ZN(cell_1717_and_out[1]) );
  XNOR2_X1 cell_1717_a_HPC2_and_U4 ( .A(
        cell_1717_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1717_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1717_a_HPC2_and_n8) );
  XNOR2_X1 cell_1717_a_HPC2_and_U3 ( .A(cell_1717_a_HPC2_and_n7), .B(
        cell_1717_a_HPC2_and_z_0__0_), .ZN(cell_1717_and_out[0]) );
  XNOR2_X1 cell_1717_a_HPC2_and_U2 ( .A(
        cell_1717_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1717_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1717_a_HPC2_and_n7) );
  DFF_X1 cell_1717_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1717_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1717_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1717_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1717_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1717_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1717_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1717_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1717_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1717_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1718_U4 ( .A(1'b0), .B(cell_1718_and_out[1]), .Z(signal_3260)
         );
  XOR2_X1 cell_1718_U3 ( .A(1'b1), .B(cell_1718_and_out[0]), .Z(signal_1986)
         );
  XOR2_X1 cell_1718_U2 ( .A(1'b0), .B(1'b0), .Z(cell_1718_and_in[1]) );
  XOR2_X1 cell_1718_U1 ( .A(1'b1), .B(1'b0), .Z(cell_1718_and_in[0]) );
  XOR2_X1 cell_1718_a_HPC2_and_U14 ( .A(Fresh[4]), .B(cell_1718_and_in[0]), 
        .Z(cell_1718_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1718_a_HPC2_and_U13 ( .A(Fresh[4]), .B(cell_1718_and_in[1]), 
        .Z(cell_1718_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1718_a_HPC2_and_U12 ( .A1(cell_1718_a_HPC2_and_a_reg[1]), .A2(
        cell_1718_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1718_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1718_a_HPC2_and_U11 ( .A1(cell_1718_a_HPC2_and_a_reg[0]), .A2(
        cell_1718_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1718_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1718_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1718_a_HPC2_and_n9), 
        .ZN(cell_1718_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1718_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1718_a_HPC2_and_n9), 
        .ZN(cell_1718_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1718_a_HPC2_and_U8 ( .A(Fresh[4]), .ZN(cell_1718_a_HPC2_and_n9)
         );
  AND2_X1 cell_1718_a_HPC2_and_U7 ( .A1(cell_1718_and_in[1]), .A2(n426), .ZN(
        cell_1718_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1718_a_HPC2_and_U6 ( .A1(cell_1718_and_in[0]), .A2(n409), .ZN(
        cell_1718_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1718_a_HPC2_and_U5 ( .A(cell_1718_a_HPC2_and_n8), .B(
        cell_1718_a_HPC2_and_z_1__1_), .ZN(cell_1718_and_out[1]) );
  XNOR2_X1 cell_1718_a_HPC2_and_U4 ( .A(
        cell_1718_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1718_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1718_a_HPC2_and_n8) );
  XNOR2_X1 cell_1718_a_HPC2_and_U3 ( .A(cell_1718_a_HPC2_and_n7), .B(
        cell_1718_a_HPC2_and_z_0__0_), .ZN(cell_1718_and_out[0]) );
  XNOR2_X1 cell_1718_a_HPC2_and_U2 ( .A(
        cell_1718_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1718_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1718_a_HPC2_and_n7) );
  DFF_X1 cell_1718_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1718_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1718_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1718_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1718_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1718_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1718_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1718_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1718_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1718_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1719_U4 ( .A(1'b0), .B(1'b0), .Z(cell_1719_and_in[1]) );
  XOR2_X1 cell_1719_U3 ( .A(1'b0), .B(1'b1), .Z(cell_1719_and_in[0]) );
  XOR2_X1 cell_1719_U2 ( .A(1'b0), .B(cell_1719_and_out[0]), .Z(signal_1987)
         );
  XOR2_X1 cell_1719_U1 ( .A(1'b0), .B(cell_1719_and_out[1]), .Z(signal_3261)
         );
  XOR2_X1 cell_1719_a_HPC2_and_U14 ( .A(Fresh[5]), .B(cell_1719_and_in[0]), 
        .Z(cell_1719_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1719_a_HPC2_and_U13 ( .A(Fresh[5]), .B(cell_1719_and_in[1]), 
        .Z(cell_1719_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1719_a_HPC2_and_U12 ( .A1(cell_1719_a_HPC2_and_a_reg[1]), .A2(
        cell_1719_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1719_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1719_a_HPC2_and_U11 ( .A1(cell_1719_a_HPC2_and_a_reg[0]), .A2(
        cell_1719_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1719_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1719_a_HPC2_and_U10 ( .A1(signal_3232), .A2(
        cell_1719_a_HPC2_and_n9), .ZN(cell_1719_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1719_a_HPC2_and_U9 ( .A1(signal_1517), .A2(
        cell_1719_a_HPC2_and_n9), .ZN(cell_1719_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1719_a_HPC2_and_U8 ( .A(Fresh[5]), .ZN(cell_1719_a_HPC2_and_n9)
         );
  AND2_X1 cell_1719_a_HPC2_and_U7 ( .A1(cell_1719_and_in[1]), .A2(signal_3232), 
        .ZN(cell_1719_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1719_a_HPC2_and_U6 ( .A1(cell_1719_and_in[0]), .A2(signal_1517), 
        .ZN(cell_1719_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1719_a_HPC2_and_U5 ( .A(cell_1719_a_HPC2_and_n8), .B(
        cell_1719_a_HPC2_and_z_1__1_), .ZN(cell_1719_and_out[1]) );
  XNOR2_X1 cell_1719_a_HPC2_and_U4 ( .A(
        cell_1719_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1719_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1719_a_HPC2_and_n8) );
  XNOR2_X1 cell_1719_a_HPC2_and_U3 ( .A(cell_1719_a_HPC2_and_n7), .B(
        cell_1719_a_HPC2_and_z_0__0_), .ZN(cell_1719_and_out[0]) );
  XNOR2_X1 cell_1719_a_HPC2_and_U2 ( .A(
        cell_1719_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1719_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1719_a_HPC2_and_n7) );
  DFF_X1 cell_1719_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1719_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1719_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1517), 
        .CK(clk), .Q(cell_1719_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1719_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1719_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3232), 
        .CK(clk), .Q(cell_1719_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1719_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1719_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1719_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1720_U4 ( .A(1'b0), .B(cell_1720_and_out[1]), .Z(signal_3402)
         );
  XOR2_X1 cell_1720_U3 ( .A(1'b1), .B(cell_1720_and_out[0]), .Z(signal_1988)
         );
  XOR2_X1 cell_1720_U2 ( .A(1'b0), .B(n389), .Z(cell_1720_and_in[1]) );
  XOR2_X1 cell_1720_U1 ( .A(1'b1), .B(n388), .Z(cell_1720_and_in[0]) );
  XOR2_X1 cell_1720_a_HPC2_and_U14 ( .A(Fresh[6]), .B(cell_1720_and_in[0]), 
        .Z(cell_1720_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1720_a_HPC2_and_U13 ( .A(Fresh[6]), .B(cell_1720_and_in[1]), 
        .Z(cell_1720_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1720_a_HPC2_and_U12 ( .A1(cell_1720_a_HPC2_and_a_reg[1]), .A2(
        cell_1720_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1720_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1720_a_HPC2_and_U11 ( .A1(cell_1720_a_HPC2_and_a_reg[0]), .A2(
        cell_1720_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1720_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1720_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1720_a_HPC2_and_n9), 
        .ZN(cell_1720_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1720_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1720_a_HPC2_and_n9), 
        .ZN(cell_1720_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1720_a_HPC2_and_U8 ( .A(Fresh[6]), .ZN(cell_1720_a_HPC2_and_n9)
         );
  AND2_X1 cell_1720_a_HPC2_and_U7 ( .A1(cell_1720_and_in[1]), .A2(n426), .ZN(
        cell_1720_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1720_a_HPC2_and_U6 ( .A1(cell_1720_and_in[0]), .A2(n409), .ZN(
        cell_1720_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1720_a_HPC2_and_U5 ( .A(cell_1720_a_HPC2_and_n8), .B(
        cell_1720_a_HPC2_and_z_1__1_), .ZN(cell_1720_and_out[1]) );
  XNOR2_X1 cell_1720_a_HPC2_and_U4 ( .A(
        cell_1720_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1720_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1720_a_HPC2_and_n8) );
  XNOR2_X1 cell_1720_a_HPC2_and_U3 ( .A(cell_1720_a_HPC2_and_n7), .B(
        cell_1720_a_HPC2_and_z_0__0_), .ZN(cell_1720_and_out[0]) );
  XNOR2_X1 cell_1720_a_HPC2_and_U2 ( .A(
        cell_1720_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1720_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1720_a_HPC2_and_n7) );
  DFF_X1 cell_1720_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1720_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1720_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1720_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1720_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1720_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1720_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1720_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1720_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1720_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1721_U4 ( .A(n383), .B(cell_1721_and_out[1]), .Z(signal_3403)
         );
  XOR2_X1 cell_1721_U3 ( .A(n382), .B(cell_1721_and_out[0]), .Z(signal_1989)
         );
  XOR2_X1 cell_1721_U2 ( .A(n383), .B(signal_3256), .Z(cell_1721_and_in[1]) );
  XOR2_X1 cell_1721_U1 ( .A(n382), .B(signal_1982), .Z(cell_1721_and_in[0]) );
  XOR2_X1 cell_1721_a_HPC2_and_U14 ( .A(Fresh[7]), .B(cell_1721_and_in[0]), 
        .Z(cell_1721_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1721_a_HPC2_and_U13 ( .A(Fresh[7]), .B(cell_1721_and_in[1]), 
        .Z(cell_1721_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1721_a_HPC2_and_U12 ( .A1(cell_1721_a_HPC2_and_a_reg[1]), .A2(
        cell_1721_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1721_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1721_a_HPC2_and_U11 ( .A1(cell_1721_a_HPC2_and_a_reg[0]), .A2(
        cell_1721_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1721_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1721_a_HPC2_and_U10 ( .A1(signal_3237), .A2(
        cell_1721_a_HPC2_and_n9), .ZN(cell_1721_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1721_a_HPC2_and_U9 ( .A1(signal_1512), .A2(
        cell_1721_a_HPC2_and_n9), .ZN(cell_1721_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1721_a_HPC2_and_U8 ( .A(Fresh[7]), .ZN(cell_1721_a_HPC2_and_n9)
         );
  AND2_X1 cell_1721_a_HPC2_and_U7 ( .A1(cell_1721_and_in[1]), .A2(signal_3237), 
        .ZN(cell_1721_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1721_a_HPC2_and_U6 ( .A1(cell_1721_and_in[0]), .A2(signal_1512), 
        .ZN(cell_1721_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1721_a_HPC2_and_U5 ( .A(cell_1721_a_HPC2_and_n8), .B(
        cell_1721_a_HPC2_and_z_1__1_), .ZN(cell_1721_and_out[1]) );
  XNOR2_X1 cell_1721_a_HPC2_and_U4 ( .A(
        cell_1721_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1721_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1721_a_HPC2_and_n8) );
  XNOR2_X1 cell_1721_a_HPC2_and_U3 ( .A(cell_1721_a_HPC2_and_n7), .B(
        cell_1721_a_HPC2_and_z_0__0_), .ZN(cell_1721_and_out[0]) );
  XNOR2_X1 cell_1721_a_HPC2_and_U2 ( .A(
        cell_1721_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1721_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1721_a_HPC2_and_n7) );
  DFF_X1 cell_1721_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1721_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1721_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1512), 
        .CK(clk), .Q(cell_1721_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1721_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1721_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3237), 
        .CK(clk), .Q(cell_1721_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1721_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1721_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1721_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1722_U4 ( .A(n389), .B(cell_1722_and_out[1]), .Z(signal_3404)
         );
  XOR2_X1 cell_1722_U3 ( .A(n388), .B(cell_1722_and_out[0]), .Z(signal_1990)
         );
  XOR2_X1 cell_1722_U2 ( .A(n389), .B(n387), .Z(cell_1722_and_in[1]) );
  XOR2_X1 cell_1722_U1 ( .A(n388), .B(n385), .Z(cell_1722_and_in[0]) );
  XOR2_X1 cell_1722_a_HPC2_and_U14 ( .A(Fresh[8]), .B(cell_1722_and_in[0]), 
        .Z(cell_1722_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1722_a_HPC2_and_U13 ( .A(Fresh[8]), .B(cell_1722_and_in[1]), 
        .Z(cell_1722_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1722_a_HPC2_and_U12 ( .A1(cell_1722_a_HPC2_and_a_reg[1]), .A2(
        cell_1722_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1722_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1722_a_HPC2_and_U11 ( .A1(cell_1722_a_HPC2_and_a_reg[0]), .A2(
        cell_1722_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1722_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1722_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1722_a_HPC2_and_n9), 
        .ZN(cell_1722_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1722_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1722_a_HPC2_and_n9), 
        .ZN(cell_1722_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1722_a_HPC2_and_U8 ( .A(Fresh[8]), .ZN(cell_1722_a_HPC2_and_n9)
         );
  AND2_X1 cell_1722_a_HPC2_and_U7 ( .A1(cell_1722_and_in[1]), .A2(n411), .ZN(
        cell_1722_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1722_a_HPC2_and_U6 ( .A1(cell_1722_and_in[0]), .A2(n394), .ZN(
        cell_1722_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1722_a_HPC2_and_U5 ( .A(cell_1722_a_HPC2_and_n8), .B(
        cell_1722_a_HPC2_and_z_1__1_), .ZN(cell_1722_and_out[1]) );
  XNOR2_X1 cell_1722_a_HPC2_and_U4 ( .A(
        cell_1722_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1722_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1722_a_HPC2_and_n8) );
  XNOR2_X1 cell_1722_a_HPC2_and_U3 ( .A(cell_1722_a_HPC2_and_n7), .B(
        cell_1722_a_HPC2_and_z_0__0_), .ZN(cell_1722_and_out[0]) );
  XNOR2_X1 cell_1722_a_HPC2_and_U2 ( .A(
        cell_1722_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1722_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1722_a_HPC2_and_n7) );
  DFF_X1 cell_1722_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1722_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1722_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1722_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1722_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1722_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1722_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1722_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1722_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1722_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1723_U4 ( .A(n383), .B(cell_1723_and_out[1]), .Z(signal_3405)
         );
  XOR2_X1 cell_1723_U3 ( .A(n382), .B(cell_1723_and_out[0]), .Z(signal_1991)
         );
  XOR2_X1 cell_1723_U2 ( .A(n383), .B(n387), .Z(cell_1723_and_in[1]) );
  XOR2_X1 cell_1723_U1 ( .A(n382), .B(n385), .Z(cell_1723_and_in[0]) );
  XOR2_X1 cell_1723_a_HPC2_and_U14 ( .A(Fresh[9]), .B(cell_1723_and_in[0]), 
        .Z(cell_1723_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1723_a_HPC2_and_U13 ( .A(Fresh[9]), .B(cell_1723_and_in[1]), 
        .Z(cell_1723_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1723_a_HPC2_and_U12 ( .A1(cell_1723_a_HPC2_and_a_reg[1]), .A2(
        cell_1723_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1723_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1723_a_HPC2_and_U11 ( .A1(cell_1723_a_HPC2_and_a_reg[0]), .A2(
        cell_1723_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1723_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1723_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1723_a_HPC2_and_n9), 
        .ZN(cell_1723_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1723_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1723_a_HPC2_and_n9), 
        .ZN(cell_1723_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1723_a_HPC2_and_U8 ( .A(Fresh[9]), .ZN(cell_1723_a_HPC2_and_n9)
         );
  AND2_X1 cell_1723_a_HPC2_and_U7 ( .A1(cell_1723_and_in[1]), .A2(n411), .ZN(
        cell_1723_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1723_a_HPC2_and_U6 ( .A1(cell_1723_and_in[0]), .A2(n394), .ZN(
        cell_1723_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1723_a_HPC2_and_U5 ( .A(cell_1723_a_HPC2_and_n8), .B(
        cell_1723_a_HPC2_and_z_1__1_), .ZN(cell_1723_and_out[1]) );
  XNOR2_X1 cell_1723_a_HPC2_and_U4 ( .A(
        cell_1723_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1723_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1723_a_HPC2_and_n8) );
  XNOR2_X1 cell_1723_a_HPC2_and_U3 ( .A(cell_1723_a_HPC2_and_n7), .B(
        cell_1723_a_HPC2_and_z_0__0_), .ZN(cell_1723_and_out[0]) );
  XNOR2_X1 cell_1723_a_HPC2_and_U2 ( .A(
        cell_1723_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1723_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1723_a_HPC2_and_n7) );
  DFF_X1 cell_1723_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1723_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1723_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1723_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1723_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1723_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1723_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1723_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1723_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1723_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1724_U6 ( .A(n389), .B(1'b0), .Z(cell_1724_and_in[1]) );
  XOR2_X1 cell_1724_U5 ( .A(n388), .B(1'b1), .Z(cell_1724_and_in[0]) );
  XOR2_X1 cell_1724_U4 ( .A(n389), .B(cell_1724_and_out[1]), .Z(cell_1724_n5)
         );
  BUF_X2 cell_1724_U3 ( .A(cell_1724_n5), .Z(signal_3406) );
  XOR2_X1 cell_1724_U2 ( .A(n388), .B(cell_1724_and_out[0]), .Z(cell_1724_n6)
         );
  BUF_X2 cell_1724_U1 ( .A(cell_1724_n6), .Z(signal_1992) );
  XOR2_X1 cell_1724_a_HPC2_and_U14 ( .A(Fresh[10]), .B(cell_1724_and_in[0]), 
        .Z(cell_1724_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1724_a_HPC2_and_U13 ( .A(Fresh[10]), .B(cell_1724_and_in[1]), 
        .Z(cell_1724_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1724_a_HPC2_and_U12 ( .A1(cell_1724_a_HPC2_and_a_reg[1]), .A2(
        cell_1724_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1724_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1724_a_HPC2_and_U11 ( .A1(cell_1724_a_HPC2_and_a_reg[0]), .A2(
        cell_1724_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1724_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1724_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1724_a_HPC2_and_n9), 
        .ZN(cell_1724_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1724_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1724_a_HPC2_and_n9), 
        .ZN(cell_1724_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1724_a_HPC2_and_U8 ( .A(Fresh[10]), .ZN(cell_1724_a_HPC2_and_n9)
         );
  AND2_X1 cell_1724_a_HPC2_and_U7 ( .A1(cell_1724_and_in[1]), .A2(n393), .ZN(
        cell_1724_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1724_a_HPC2_and_U6 ( .A1(cell_1724_and_in[0]), .A2(n392), .ZN(
        cell_1724_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1724_a_HPC2_and_U5 ( .A(cell_1724_a_HPC2_and_n8), .B(
        cell_1724_a_HPC2_and_z_1__1_), .ZN(cell_1724_and_out[1]) );
  XNOR2_X1 cell_1724_a_HPC2_and_U4 ( .A(
        cell_1724_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1724_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1724_a_HPC2_and_n8) );
  XNOR2_X1 cell_1724_a_HPC2_and_U3 ( .A(cell_1724_a_HPC2_and_n7), .B(
        cell_1724_a_HPC2_and_z_0__0_), .ZN(cell_1724_and_out[0]) );
  XNOR2_X1 cell_1724_a_HPC2_and_U2 ( .A(
        cell_1724_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1724_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1724_a_HPC2_and_n7) );
  DFF_X1 cell_1724_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1724_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1724_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1724_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1724_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1724_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1724_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1724_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1724_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1724_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1725_U4 ( .A(1'b0), .B(n389), .Z(cell_1725_and_in[1]) );
  XOR2_X1 cell_1725_U3 ( .A(1'b1), .B(n388), .Z(cell_1725_and_in[0]) );
  XOR2_X1 cell_1725_U2 ( .A(1'b0), .B(cell_1725_and_out[1]), .Z(signal_3407)
         );
  XOR2_X1 cell_1725_U1 ( .A(1'b1), .B(cell_1725_and_out[0]), .Z(signal_1993)
         );
  XOR2_X1 cell_1725_a_HPC2_and_U14 ( .A(Fresh[11]), .B(cell_1725_and_in[0]), 
        .Z(cell_1725_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1725_a_HPC2_and_U13 ( .A(Fresh[11]), .B(cell_1725_and_in[1]), 
        .Z(cell_1725_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1725_a_HPC2_and_U12 ( .A1(cell_1725_a_HPC2_and_a_reg[1]), .A2(
        cell_1725_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1725_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1725_a_HPC2_and_U11 ( .A1(cell_1725_a_HPC2_and_a_reg[0]), .A2(
        cell_1725_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1725_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1725_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1725_a_HPC2_and_n9), 
        .ZN(cell_1725_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1725_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1725_a_HPC2_and_n9), 
        .ZN(cell_1725_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1725_a_HPC2_and_U8 ( .A(Fresh[11]), .ZN(cell_1725_a_HPC2_and_n9)
         );
  AND2_X1 cell_1725_a_HPC2_and_U7 ( .A1(cell_1725_and_in[1]), .A2(n393), .ZN(
        cell_1725_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1725_a_HPC2_and_U6 ( .A1(cell_1725_and_in[0]), .A2(n392), .ZN(
        cell_1725_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1725_a_HPC2_and_U5 ( .A(cell_1725_a_HPC2_and_n8), .B(
        cell_1725_a_HPC2_and_z_1__1_), .ZN(cell_1725_and_out[1]) );
  XNOR2_X1 cell_1725_a_HPC2_and_U4 ( .A(
        cell_1725_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1725_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1725_a_HPC2_and_n8) );
  XNOR2_X1 cell_1725_a_HPC2_and_U3 ( .A(cell_1725_a_HPC2_and_n7), .B(
        cell_1725_a_HPC2_and_z_0__0_), .ZN(cell_1725_and_out[0]) );
  XNOR2_X1 cell_1725_a_HPC2_and_U2 ( .A(
        cell_1725_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1725_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1725_a_HPC2_and_n7) );
  DFF_X1 cell_1725_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1725_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1725_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1725_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1725_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1725_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1725_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1725_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1725_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1725_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1726_U4 ( .A(1'b0), .B(cell_1726_and_out[1]), .Z(signal_3408)
         );
  XOR2_X1 cell_1726_U3 ( .A(1'b0), .B(cell_1726_and_out[0]), .Z(signal_1994)
         );
  XOR2_X1 cell_1726_U2 ( .A(1'b0), .B(n387), .Z(cell_1726_and_in[1]) );
  XOR2_X1 cell_1726_U1 ( .A(1'b0), .B(n385), .Z(cell_1726_and_in[0]) );
  XOR2_X1 cell_1726_a_HPC2_and_U14 ( .A(Fresh[12]), .B(cell_1726_and_in[0]), 
        .Z(cell_1726_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1726_a_HPC2_and_U13 ( .A(Fresh[12]), .B(cell_1726_and_in[1]), 
        .Z(cell_1726_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1726_a_HPC2_and_U12 ( .A1(cell_1726_a_HPC2_and_a_reg[1]), .A2(
        cell_1726_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1726_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1726_a_HPC2_and_U11 ( .A1(cell_1726_a_HPC2_and_a_reg[0]), .A2(
        cell_1726_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1726_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1726_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1726_a_HPC2_and_n9), 
        .ZN(cell_1726_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1726_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1726_a_HPC2_and_n9), 
        .ZN(cell_1726_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1726_a_HPC2_and_U8 ( .A(Fresh[12]), .ZN(cell_1726_a_HPC2_and_n9)
         );
  AND2_X1 cell_1726_a_HPC2_and_U7 ( .A1(cell_1726_and_in[1]), .A2(n426), .ZN(
        cell_1726_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1726_a_HPC2_and_U6 ( .A1(cell_1726_and_in[0]), .A2(n409), .ZN(
        cell_1726_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1726_a_HPC2_and_U5 ( .A(cell_1726_a_HPC2_and_n8), .B(
        cell_1726_a_HPC2_and_z_1__1_), .ZN(cell_1726_and_out[1]) );
  XNOR2_X1 cell_1726_a_HPC2_and_U4 ( .A(
        cell_1726_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1726_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1726_a_HPC2_and_n8) );
  XNOR2_X1 cell_1726_a_HPC2_and_U3 ( .A(cell_1726_a_HPC2_and_n7), .B(
        cell_1726_a_HPC2_and_z_0__0_), .ZN(cell_1726_and_out[0]) );
  XNOR2_X1 cell_1726_a_HPC2_and_U2 ( .A(
        cell_1726_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1726_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1726_a_HPC2_and_n7) );
  DFF_X1 cell_1726_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1726_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1726_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1726_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1726_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1726_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1726_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1726_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1726_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1726_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1727_U4 ( .A(n389), .B(cell_1727_and_out[1]), .Z(signal_3409)
         );
  XOR2_X1 cell_1727_U3 ( .A(n388), .B(cell_1727_and_out[0]), .Z(signal_1995)
         );
  XOR2_X1 cell_1727_U2 ( .A(n389), .B(1'b0), .Z(cell_1727_and_in[1]) );
  XOR2_X1 cell_1727_U1 ( .A(n388), .B(1'b0), .Z(cell_1727_and_in[0]) );
  XOR2_X1 cell_1727_a_HPC2_and_U14 ( .A(Fresh[13]), .B(cell_1727_and_in[0]), 
        .Z(cell_1727_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1727_a_HPC2_and_U13 ( .A(Fresh[13]), .B(cell_1727_and_in[1]), 
        .Z(cell_1727_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1727_a_HPC2_and_U12 ( .A1(cell_1727_a_HPC2_and_a_reg[1]), .A2(
        cell_1727_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1727_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1727_a_HPC2_and_U11 ( .A1(cell_1727_a_HPC2_and_a_reg[0]), .A2(
        cell_1727_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1727_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1727_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1727_a_HPC2_and_n9), 
        .ZN(cell_1727_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1727_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1727_a_HPC2_and_n9), 
        .ZN(cell_1727_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1727_a_HPC2_and_U8 ( .A(Fresh[13]), .ZN(cell_1727_a_HPC2_and_n9)
         );
  AND2_X1 cell_1727_a_HPC2_and_U7 ( .A1(cell_1727_and_in[1]), .A2(n426), .ZN(
        cell_1727_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1727_a_HPC2_and_U6 ( .A1(cell_1727_and_in[0]), .A2(n409), .ZN(
        cell_1727_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1727_a_HPC2_and_U5 ( .A(cell_1727_a_HPC2_and_n8), .B(
        cell_1727_a_HPC2_and_z_1__1_), .ZN(cell_1727_and_out[1]) );
  XNOR2_X1 cell_1727_a_HPC2_and_U4 ( .A(
        cell_1727_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1727_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1727_a_HPC2_and_n8) );
  XNOR2_X1 cell_1727_a_HPC2_and_U3 ( .A(cell_1727_a_HPC2_and_n7), .B(
        cell_1727_a_HPC2_and_z_0__0_), .ZN(cell_1727_and_out[0]) );
  XNOR2_X1 cell_1727_a_HPC2_and_U2 ( .A(
        cell_1727_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1727_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1727_a_HPC2_and_n7) );
  DFF_X1 cell_1727_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1727_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1727_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1727_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1727_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1727_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1727_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1727_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1727_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1727_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1728_U4 ( .A(n381), .B(cell_1728_and_out[1]), .Z(signal_3410)
         );
  XOR2_X1 cell_1728_U3 ( .A(n380), .B(cell_1728_and_out[0]), .Z(signal_1996)
         );
  XOR2_X1 cell_1728_U2 ( .A(n381), .B(signal_3256), .Z(cell_1728_and_in[1]) );
  XOR2_X1 cell_1728_U1 ( .A(n380), .B(signal_1982), .Z(cell_1728_and_in[0]) );
  XOR2_X1 cell_1728_a_HPC2_and_U14 ( .A(Fresh[14]), .B(cell_1728_and_in[0]), 
        .Z(cell_1728_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1728_a_HPC2_and_U13 ( .A(Fresh[14]), .B(cell_1728_and_in[1]), 
        .Z(cell_1728_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1728_a_HPC2_and_U12 ( .A1(cell_1728_a_HPC2_and_a_reg[1]), .A2(
        cell_1728_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1728_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1728_a_HPC2_and_U11 ( .A1(cell_1728_a_HPC2_and_a_reg[0]), .A2(
        cell_1728_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1728_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1728_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1728_a_HPC2_and_n9), 
        .ZN(cell_1728_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1728_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1728_a_HPC2_and_n9), 
        .ZN(cell_1728_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1728_a_HPC2_and_U8 ( .A(Fresh[14]), .ZN(cell_1728_a_HPC2_and_n9)
         );
  AND2_X1 cell_1728_a_HPC2_and_U7 ( .A1(cell_1728_and_in[1]), .A2(n393), .ZN(
        cell_1728_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1728_a_HPC2_and_U6 ( .A1(cell_1728_and_in[0]), .A2(n392), .ZN(
        cell_1728_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1728_a_HPC2_and_U5 ( .A(cell_1728_a_HPC2_and_n8), .B(
        cell_1728_a_HPC2_and_z_1__1_), .ZN(cell_1728_and_out[1]) );
  XNOR2_X1 cell_1728_a_HPC2_and_U4 ( .A(
        cell_1728_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1728_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1728_a_HPC2_and_n8) );
  XNOR2_X1 cell_1728_a_HPC2_and_U3 ( .A(cell_1728_a_HPC2_and_n7), .B(
        cell_1728_a_HPC2_and_z_0__0_), .ZN(cell_1728_and_out[0]) );
  XNOR2_X1 cell_1728_a_HPC2_and_U2 ( .A(
        cell_1728_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1728_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1728_a_HPC2_and_n7) );
  DFF_X1 cell_1728_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1728_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1728_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1728_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1728_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1728_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1728_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1728_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1728_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1728_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1729_U4 ( .A(1'b0), .B(cell_1729_and_out[1]), .Z(signal_3411)
         );
  XOR2_X1 cell_1729_U3 ( .A(1'b0), .B(cell_1729_and_out[0]), .Z(signal_1997)
         );
  XOR2_X1 cell_1729_U2 ( .A(1'b0), .B(n389), .Z(cell_1729_and_in[1]) );
  XOR2_X1 cell_1729_U1 ( .A(1'b0), .B(n388), .Z(cell_1729_and_in[0]) );
  XOR2_X1 cell_1729_a_HPC2_and_U14 ( .A(Fresh[15]), .B(cell_1729_and_in[0]), 
        .Z(cell_1729_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1729_a_HPC2_and_U13 ( .A(Fresh[15]), .B(cell_1729_and_in[1]), 
        .Z(cell_1729_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1729_a_HPC2_and_U12 ( .A1(cell_1729_a_HPC2_and_a_reg[1]), .A2(
        cell_1729_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1729_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1729_a_HPC2_and_U11 ( .A1(cell_1729_a_HPC2_and_a_reg[0]), .A2(
        cell_1729_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1729_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1729_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1729_a_HPC2_and_n9), 
        .ZN(cell_1729_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1729_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1729_a_HPC2_and_n9), 
        .ZN(cell_1729_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1729_a_HPC2_and_U8 ( .A(Fresh[15]), .ZN(cell_1729_a_HPC2_and_n9)
         );
  AND2_X1 cell_1729_a_HPC2_and_U7 ( .A1(cell_1729_and_in[1]), .A2(n393), .ZN(
        cell_1729_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1729_a_HPC2_and_U6 ( .A1(cell_1729_and_in[0]), .A2(n392), .ZN(
        cell_1729_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1729_a_HPC2_and_U5 ( .A(cell_1729_a_HPC2_and_n8), .B(
        cell_1729_a_HPC2_and_z_1__1_), .ZN(cell_1729_and_out[1]) );
  XNOR2_X1 cell_1729_a_HPC2_and_U4 ( .A(
        cell_1729_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1729_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1729_a_HPC2_and_n8) );
  XNOR2_X1 cell_1729_a_HPC2_and_U3 ( .A(cell_1729_a_HPC2_and_n7), .B(
        cell_1729_a_HPC2_and_z_0__0_), .ZN(cell_1729_and_out[0]) );
  XNOR2_X1 cell_1729_a_HPC2_and_U2 ( .A(
        cell_1729_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1729_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1729_a_HPC2_and_n7) );
  DFF_X1 cell_1729_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1729_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1729_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1729_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1729_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1729_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1729_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1729_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1729_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1729_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1730_U4 ( .A(1'b0), .B(cell_1730_and_out[1]), .Z(signal_3412)
         );
  XOR2_X1 cell_1730_U3 ( .A(1'b1), .B(cell_1730_and_out[0]), .Z(signal_1998)
         );
  XOR2_X1 cell_1730_U2 ( .A(1'b0), .B(n383), .Z(cell_1730_and_in[1]) );
  XOR2_X1 cell_1730_U1 ( .A(1'b1), .B(n382), .Z(cell_1730_and_in[0]) );
  XOR2_X1 cell_1730_a_HPC2_and_U14 ( .A(Fresh[16]), .B(cell_1730_and_in[0]), 
        .Z(cell_1730_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1730_a_HPC2_and_U13 ( .A(Fresh[16]), .B(cell_1730_and_in[1]), 
        .Z(cell_1730_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1730_a_HPC2_and_U12 ( .A1(cell_1730_a_HPC2_and_a_reg[1]), .A2(
        cell_1730_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1730_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1730_a_HPC2_and_U11 ( .A1(cell_1730_a_HPC2_and_a_reg[0]), .A2(
        cell_1730_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1730_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1730_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1730_a_HPC2_and_n9), 
        .ZN(cell_1730_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1730_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1730_a_HPC2_and_n9), 
        .ZN(cell_1730_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1730_a_HPC2_and_U8 ( .A(Fresh[16]), .ZN(cell_1730_a_HPC2_and_n9)
         );
  AND2_X1 cell_1730_a_HPC2_and_U7 ( .A1(cell_1730_and_in[1]), .A2(n427), .ZN(
        cell_1730_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1730_a_HPC2_and_U6 ( .A1(cell_1730_and_in[0]), .A2(n410), .ZN(
        cell_1730_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1730_a_HPC2_and_U5 ( .A(cell_1730_a_HPC2_and_n8), .B(
        cell_1730_a_HPC2_and_z_1__1_), .ZN(cell_1730_and_out[1]) );
  XNOR2_X1 cell_1730_a_HPC2_and_U4 ( .A(
        cell_1730_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1730_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1730_a_HPC2_and_n8) );
  XNOR2_X1 cell_1730_a_HPC2_and_U3 ( .A(cell_1730_a_HPC2_and_n7), .B(
        cell_1730_a_HPC2_and_z_0__0_), .ZN(cell_1730_and_out[0]) );
  XNOR2_X1 cell_1730_a_HPC2_and_U2 ( .A(
        cell_1730_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1730_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1730_a_HPC2_and_n7) );
  DFF_X1 cell_1730_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1730_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1730_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1730_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1730_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1730_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1730_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1730_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1730_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1730_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1731_U4 ( .A(1'b0), .B(n381), .Z(cell_1731_and_in[1]) );
  XOR2_X1 cell_1731_U3 ( .A(1'b1), .B(n380), .Z(cell_1731_and_in[0]) );
  XOR2_X1 cell_1731_U2 ( .A(1'b1), .B(cell_1731_and_out[0]), .Z(signal_1999)
         );
  XOR2_X1 cell_1731_U1 ( .A(1'b0), .B(cell_1731_and_out[1]), .Z(signal_3413)
         );
  XOR2_X1 cell_1731_a_HPC2_and_U14 ( .A(Fresh[17]), .B(cell_1731_and_in[0]), 
        .Z(cell_1731_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1731_a_HPC2_and_U13 ( .A(Fresh[17]), .B(cell_1731_and_in[1]), 
        .Z(cell_1731_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1731_a_HPC2_and_U12 ( .A1(cell_1731_a_HPC2_and_a_reg[1]), .A2(
        cell_1731_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1731_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1731_a_HPC2_and_U11 ( .A1(cell_1731_a_HPC2_and_a_reg[0]), .A2(
        cell_1731_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1731_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1731_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1731_a_HPC2_and_n9), 
        .ZN(cell_1731_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1731_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1731_a_HPC2_and_n9), 
        .ZN(cell_1731_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1731_a_HPC2_and_U8 ( .A(Fresh[17]), .ZN(cell_1731_a_HPC2_and_n9)
         );
  AND2_X1 cell_1731_a_HPC2_and_U7 ( .A1(cell_1731_and_in[1]), .A2(n393), .ZN(
        cell_1731_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1731_a_HPC2_and_U6 ( .A1(cell_1731_and_in[0]), .A2(n392), .ZN(
        cell_1731_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1731_a_HPC2_and_U5 ( .A(cell_1731_a_HPC2_and_n8), .B(
        cell_1731_a_HPC2_and_z_1__1_), .ZN(cell_1731_and_out[1]) );
  XNOR2_X1 cell_1731_a_HPC2_and_U4 ( .A(
        cell_1731_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1731_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1731_a_HPC2_and_n8) );
  XNOR2_X1 cell_1731_a_HPC2_and_U3 ( .A(cell_1731_a_HPC2_and_n7), .B(
        cell_1731_a_HPC2_and_z_0__0_), .ZN(cell_1731_and_out[0]) );
  XNOR2_X1 cell_1731_a_HPC2_and_U2 ( .A(
        cell_1731_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1731_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1731_a_HPC2_and_n7) );
  DFF_X1 cell_1731_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1731_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1731_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1731_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1731_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1731_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1731_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1731_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1731_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1731_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1732_U4 ( .A(1'b0), .B(cell_1732_and_out[1]), .Z(signal_3414)
         );
  XOR2_X1 cell_1732_U3 ( .A(1'b0), .B(cell_1732_and_out[0]), .Z(signal_2000)
         );
  XOR2_X1 cell_1732_U2 ( .A(1'b0), .B(n381), .Z(cell_1732_and_in[1]) );
  XOR2_X1 cell_1732_U1 ( .A(1'b0), .B(n380), .Z(cell_1732_and_in[0]) );
  XOR2_X1 cell_1732_a_HPC2_and_U14 ( .A(Fresh[18]), .B(cell_1732_and_in[0]), 
        .Z(cell_1732_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1732_a_HPC2_and_U13 ( .A(Fresh[18]), .B(cell_1732_and_in[1]), 
        .Z(cell_1732_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1732_a_HPC2_and_U12 ( .A1(cell_1732_a_HPC2_and_a_reg[1]), .A2(
        cell_1732_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1732_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1732_a_HPC2_and_U11 ( .A1(cell_1732_a_HPC2_and_a_reg[0]), .A2(
        cell_1732_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1732_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1732_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1732_a_HPC2_and_n9), 
        .ZN(cell_1732_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1732_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1732_a_HPC2_and_n9), 
        .ZN(cell_1732_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1732_a_HPC2_and_U8 ( .A(Fresh[18]), .ZN(cell_1732_a_HPC2_and_n9)
         );
  AND2_X1 cell_1732_a_HPC2_and_U7 ( .A1(cell_1732_and_in[1]), .A2(n393), .ZN(
        cell_1732_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1732_a_HPC2_and_U6 ( .A1(cell_1732_and_in[0]), .A2(n392), .ZN(
        cell_1732_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1732_a_HPC2_and_U5 ( .A(cell_1732_a_HPC2_and_n8), .B(
        cell_1732_a_HPC2_and_z_1__1_), .ZN(cell_1732_and_out[1]) );
  XNOR2_X1 cell_1732_a_HPC2_and_U4 ( .A(
        cell_1732_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1732_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1732_a_HPC2_and_n8) );
  XNOR2_X1 cell_1732_a_HPC2_and_U3 ( .A(cell_1732_a_HPC2_and_n7), .B(
        cell_1732_a_HPC2_and_z_0__0_), .ZN(cell_1732_and_out[0]) );
  XNOR2_X1 cell_1732_a_HPC2_and_U2 ( .A(
        cell_1732_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1732_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1732_a_HPC2_and_n7) );
  DFF_X1 cell_1732_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1732_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1732_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1732_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1732_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1732_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1732_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1732_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1732_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1732_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1733_U4 ( .A(n389), .B(cell_1733_and_out[1]), .Z(signal_3415)
         );
  XOR2_X1 cell_1733_U3 ( .A(n388), .B(cell_1733_and_out[0]), .Z(signal_2001)
         );
  XOR2_X1 cell_1733_U2 ( .A(n389), .B(n383), .Z(cell_1733_and_in[1]) );
  XOR2_X1 cell_1733_U1 ( .A(n388), .B(n382), .Z(cell_1733_and_in[0]) );
  XOR2_X1 cell_1733_a_HPC2_and_U14 ( .A(Fresh[19]), .B(cell_1733_and_in[0]), 
        .Z(cell_1733_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1733_a_HPC2_and_U13 ( .A(Fresh[19]), .B(cell_1733_and_in[1]), 
        .Z(cell_1733_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1733_a_HPC2_and_U12 ( .A1(cell_1733_a_HPC2_and_a_reg[1]), .A2(
        cell_1733_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1733_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1733_a_HPC2_and_U11 ( .A1(cell_1733_a_HPC2_and_a_reg[0]), .A2(
        cell_1733_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1733_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1733_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1733_a_HPC2_and_n9), 
        .ZN(cell_1733_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1733_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1733_a_HPC2_and_n9), 
        .ZN(cell_1733_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1733_a_HPC2_and_U8 ( .A(Fresh[19]), .ZN(cell_1733_a_HPC2_and_n9)
         );
  AND2_X1 cell_1733_a_HPC2_and_U7 ( .A1(cell_1733_and_in[1]), .A2(n411), .ZN(
        cell_1733_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1733_a_HPC2_and_U6 ( .A1(cell_1733_and_in[0]), .A2(n394), .ZN(
        cell_1733_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1733_a_HPC2_and_U5 ( .A(cell_1733_a_HPC2_and_n8), .B(
        cell_1733_a_HPC2_and_z_1__1_), .ZN(cell_1733_and_out[1]) );
  XNOR2_X1 cell_1733_a_HPC2_and_U4 ( .A(
        cell_1733_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1733_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1733_a_HPC2_and_n8) );
  XNOR2_X1 cell_1733_a_HPC2_and_U3 ( .A(cell_1733_a_HPC2_and_n7), .B(
        cell_1733_a_HPC2_and_z_0__0_), .ZN(cell_1733_and_out[0]) );
  XNOR2_X1 cell_1733_a_HPC2_and_U2 ( .A(
        cell_1733_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1733_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1733_a_HPC2_and_n7) );
  DFF_X1 cell_1733_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1733_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1733_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1733_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1733_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1733_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1733_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1733_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1733_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1733_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1734_U4 ( .A(n381), .B(cell_1734_and_out[1]), .Z(signal_3416)
         );
  XOR2_X1 cell_1734_U3 ( .A(n380), .B(cell_1734_and_out[0]), .Z(signal_2002)
         );
  XOR2_X1 cell_1734_U2 ( .A(n381), .B(signal_3258), .Z(cell_1734_and_in[1]) );
  XOR2_X1 cell_1734_U1 ( .A(n380), .B(signal_1984), .Z(cell_1734_and_in[0]) );
  XOR2_X1 cell_1734_a_HPC2_and_U14 ( .A(Fresh[20]), .B(cell_1734_and_in[0]), 
        .Z(cell_1734_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1734_a_HPC2_and_U13 ( .A(Fresh[20]), .B(cell_1734_and_in[1]), 
        .Z(cell_1734_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1734_a_HPC2_and_U12 ( .A1(cell_1734_a_HPC2_and_a_reg[1]), .A2(
        cell_1734_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1734_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1734_a_HPC2_and_U11 ( .A1(cell_1734_a_HPC2_and_a_reg[0]), .A2(
        cell_1734_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1734_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1734_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1734_a_HPC2_and_n9), 
        .ZN(cell_1734_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1734_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1734_a_HPC2_and_n9), 
        .ZN(cell_1734_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1734_a_HPC2_and_U8 ( .A(Fresh[20]), .ZN(cell_1734_a_HPC2_and_n9)
         );
  AND2_X1 cell_1734_a_HPC2_and_U7 ( .A1(cell_1734_and_in[1]), .A2(n411), .ZN(
        cell_1734_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1734_a_HPC2_and_U6 ( .A1(cell_1734_and_in[0]), .A2(n394), .ZN(
        cell_1734_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1734_a_HPC2_and_U5 ( .A(cell_1734_a_HPC2_and_n8), .B(
        cell_1734_a_HPC2_and_z_1__1_), .ZN(cell_1734_and_out[1]) );
  XNOR2_X1 cell_1734_a_HPC2_and_U4 ( .A(
        cell_1734_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1734_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1734_a_HPC2_and_n8) );
  XNOR2_X1 cell_1734_a_HPC2_and_U3 ( .A(cell_1734_a_HPC2_and_n7), .B(
        cell_1734_a_HPC2_and_z_0__0_), .ZN(cell_1734_and_out[0]) );
  XNOR2_X1 cell_1734_a_HPC2_and_U2 ( .A(
        cell_1734_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1734_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1734_a_HPC2_and_n7) );
  DFF_X1 cell_1734_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1734_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1734_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1734_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1734_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1734_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1734_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1734_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1734_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1734_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1735_U4 ( .A(1'b0), .B(cell_1735_and_out[1]), .Z(signal_3417)
         );
  XOR2_X1 cell_1735_U3 ( .A(1'b0), .B(cell_1735_and_out[0]), .Z(signal_2003)
         );
  XOR2_X1 cell_1735_U2 ( .A(1'b0), .B(n389), .Z(cell_1735_and_in[1]) );
  XOR2_X1 cell_1735_U1 ( .A(1'b0), .B(n388), .Z(cell_1735_and_in[0]) );
  XOR2_X1 cell_1735_a_HPC2_and_U14 ( .A(Fresh[21]), .B(cell_1735_and_in[0]), 
        .Z(cell_1735_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1735_a_HPC2_and_U13 ( .A(Fresh[21]), .B(cell_1735_and_in[1]), 
        .Z(cell_1735_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1735_a_HPC2_and_U12 ( .A1(cell_1735_a_HPC2_and_a_reg[1]), .A2(
        cell_1735_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1735_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1735_a_HPC2_and_U11 ( .A1(cell_1735_a_HPC2_and_a_reg[0]), .A2(
        cell_1735_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1735_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1735_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1735_a_HPC2_and_n9), 
        .ZN(cell_1735_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1735_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1735_a_HPC2_and_n9), 
        .ZN(cell_1735_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1735_a_HPC2_and_U8 ( .A(Fresh[21]), .ZN(cell_1735_a_HPC2_and_n9)
         );
  AND2_X1 cell_1735_a_HPC2_and_U7 ( .A1(cell_1735_and_in[1]), .A2(n427), .ZN(
        cell_1735_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1735_a_HPC2_and_U6 ( .A1(cell_1735_and_in[0]), .A2(n410), .ZN(
        cell_1735_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1735_a_HPC2_and_U5 ( .A(cell_1735_a_HPC2_and_n8), .B(
        cell_1735_a_HPC2_and_z_1__1_), .ZN(cell_1735_and_out[1]) );
  XNOR2_X1 cell_1735_a_HPC2_and_U4 ( .A(
        cell_1735_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1735_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1735_a_HPC2_and_n8) );
  XNOR2_X1 cell_1735_a_HPC2_and_U3 ( .A(cell_1735_a_HPC2_and_n7), .B(
        cell_1735_a_HPC2_and_z_0__0_), .ZN(cell_1735_and_out[0]) );
  XNOR2_X1 cell_1735_a_HPC2_and_U2 ( .A(
        cell_1735_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1735_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1735_a_HPC2_and_n7) );
  DFF_X1 cell_1735_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1735_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1735_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1735_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1735_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1735_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1735_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1735_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1735_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1735_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1736_U4 ( .A(n389), .B(cell_1736_and_out[1]), .Z(signal_3418)
         );
  XOR2_X1 cell_1736_U3 ( .A(n388), .B(cell_1736_and_out[0]), .Z(signal_2004)
         );
  XOR2_X1 cell_1736_U2 ( .A(n389), .B(1'b0), .Z(cell_1736_and_in[1]) );
  XOR2_X1 cell_1736_U1 ( .A(n388), .B(1'b1), .Z(cell_1736_and_in[0]) );
  XOR2_X1 cell_1736_a_HPC2_and_U14 ( .A(Fresh[22]), .B(cell_1736_and_in[0]), 
        .Z(cell_1736_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1736_a_HPC2_and_U13 ( .A(Fresh[22]), .B(cell_1736_and_in[1]), 
        .Z(cell_1736_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1736_a_HPC2_and_U12 ( .A1(cell_1736_a_HPC2_and_a_reg[1]), .A2(
        cell_1736_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1736_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1736_a_HPC2_and_U11 ( .A1(cell_1736_a_HPC2_and_a_reg[0]), .A2(
        cell_1736_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1736_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1736_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1736_a_HPC2_and_n9), 
        .ZN(cell_1736_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1736_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1736_a_HPC2_and_n9), 
        .ZN(cell_1736_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1736_a_HPC2_and_U8 ( .A(Fresh[22]), .ZN(cell_1736_a_HPC2_and_n9)
         );
  AND2_X1 cell_1736_a_HPC2_and_U7 ( .A1(cell_1736_and_in[1]), .A2(n427), .ZN(
        cell_1736_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1736_a_HPC2_and_U6 ( .A1(cell_1736_and_in[0]), .A2(n410), .ZN(
        cell_1736_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1736_a_HPC2_and_U5 ( .A(cell_1736_a_HPC2_and_n8), .B(
        cell_1736_a_HPC2_and_z_1__1_), .ZN(cell_1736_and_out[1]) );
  XNOR2_X1 cell_1736_a_HPC2_and_U4 ( .A(
        cell_1736_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1736_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1736_a_HPC2_and_n8) );
  XNOR2_X1 cell_1736_a_HPC2_and_U3 ( .A(cell_1736_a_HPC2_and_n7), .B(
        cell_1736_a_HPC2_and_z_0__0_), .ZN(cell_1736_and_out[0]) );
  XNOR2_X1 cell_1736_a_HPC2_and_U2 ( .A(
        cell_1736_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1736_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1736_a_HPC2_and_n7) );
  DFF_X1 cell_1736_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1736_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1736_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1736_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1736_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1736_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1736_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1736_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1736_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1736_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1737_U4 ( .A(1'b0), .B(cell_1737_and_out[1]), .Z(signal_3419)
         );
  XOR2_X1 cell_1737_U3 ( .A(1'b0), .B(cell_1737_and_out[0]), .Z(signal_2005)
         );
  XOR2_X1 cell_1737_U2 ( .A(1'b0), .B(n381), .Z(cell_1737_and_in[1]) );
  XOR2_X1 cell_1737_U1 ( .A(1'b0), .B(n380), .Z(cell_1737_and_in[0]) );
  XOR2_X1 cell_1737_a_HPC2_and_U14 ( .A(Fresh[23]), .B(cell_1737_and_in[0]), 
        .Z(cell_1737_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1737_a_HPC2_and_U13 ( .A(Fresh[23]), .B(cell_1737_and_in[1]), 
        .Z(cell_1737_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1737_a_HPC2_and_U12 ( .A1(cell_1737_a_HPC2_and_a_reg[1]), .A2(
        cell_1737_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1737_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1737_a_HPC2_and_U11 ( .A1(cell_1737_a_HPC2_and_a_reg[0]), .A2(
        cell_1737_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1737_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1737_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1737_a_HPC2_and_n9), 
        .ZN(cell_1737_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1737_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1737_a_HPC2_and_n9), 
        .ZN(cell_1737_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1737_a_HPC2_and_U8 ( .A(Fresh[23]), .ZN(cell_1737_a_HPC2_and_n9)
         );
  AND2_X1 cell_1737_a_HPC2_and_U7 ( .A1(cell_1737_and_in[1]), .A2(n427), .ZN(
        cell_1737_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1737_a_HPC2_and_U6 ( .A1(cell_1737_and_in[0]), .A2(n410), .ZN(
        cell_1737_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1737_a_HPC2_and_U5 ( .A(cell_1737_a_HPC2_and_n8), .B(
        cell_1737_a_HPC2_and_z_1__1_), .ZN(cell_1737_and_out[1]) );
  XNOR2_X1 cell_1737_a_HPC2_and_U4 ( .A(
        cell_1737_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1737_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1737_a_HPC2_and_n8) );
  XNOR2_X1 cell_1737_a_HPC2_and_U3 ( .A(cell_1737_a_HPC2_and_n7), .B(
        cell_1737_a_HPC2_and_z_0__0_), .ZN(cell_1737_and_out[0]) );
  XNOR2_X1 cell_1737_a_HPC2_and_U2 ( .A(
        cell_1737_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1737_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1737_a_HPC2_and_n7) );
  DFF_X1 cell_1737_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1737_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1737_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1737_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1737_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1737_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1737_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1737_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1737_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1737_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1738_U4 ( .A(1'b0), .B(cell_1738_and_out[1]), .Z(signal_3420)
         );
  XOR2_X1 cell_1738_U3 ( .A(1'b1), .B(cell_1738_and_out[0]), .Z(signal_2006)
         );
  XOR2_X1 cell_1738_U2 ( .A(1'b0), .B(n381), .Z(cell_1738_and_in[1]) );
  XOR2_X1 cell_1738_U1 ( .A(1'b1), .B(n380), .Z(cell_1738_and_in[0]) );
  XOR2_X1 cell_1738_a_HPC2_and_U14 ( .A(Fresh[24]), .B(cell_1738_and_in[0]), 
        .Z(cell_1738_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1738_a_HPC2_and_U13 ( .A(Fresh[24]), .B(cell_1738_and_in[1]), 
        .Z(cell_1738_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1738_a_HPC2_and_U12 ( .A1(cell_1738_a_HPC2_and_a_reg[1]), .A2(
        cell_1738_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1738_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1738_a_HPC2_and_U11 ( .A1(cell_1738_a_HPC2_and_a_reg[0]), .A2(
        cell_1738_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1738_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1738_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1738_a_HPC2_and_n9), 
        .ZN(cell_1738_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1738_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1738_a_HPC2_and_n9), 
        .ZN(cell_1738_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1738_a_HPC2_and_U8 ( .A(Fresh[24]), .ZN(cell_1738_a_HPC2_and_n9)
         );
  AND2_X1 cell_1738_a_HPC2_and_U7 ( .A1(cell_1738_and_in[1]), .A2(n427), .ZN(
        cell_1738_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1738_a_HPC2_and_U6 ( .A1(cell_1738_and_in[0]), .A2(n410), .ZN(
        cell_1738_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1738_a_HPC2_and_U5 ( .A(cell_1738_a_HPC2_and_n8), .B(
        cell_1738_a_HPC2_and_z_1__1_), .ZN(cell_1738_and_out[1]) );
  XNOR2_X1 cell_1738_a_HPC2_and_U4 ( .A(
        cell_1738_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1738_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1738_a_HPC2_and_n8) );
  XNOR2_X1 cell_1738_a_HPC2_and_U3 ( .A(cell_1738_a_HPC2_and_n7), .B(
        cell_1738_a_HPC2_and_z_0__0_), .ZN(cell_1738_and_out[0]) );
  XNOR2_X1 cell_1738_a_HPC2_and_U2 ( .A(
        cell_1738_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1738_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1738_a_HPC2_and_n7) );
  DFF_X1 cell_1738_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1738_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1738_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1738_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1738_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1738_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1738_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1738_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1738_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1738_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1739_U4 ( .A(n386), .B(cell_1739_and_out[1]), .Z(signal_3421)
         );
  XOR2_X1 cell_1739_U3 ( .A(n384), .B(cell_1739_and_out[0]), .Z(signal_2007)
         );
  XOR2_X1 cell_1739_U2 ( .A(n386), .B(1'b0), .Z(cell_1739_and_in[1]) );
  XOR2_X1 cell_1739_U1 ( .A(n384), .B(1'b0), .Z(cell_1739_and_in[0]) );
  XOR2_X1 cell_1739_a_HPC2_and_U14 ( .A(Fresh[25]), .B(cell_1739_and_in[0]), 
        .Z(cell_1739_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1739_a_HPC2_and_U13 ( .A(Fresh[25]), .B(cell_1739_and_in[1]), 
        .Z(cell_1739_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1739_a_HPC2_and_U12 ( .A1(cell_1739_a_HPC2_and_a_reg[1]), .A2(
        cell_1739_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1739_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1739_a_HPC2_and_U11 ( .A1(cell_1739_a_HPC2_and_a_reg[0]), .A2(
        cell_1739_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1739_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1739_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1739_a_HPC2_and_n9), 
        .ZN(cell_1739_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1739_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1739_a_HPC2_and_n9), 
        .ZN(cell_1739_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1739_a_HPC2_and_U8 ( .A(Fresh[25]), .ZN(cell_1739_a_HPC2_and_n9)
         );
  AND2_X1 cell_1739_a_HPC2_and_U7 ( .A1(cell_1739_and_in[1]), .A2(n427), .ZN(
        cell_1739_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1739_a_HPC2_and_U6 ( .A1(cell_1739_and_in[0]), .A2(n410), .ZN(
        cell_1739_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1739_a_HPC2_and_U5 ( .A(cell_1739_a_HPC2_and_n8), .B(
        cell_1739_a_HPC2_and_z_1__1_), .ZN(cell_1739_and_out[1]) );
  XNOR2_X1 cell_1739_a_HPC2_and_U4 ( .A(
        cell_1739_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1739_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1739_a_HPC2_and_n8) );
  XNOR2_X1 cell_1739_a_HPC2_and_U3 ( .A(cell_1739_a_HPC2_and_n7), .B(
        cell_1739_a_HPC2_and_z_0__0_), .ZN(cell_1739_and_out[0]) );
  XNOR2_X1 cell_1739_a_HPC2_and_U2 ( .A(
        cell_1739_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1739_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1739_a_HPC2_and_n7) );
  DFF_X1 cell_1739_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1739_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1739_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1739_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1739_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1739_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1739_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1739_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1739_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1739_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1740_U4 ( .A(n383), .B(cell_1740_and_out[1]), .Z(signal_3422)
         );
  XOR2_X1 cell_1740_U3 ( .A(n382), .B(cell_1740_and_out[0]), .Z(signal_2008)
         );
  XOR2_X1 cell_1740_U2 ( .A(n383), .B(1'b0), .Z(cell_1740_and_in[1]) );
  XOR2_X1 cell_1740_U1 ( .A(n382), .B(1'b0), .Z(cell_1740_and_in[0]) );
  XOR2_X1 cell_1740_a_HPC2_and_U14 ( .A(Fresh[26]), .B(cell_1740_and_in[0]), 
        .Z(cell_1740_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1740_a_HPC2_and_U13 ( .A(Fresh[26]), .B(cell_1740_and_in[1]), 
        .Z(cell_1740_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1740_a_HPC2_and_U12 ( .A1(cell_1740_a_HPC2_and_a_reg[1]), .A2(
        cell_1740_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1740_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1740_a_HPC2_and_U11 ( .A1(cell_1740_a_HPC2_and_a_reg[0]), .A2(
        cell_1740_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1740_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1740_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1740_a_HPC2_and_n9), 
        .ZN(cell_1740_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1740_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1740_a_HPC2_and_n9), 
        .ZN(cell_1740_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1740_a_HPC2_and_U8 ( .A(Fresh[26]), .ZN(cell_1740_a_HPC2_and_n9)
         );
  AND2_X1 cell_1740_a_HPC2_and_U7 ( .A1(cell_1740_and_in[1]), .A2(n427), .ZN(
        cell_1740_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1740_a_HPC2_and_U6 ( .A1(cell_1740_and_in[0]), .A2(n410), .ZN(
        cell_1740_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1740_a_HPC2_and_U5 ( .A(cell_1740_a_HPC2_and_n8), .B(
        cell_1740_a_HPC2_and_z_1__1_), .ZN(cell_1740_and_out[1]) );
  XNOR2_X1 cell_1740_a_HPC2_and_U4 ( .A(
        cell_1740_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1740_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1740_a_HPC2_and_n8) );
  XNOR2_X1 cell_1740_a_HPC2_and_U3 ( .A(cell_1740_a_HPC2_and_n7), .B(
        cell_1740_a_HPC2_and_z_0__0_), .ZN(cell_1740_and_out[0]) );
  XNOR2_X1 cell_1740_a_HPC2_and_U2 ( .A(
        cell_1740_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1740_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1740_a_HPC2_and_n7) );
  DFF_X1 cell_1740_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1740_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1740_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1740_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1740_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1740_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1740_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1740_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1740_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1740_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1741_U4 ( .A(n387), .B(cell_1741_and_out[1]), .Z(signal_3423)
         );
  XOR2_X1 cell_1741_U3 ( .A(n385), .B(cell_1741_and_out[0]), .Z(signal_2009)
         );
  XOR2_X1 cell_1741_U2 ( .A(n387), .B(n383), .Z(cell_1741_and_in[1]) );
  XOR2_X1 cell_1741_U1 ( .A(n385), .B(n382), .Z(cell_1741_and_in[0]) );
  XOR2_X1 cell_1741_a_HPC2_and_U14 ( .A(Fresh[27]), .B(cell_1741_and_in[0]), 
        .Z(cell_1741_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1741_a_HPC2_and_U13 ( .A(Fresh[27]), .B(cell_1741_and_in[1]), 
        .Z(cell_1741_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1741_a_HPC2_and_U12 ( .A1(cell_1741_a_HPC2_and_a_reg[1]), .A2(
        cell_1741_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1741_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1741_a_HPC2_and_U11 ( .A1(cell_1741_a_HPC2_and_a_reg[0]), .A2(
        cell_1741_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1741_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1741_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1741_a_HPC2_and_n9), 
        .ZN(cell_1741_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1741_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1741_a_HPC2_and_n9), 
        .ZN(cell_1741_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1741_a_HPC2_and_U8 ( .A(Fresh[27]), .ZN(cell_1741_a_HPC2_and_n9)
         );
  AND2_X1 cell_1741_a_HPC2_and_U7 ( .A1(cell_1741_and_in[1]), .A2(n411), .ZN(
        cell_1741_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1741_a_HPC2_and_U6 ( .A1(cell_1741_and_in[0]), .A2(n394), .ZN(
        cell_1741_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1741_a_HPC2_and_U5 ( .A(cell_1741_a_HPC2_and_n8), .B(
        cell_1741_a_HPC2_and_z_1__1_), .ZN(cell_1741_and_out[1]) );
  XNOR2_X1 cell_1741_a_HPC2_and_U4 ( .A(
        cell_1741_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1741_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1741_a_HPC2_and_n8) );
  XNOR2_X1 cell_1741_a_HPC2_and_U3 ( .A(cell_1741_a_HPC2_and_n7), .B(
        cell_1741_a_HPC2_and_z_0__0_), .ZN(cell_1741_and_out[0]) );
  XNOR2_X1 cell_1741_a_HPC2_and_U2 ( .A(
        cell_1741_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1741_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1741_a_HPC2_and_n7) );
  DFF_X1 cell_1741_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1741_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1741_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1741_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1741_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1741_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1741_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1741_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1741_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1741_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1742_U4 ( .A(n381), .B(1'b0), .Z(cell_1742_and_in[1]) );
  XOR2_X1 cell_1742_U3 ( .A(n380), .B(1'b1), .Z(cell_1742_and_in[0]) );
  XOR2_X1 cell_1742_U2 ( .A(n381), .B(cell_1742_and_out[1]), .Z(signal_3424)
         );
  XOR2_X1 cell_1742_U1 ( .A(n380), .B(cell_1742_and_out[0]), .Z(signal_2010)
         );
  XOR2_X1 cell_1742_a_HPC2_and_U14 ( .A(Fresh[28]), .B(cell_1742_and_in[0]), 
        .Z(cell_1742_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1742_a_HPC2_and_U13 ( .A(Fresh[28]), .B(cell_1742_and_in[1]), 
        .Z(cell_1742_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1742_a_HPC2_and_U12 ( .A1(cell_1742_a_HPC2_and_a_reg[1]), .A2(
        cell_1742_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1742_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1742_a_HPC2_and_U11 ( .A1(cell_1742_a_HPC2_and_a_reg[0]), .A2(
        cell_1742_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1742_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1742_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1742_a_HPC2_and_n9), 
        .ZN(cell_1742_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1742_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1742_a_HPC2_and_n9), 
        .ZN(cell_1742_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1742_a_HPC2_and_U8 ( .A(Fresh[28]), .ZN(cell_1742_a_HPC2_and_n9)
         );
  AND2_X1 cell_1742_a_HPC2_and_U7 ( .A1(cell_1742_and_in[1]), .A2(n393), .ZN(
        cell_1742_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1742_a_HPC2_and_U6 ( .A1(cell_1742_and_in[0]), .A2(n392), .ZN(
        cell_1742_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1742_a_HPC2_and_U5 ( .A(cell_1742_a_HPC2_and_n8), .B(
        cell_1742_a_HPC2_and_z_1__1_), .ZN(cell_1742_and_out[1]) );
  XNOR2_X1 cell_1742_a_HPC2_and_U4 ( .A(
        cell_1742_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1742_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1742_a_HPC2_and_n8) );
  XNOR2_X1 cell_1742_a_HPC2_and_U3 ( .A(cell_1742_a_HPC2_and_n7), .B(
        cell_1742_a_HPC2_and_z_0__0_), .ZN(cell_1742_and_out[0]) );
  XNOR2_X1 cell_1742_a_HPC2_and_U2 ( .A(
        cell_1742_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1742_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1742_a_HPC2_and_n7) );
  DFF_X1 cell_1742_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1742_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1742_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1742_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1742_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1742_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1742_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1742_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1742_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1742_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1743_U4 ( .A(n389), .B(cell_1743_and_out[1]), .Z(signal_3425)
         );
  XOR2_X1 cell_1743_U3 ( .A(n388), .B(cell_1743_and_out[0]), .Z(signal_2011)
         );
  XOR2_X1 cell_1743_U2 ( .A(n389), .B(signal_3261), .Z(cell_1743_and_in[1]) );
  XOR2_X1 cell_1743_U1 ( .A(n388), .B(signal_1987), .Z(cell_1743_and_in[0]) );
  XOR2_X1 cell_1743_a_HPC2_and_U14 ( .A(Fresh[29]), .B(cell_1743_and_in[0]), 
        .Z(cell_1743_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1743_a_HPC2_and_U13 ( .A(Fresh[29]), .B(cell_1743_and_in[1]), 
        .Z(cell_1743_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1743_a_HPC2_and_U12 ( .A1(cell_1743_a_HPC2_and_a_reg[1]), .A2(
        cell_1743_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1743_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1743_a_HPC2_and_U11 ( .A1(cell_1743_a_HPC2_and_a_reg[0]), .A2(
        cell_1743_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1743_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1743_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1743_a_HPC2_and_n9), 
        .ZN(cell_1743_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1743_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1743_a_HPC2_and_n9), 
        .ZN(cell_1743_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1743_a_HPC2_and_U8 ( .A(Fresh[29]), .ZN(cell_1743_a_HPC2_and_n9)
         );
  AND2_X1 cell_1743_a_HPC2_and_U7 ( .A1(cell_1743_and_in[1]), .A2(n412), .ZN(
        cell_1743_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1743_a_HPC2_and_U6 ( .A1(cell_1743_and_in[0]), .A2(n395), .ZN(
        cell_1743_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1743_a_HPC2_and_U5 ( .A(cell_1743_a_HPC2_and_n8), .B(
        cell_1743_a_HPC2_and_z_1__1_), .ZN(cell_1743_and_out[1]) );
  XNOR2_X1 cell_1743_a_HPC2_and_U4 ( .A(
        cell_1743_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1743_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1743_a_HPC2_and_n8) );
  XNOR2_X1 cell_1743_a_HPC2_and_U3 ( .A(cell_1743_a_HPC2_and_n7), .B(
        cell_1743_a_HPC2_and_z_0__0_), .ZN(cell_1743_and_out[0]) );
  XNOR2_X1 cell_1743_a_HPC2_and_U2 ( .A(
        cell_1743_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1743_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1743_a_HPC2_and_n7) );
  DFF_X1 cell_1743_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1743_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1743_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1743_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1743_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1743_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1743_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1743_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1743_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1743_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1744_U4 ( .A(n389), .B(1'b0), .Z(cell_1744_and_in[1]) );
  XOR2_X1 cell_1744_U3 ( .A(n388), .B(1'b0), .Z(cell_1744_and_in[0]) );
  XOR2_X2 cell_1744_U2 ( .A(n389), .B(cell_1744_and_out[1]), .Z(signal_3426)
         );
  XOR2_X2 cell_1744_U1 ( .A(n388), .B(cell_1744_and_out[0]), .Z(signal_2012)
         );
  XOR2_X1 cell_1744_a_HPC2_and_U14 ( .A(Fresh[30]), .B(cell_1744_and_in[0]), 
        .Z(cell_1744_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1744_a_HPC2_and_U13 ( .A(Fresh[30]), .B(cell_1744_and_in[1]), 
        .Z(cell_1744_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1744_a_HPC2_and_U12 ( .A1(cell_1744_a_HPC2_and_a_reg[1]), .A2(
        cell_1744_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1744_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1744_a_HPC2_and_U11 ( .A1(cell_1744_a_HPC2_and_a_reg[0]), .A2(
        cell_1744_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1744_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1744_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1744_a_HPC2_and_n9), 
        .ZN(cell_1744_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1744_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1744_a_HPC2_and_n9), 
        .ZN(cell_1744_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1744_a_HPC2_and_U8 ( .A(Fresh[30]), .ZN(cell_1744_a_HPC2_and_n9)
         );
  AND2_X1 cell_1744_a_HPC2_and_U7 ( .A1(cell_1744_and_in[1]), .A2(n393), .ZN(
        cell_1744_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1744_a_HPC2_and_U6 ( .A1(cell_1744_and_in[0]), .A2(n392), .ZN(
        cell_1744_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1744_a_HPC2_and_U5 ( .A(cell_1744_a_HPC2_and_n8), .B(
        cell_1744_a_HPC2_and_z_1__1_), .ZN(cell_1744_and_out[1]) );
  XNOR2_X1 cell_1744_a_HPC2_and_U4 ( .A(
        cell_1744_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1744_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1744_a_HPC2_and_n8) );
  XNOR2_X1 cell_1744_a_HPC2_and_U3 ( .A(cell_1744_a_HPC2_and_n7), .B(
        cell_1744_a_HPC2_and_z_0__0_), .ZN(cell_1744_and_out[0]) );
  XNOR2_X1 cell_1744_a_HPC2_and_U2 ( .A(
        cell_1744_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1744_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1744_a_HPC2_and_n7) );
  DFF_X1 cell_1744_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1744_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1744_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1744_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1744_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1744_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1744_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1744_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1744_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1744_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1745_U4 ( .A(n389), .B(n381), .Z(cell_1745_and_in[1]) );
  XOR2_X1 cell_1745_U3 ( .A(n388), .B(n380), .Z(cell_1745_and_in[0]) );
  XOR2_X1 cell_1745_U2 ( .A(n388), .B(cell_1745_and_out[0]), .Z(signal_2013)
         );
  XOR2_X1 cell_1745_U1 ( .A(n389), .B(cell_1745_and_out[1]), .Z(signal_3427)
         );
  XOR2_X1 cell_1745_a_HPC2_and_U14 ( .A(Fresh[31]), .B(cell_1745_and_in[0]), 
        .Z(cell_1745_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1745_a_HPC2_and_U13 ( .A(Fresh[31]), .B(cell_1745_and_in[1]), 
        .Z(cell_1745_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1745_a_HPC2_and_U12 ( .A1(cell_1745_a_HPC2_and_a_reg[1]), .A2(
        cell_1745_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1745_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1745_a_HPC2_and_U11 ( .A1(cell_1745_a_HPC2_and_a_reg[0]), .A2(
        cell_1745_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1745_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1745_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1745_a_HPC2_and_n9), 
        .ZN(cell_1745_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1745_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1745_a_HPC2_and_n9), 
        .ZN(cell_1745_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1745_a_HPC2_and_U8 ( .A(Fresh[31]), .ZN(cell_1745_a_HPC2_and_n9)
         );
  AND2_X1 cell_1745_a_HPC2_and_U7 ( .A1(cell_1745_and_in[1]), .A2(n393), .ZN(
        cell_1745_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1745_a_HPC2_and_U6 ( .A1(cell_1745_and_in[0]), .A2(n392), .ZN(
        cell_1745_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1745_a_HPC2_and_U5 ( .A(cell_1745_a_HPC2_and_n8), .B(
        cell_1745_a_HPC2_and_z_1__1_), .ZN(cell_1745_and_out[1]) );
  XNOR2_X1 cell_1745_a_HPC2_and_U4 ( .A(
        cell_1745_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1745_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1745_a_HPC2_and_n8) );
  XNOR2_X1 cell_1745_a_HPC2_and_U3 ( .A(cell_1745_a_HPC2_and_n7), .B(
        cell_1745_a_HPC2_and_z_0__0_), .ZN(cell_1745_and_out[0]) );
  XNOR2_X1 cell_1745_a_HPC2_and_U2 ( .A(
        cell_1745_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1745_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1745_a_HPC2_and_n7) );
  DFF_X1 cell_1745_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1745_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1745_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1745_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1745_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1745_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1745_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1745_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1745_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1745_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1746_U4 ( .A(n383), .B(cell_1746_and_out[1]), .Z(signal_3428)
         );
  XOR2_X1 cell_1746_U3 ( .A(n382), .B(cell_1746_and_out[0]), .Z(signal_2014)
         );
  XOR2_X1 cell_1746_U2 ( .A(n383), .B(n381), .Z(cell_1746_and_in[1]) );
  XOR2_X1 cell_1746_U1 ( .A(n382), .B(n380), .Z(cell_1746_and_in[0]) );
  XOR2_X1 cell_1746_a_HPC2_and_U14 ( .A(Fresh[32]), .B(cell_1746_and_in[0]), 
        .Z(cell_1746_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1746_a_HPC2_and_U13 ( .A(Fresh[32]), .B(cell_1746_and_in[1]), 
        .Z(cell_1746_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1746_a_HPC2_and_U12 ( .A1(cell_1746_a_HPC2_and_a_reg[1]), .A2(
        cell_1746_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1746_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1746_a_HPC2_and_U11 ( .A1(cell_1746_a_HPC2_and_a_reg[0]), .A2(
        cell_1746_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1746_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1746_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1746_a_HPC2_and_n9), 
        .ZN(cell_1746_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1746_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1746_a_HPC2_and_n9), 
        .ZN(cell_1746_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1746_a_HPC2_and_U8 ( .A(Fresh[32]), .ZN(cell_1746_a_HPC2_and_n9)
         );
  AND2_X1 cell_1746_a_HPC2_and_U7 ( .A1(cell_1746_and_in[1]), .A2(n412), .ZN(
        cell_1746_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1746_a_HPC2_and_U6 ( .A1(cell_1746_and_in[0]), .A2(n395), .ZN(
        cell_1746_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1746_a_HPC2_and_U5 ( .A(cell_1746_a_HPC2_and_n8), .B(
        cell_1746_a_HPC2_and_z_1__1_), .ZN(cell_1746_and_out[1]) );
  XNOR2_X1 cell_1746_a_HPC2_and_U4 ( .A(
        cell_1746_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1746_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1746_a_HPC2_and_n8) );
  XNOR2_X1 cell_1746_a_HPC2_and_U3 ( .A(cell_1746_a_HPC2_and_n7), .B(
        cell_1746_a_HPC2_and_z_0__0_), .ZN(cell_1746_and_out[0]) );
  XNOR2_X1 cell_1746_a_HPC2_and_U2 ( .A(
        cell_1746_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1746_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1746_a_HPC2_and_n7) );
  DFF_X1 cell_1746_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1746_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1746_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1746_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1746_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1746_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1746_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1746_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1746_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1746_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1747_U4 ( .A(n381), .B(1'b0), .Z(cell_1747_and_in[1]) );
  XOR2_X1 cell_1747_U3 ( .A(n380), .B(1'b0), .Z(cell_1747_and_in[0]) );
  XOR2_X1 cell_1747_U2 ( .A(n381), .B(cell_1747_and_out[1]), .Z(signal_3429)
         );
  XOR2_X1 cell_1747_U1 ( .A(n380), .B(cell_1747_and_out[0]), .Z(signal_2015)
         );
  XOR2_X1 cell_1747_a_HPC2_and_U14 ( .A(Fresh[33]), .B(cell_1747_and_in[0]), 
        .Z(cell_1747_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1747_a_HPC2_and_U13 ( .A(Fresh[33]), .B(cell_1747_and_in[1]), 
        .Z(cell_1747_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1747_a_HPC2_and_U12 ( .A1(cell_1747_a_HPC2_and_a_reg[1]), .A2(
        cell_1747_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1747_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1747_a_HPC2_and_U11 ( .A1(cell_1747_a_HPC2_and_a_reg[0]), .A2(
        cell_1747_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1747_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1747_a_HPC2_and_U10 ( .A1(n393), .A2(cell_1747_a_HPC2_and_n9), 
        .ZN(cell_1747_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1747_a_HPC2_and_U9 ( .A1(n392), .A2(cell_1747_a_HPC2_and_n9), 
        .ZN(cell_1747_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1747_a_HPC2_and_U8 ( .A(Fresh[33]), .ZN(cell_1747_a_HPC2_and_n9)
         );
  AND2_X1 cell_1747_a_HPC2_and_U7 ( .A1(cell_1747_and_in[1]), .A2(n393), .ZN(
        cell_1747_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1747_a_HPC2_and_U6 ( .A1(cell_1747_and_in[0]), .A2(n392), .ZN(
        cell_1747_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1747_a_HPC2_and_U5 ( .A(cell_1747_a_HPC2_and_n8), .B(
        cell_1747_a_HPC2_and_z_1__1_), .ZN(cell_1747_and_out[1]) );
  XNOR2_X1 cell_1747_a_HPC2_and_U4 ( .A(
        cell_1747_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1747_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1747_a_HPC2_and_n8) );
  XNOR2_X1 cell_1747_a_HPC2_and_U3 ( .A(cell_1747_a_HPC2_and_n7), .B(
        cell_1747_a_HPC2_and_z_0__0_), .ZN(cell_1747_and_out[0]) );
  XNOR2_X1 cell_1747_a_HPC2_and_U2 ( .A(
        cell_1747_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1747_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1747_a_HPC2_and_n7) );
  DFF_X1 cell_1747_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1747_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1747_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n392), .CK(clk), 
        .Q(cell_1747_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1747_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1747_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n393), .CK(clk), 
        .Q(cell_1747_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1747_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1747_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1747_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1748_U4 ( .A(n381), .B(cell_1748_and_out[1]), .Z(signal_3430)
         );
  XOR2_X1 cell_1748_U3 ( .A(n380), .B(cell_1748_and_out[0]), .Z(signal_2016)
         );
  XOR2_X1 cell_1748_U2 ( .A(n381), .B(signal_3256), .Z(cell_1748_and_in[1]) );
  XOR2_X1 cell_1748_U1 ( .A(n380), .B(signal_1982), .Z(cell_1748_and_in[0]) );
  XOR2_X1 cell_1748_a_HPC2_and_U14 ( .A(Fresh[34]), .B(cell_1748_and_in[0]), 
        .Z(cell_1748_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1748_a_HPC2_and_U13 ( .A(Fresh[34]), .B(cell_1748_and_in[1]), 
        .Z(cell_1748_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1748_a_HPC2_and_U12 ( .A1(cell_1748_a_HPC2_and_a_reg[1]), .A2(
        cell_1748_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1748_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1748_a_HPC2_and_U11 ( .A1(cell_1748_a_HPC2_and_a_reg[0]), .A2(
        cell_1748_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1748_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1748_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1748_a_HPC2_and_n9), 
        .ZN(cell_1748_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1748_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1748_a_HPC2_and_n9), 
        .ZN(cell_1748_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1748_a_HPC2_and_U8 ( .A(Fresh[34]), .ZN(cell_1748_a_HPC2_and_n9)
         );
  AND2_X1 cell_1748_a_HPC2_and_U7 ( .A1(cell_1748_and_in[1]), .A2(n412), .ZN(
        cell_1748_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1748_a_HPC2_and_U6 ( .A1(cell_1748_and_in[0]), .A2(n395), .ZN(
        cell_1748_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1748_a_HPC2_and_U5 ( .A(cell_1748_a_HPC2_and_n8), .B(
        cell_1748_a_HPC2_and_z_1__1_), .ZN(cell_1748_and_out[1]) );
  XNOR2_X1 cell_1748_a_HPC2_and_U4 ( .A(
        cell_1748_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1748_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1748_a_HPC2_and_n8) );
  XNOR2_X1 cell_1748_a_HPC2_and_U3 ( .A(cell_1748_a_HPC2_and_n7), .B(
        cell_1748_a_HPC2_and_z_0__0_), .ZN(cell_1748_and_out[0]) );
  XNOR2_X1 cell_1748_a_HPC2_and_U2 ( .A(
        cell_1748_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1748_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1748_a_HPC2_and_n7) );
  DFF_X1 cell_1748_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1748_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1748_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1748_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1748_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1748_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1748_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1748_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1748_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1748_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1749_U4 ( .A(n387), .B(cell_1749_and_out[1]), .Z(signal_3431)
         );
  XOR2_X1 cell_1749_U3 ( .A(n385), .B(cell_1749_and_out[0]), .Z(signal_2017)
         );
  XOR2_X1 cell_1749_U2 ( .A(n387), .B(n381), .Z(cell_1749_and_in[1]) );
  XOR2_X1 cell_1749_U1 ( .A(n385), .B(n380), .Z(cell_1749_and_in[0]) );
  XOR2_X1 cell_1749_a_HPC2_and_U14 ( .A(Fresh[35]), .B(cell_1749_and_in[0]), 
        .Z(cell_1749_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1749_a_HPC2_and_U13 ( .A(Fresh[35]), .B(cell_1749_and_in[1]), 
        .Z(cell_1749_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1749_a_HPC2_and_U12 ( .A1(cell_1749_a_HPC2_and_a_reg[1]), .A2(
        cell_1749_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1749_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1749_a_HPC2_and_U11 ( .A1(cell_1749_a_HPC2_and_a_reg[0]), .A2(
        cell_1749_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1749_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1749_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1749_a_HPC2_and_n9), 
        .ZN(cell_1749_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1749_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1749_a_HPC2_and_n9), 
        .ZN(cell_1749_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1749_a_HPC2_and_U8 ( .A(Fresh[35]), .ZN(cell_1749_a_HPC2_and_n9)
         );
  AND2_X1 cell_1749_a_HPC2_and_U7 ( .A1(cell_1749_and_in[1]), .A2(n412), .ZN(
        cell_1749_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1749_a_HPC2_and_U6 ( .A1(cell_1749_and_in[0]), .A2(n395), .ZN(
        cell_1749_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1749_a_HPC2_and_U5 ( .A(cell_1749_a_HPC2_and_n8), .B(
        cell_1749_a_HPC2_and_z_1__1_), .ZN(cell_1749_and_out[1]) );
  XNOR2_X1 cell_1749_a_HPC2_and_U4 ( .A(
        cell_1749_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1749_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1749_a_HPC2_and_n8) );
  XNOR2_X1 cell_1749_a_HPC2_and_U3 ( .A(cell_1749_a_HPC2_and_n7), .B(
        cell_1749_a_HPC2_and_z_0__0_), .ZN(cell_1749_and_out[0]) );
  XNOR2_X1 cell_1749_a_HPC2_and_U2 ( .A(
        cell_1749_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1749_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1749_a_HPC2_and_n7) );
  DFF_X1 cell_1749_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1749_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1749_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1749_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1749_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1749_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1749_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1749_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1749_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1749_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1750_U4 ( .A(n386), .B(cell_1750_and_out[1]), .Z(signal_3432)
         );
  XOR2_X1 cell_1750_U3 ( .A(n384), .B(cell_1750_and_out[0]), .Z(signal_2018)
         );
  XOR2_X1 cell_1750_U2 ( .A(n386), .B(1'b0), .Z(cell_1750_and_in[1]) );
  XOR2_X1 cell_1750_U1 ( .A(n384), .B(1'b1), .Z(cell_1750_and_in[0]) );
  XOR2_X1 cell_1750_a_HPC2_and_U14 ( .A(Fresh[36]), .B(cell_1750_and_in[0]), 
        .Z(cell_1750_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1750_a_HPC2_and_U13 ( .A(Fresh[36]), .B(cell_1750_and_in[1]), 
        .Z(cell_1750_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1750_a_HPC2_and_U12 ( .A1(cell_1750_a_HPC2_and_a_reg[1]), .A2(
        cell_1750_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1750_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1750_a_HPC2_and_U11 ( .A1(cell_1750_a_HPC2_and_a_reg[0]), .A2(
        cell_1750_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1750_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1750_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1750_a_HPC2_and_n9), 
        .ZN(cell_1750_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1750_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1750_a_HPC2_and_n9), 
        .ZN(cell_1750_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1750_a_HPC2_and_U8 ( .A(Fresh[36]), .ZN(cell_1750_a_HPC2_and_n9)
         );
  AND2_X1 cell_1750_a_HPC2_and_U7 ( .A1(cell_1750_and_in[1]), .A2(n421), .ZN(
        cell_1750_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1750_a_HPC2_and_U6 ( .A1(cell_1750_and_in[0]), .A2(n404), .ZN(
        cell_1750_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1750_a_HPC2_and_U5 ( .A(cell_1750_a_HPC2_and_n8), .B(
        cell_1750_a_HPC2_and_z_1__1_), .ZN(cell_1750_and_out[1]) );
  XNOR2_X1 cell_1750_a_HPC2_and_U4 ( .A(
        cell_1750_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1750_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1750_a_HPC2_and_n8) );
  XNOR2_X1 cell_1750_a_HPC2_and_U3 ( .A(cell_1750_a_HPC2_and_n7), .B(
        cell_1750_a_HPC2_and_z_0__0_), .ZN(cell_1750_and_out[0]) );
  XNOR2_X1 cell_1750_a_HPC2_and_U2 ( .A(
        cell_1750_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1750_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1750_a_HPC2_and_n7) );
  DFF_X1 cell_1750_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1750_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1750_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1750_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1750_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1750_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1750_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1750_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1750_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1750_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1751_U4 ( .A(n383), .B(cell_1751_and_out[1]), .Z(signal_3433)
         );
  XOR2_X1 cell_1751_U3 ( .A(n382), .B(cell_1751_and_out[0]), .Z(signal_2019)
         );
  XOR2_X1 cell_1751_U2 ( .A(n383), .B(1'b0), .Z(cell_1751_and_in[1]) );
  XOR2_X1 cell_1751_U1 ( .A(n382), .B(1'b1), .Z(cell_1751_and_in[0]) );
  XOR2_X1 cell_1751_a_HPC2_and_U14 ( .A(Fresh[37]), .B(cell_1751_and_in[0]), 
        .Z(cell_1751_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1751_a_HPC2_and_U13 ( .A(Fresh[37]), .B(cell_1751_and_in[1]), 
        .Z(cell_1751_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1751_a_HPC2_and_U12 ( .A1(cell_1751_a_HPC2_and_a_reg[1]), .A2(
        cell_1751_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1751_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1751_a_HPC2_and_U11 ( .A1(cell_1751_a_HPC2_and_a_reg[0]), .A2(
        cell_1751_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1751_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1751_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1751_a_HPC2_and_n9), 
        .ZN(cell_1751_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1751_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1751_a_HPC2_and_n9), 
        .ZN(cell_1751_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1751_a_HPC2_and_U8 ( .A(Fresh[37]), .ZN(cell_1751_a_HPC2_and_n9)
         );
  AND2_X1 cell_1751_a_HPC2_and_U7 ( .A1(cell_1751_and_in[1]), .A2(n417), .ZN(
        cell_1751_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1751_a_HPC2_and_U6 ( .A1(cell_1751_and_in[0]), .A2(n400), .ZN(
        cell_1751_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1751_a_HPC2_and_U5 ( .A(cell_1751_a_HPC2_and_n8), .B(
        cell_1751_a_HPC2_and_z_1__1_), .ZN(cell_1751_and_out[1]) );
  XNOR2_X1 cell_1751_a_HPC2_and_U4 ( .A(
        cell_1751_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1751_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1751_a_HPC2_and_n8) );
  XNOR2_X1 cell_1751_a_HPC2_and_U3 ( .A(cell_1751_a_HPC2_and_n7), .B(
        cell_1751_a_HPC2_and_z_0__0_), .ZN(cell_1751_and_out[0]) );
  XNOR2_X1 cell_1751_a_HPC2_and_U2 ( .A(
        cell_1751_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1751_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1751_a_HPC2_and_n7) );
  DFF_X1 cell_1751_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1751_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1751_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1751_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1751_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1751_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1751_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1751_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1751_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1751_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1752_U4 ( .A(n389), .B(cell_1752_and_out[1]), .Z(signal_3458)
         );
  XOR2_X1 cell_1752_U3 ( .A(n388), .B(cell_1752_and_out[0]), .Z(signal_2020)
         );
  XOR2_X1 cell_1752_U2 ( .A(n389), .B(n379), .Z(cell_1752_and_in[1]) );
  XOR2_X1 cell_1752_U1 ( .A(n388), .B(n377), .Z(cell_1752_and_in[0]) );
  XOR2_X1 cell_1752_a_HPC2_and_U14 ( .A(Fresh[38]), .B(cell_1752_and_in[0]), 
        .Z(cell_1752_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1752_a_HPC2_and_U13 ( .A(Fresh[38]), .B(cell_1752_and_in[1]), 
        .Z(cell_1752_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1752_a_HPC2_and_U12 ( .A1(cell_1752_a_HPC2_and_a_reg[1]), .A2(
        cell_1752_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1752_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1752_a_HPC2_and_U11 ( .A1(cell_1752_a_HPC2_and_a_reg[0]), .A2(
        cell_1752_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1752_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1752_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1752_a_HPC2_and_n9), 
        .ZN(cell_1752_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1752_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1752_a_HPC2_and_n9), 
        .ZN(cell_1752_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1752_a_HPC2_and_U8 ( .A(Fresh[38]), .ZN(cell_1752_a_HPC2_and_n9)
         );
  AND2_X1 cell_1752_a_HPC2_and_U7 ( .A1(cell_1752_and_in[1]), .A2(n412), .ZN(
        cell_1752_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1752_a_HPC2_and_U6 ( .A1(cell_1752_and_in[0]), .A2(n395), .ZN(
        cell_1752_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1752_a_HPC2_and_U5 ( .A(cell_1752_a_HPC2_and_n8), .B(
        cell_1752_a_HPC2_and_z_1__1_), .ZN(cell_1752_and_out[1]) );
  XNOR2_X1 cell_1752_a_HPC2_and_U4 ( .A(
        cell_1752_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1752_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1752_a_HPC2_and_n8) );
  XNOR2_X1 cell_1752_a_HPC2_and_U3 ( .A(cell_1752_a_HPC2_and_n7), .B(
        cell_1752_a_HPC2_and_z_0__0_), .ZN(cell_1752_and_out[0]) );
  XNOR2_X1 cell_1752_a_HPC2_and_U2 ( .A(
        cell_1752_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1752_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1752_a_HPC2_and_n7) );
  DFF_X1 cell_1752_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1752_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1752_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1752_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1752_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1752_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1752_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1752_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1752_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1752_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1753_U4 ( .A(1'b0), .B(cell_1753_and_out[1]), .Z(signal_3459)
         );
  XOR2_X1 cell_1753_U3 ( .A(1'b1), .B(cell_1753_and_out[0]), .Z(signal_2021)
         );
  XOR2_X1 cell_1753_U2 ( .A(1'b0), .B(signal_3426), .Z(cell_1753_and_in[1]) );
  XOR2_X1 cell_1753_U1 ( .A(1'b1), .B(signal_2012), .Z(cell_1753_and_in[0]) );
  XOR2_X1 cell_1753_a_HPC2_and_U14 ( .A(Fresh[39]), .B(cell_1753_and_in[0]), 
        .Z(cell_1753_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1753_a_HPC2_and_U13 ( .A(Fresh[39]), .B(cell_1753_and_in[1]), 
        .Z(cell_1753_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1753_a_HPC2_and_U12 ( .A1(cell_1753_a_HPC2_and_a_reg[1]), .A2(
        cell_1753_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1753_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1753_a_HPC2_and_U11 ( .A1(cell_1753_a_HPC2_and_a_reg[0]), .A2(
        cell_1753_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1753_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1753_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1753_a_HPC2_and_n9), 
        .ZN(cell_1753_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1753_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1753_a_HPC2_and_n9), 
        .ZN(cell_1753_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1753_a_HPC2_and_U8 ( .A(Fresh[39]), .ZN(cell_1753_a_HPC2_and_n9)
         );
  AND2_X1 cell_1753_a_HPC2_and_U7 ( .A1(cell_1753_and_in[1]), .A2(n416), .ZN(
        cell_1753_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1753_a_HPC2_and_U6 ( .A1(cell_1753_and_in[0]), .A2(n399), .ZN(
        cell_1753_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1753_a_HPC2_and_U5 ( .A(cell_1753_a_HPC2_and_n8), .B(
        cell_1753_a_HPC2_and_z_1__1_), .ZN(cell_1753_and_out[1]) );
  XNOR2_X1 cell_1753_a_HPC2_and_U4 ( .A(
        cell_1753_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1753_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1753_a_HPC2_and_n8) );
  XNOR2_X1 cell_1753_a_HPC2_and_U3 ( .A(cell_1753_a_HPC2_and_n7), .B(
        cell_1753_a_HPC2_and_z_0__0_), .ZN(cell_1753_and_out[0]) );
  XNOR2_X1 cell_1753_a_HPC2_and_U2 ( .A(
        cell_1753_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1753_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1753_a_HPC2_and_n7) );
  DFF_X1 cell_1753_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1753_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1753_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1753_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1753_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1753_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1753_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1753_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1753_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1753_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1754_U4 ( .A(n374), .B(cell_1754_and_out[1]), .Z(signal_3460)
         );
  XOR2_X1 cell_1754_U3 ( .A(n372), .B(cell_1754_and_out[0]), .Z(signal_2022)
         );
  XOR2_X1 cell_1754_U2 ( .A(n374), .B(n383), .Z(cell_1754_and_in[1]) );
  XOR2_X1 cell_1754_U1 ( .A(n372), .B(n382), .Z(cell_1754_and_in[0]) );
  XOR2_X1 cell_1754_a_HPC2_and_U14 ( .A(Fresh[40]), .B(cell_1754_and_in[0]), 
        .Z(cell_1754_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1754_a_HPC2_and_U13 ( .A(Fresh[40]), .B(cell_1754_and_in[1]), 
        .Z(cell_1754_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1754_a_HPC2_and_U12 ( .A1(cell_1754_a_HPC2_and_a_reg[1]), .A2(
        cell_1754_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1754_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1754_a_HPC2_and_U11 ( .A1(cell_1754_a_HPC2_and_a_reg[0]), .A2(
        cell_1754_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1754_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1754_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1754_a_HPC2_and_n9), 
        .ZN(cell_1754_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1754_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1754_a_HPC2_and_n9), 
        .ZN(cell_1754_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1754_a_HPC2_and_U8 ( .A(Fresh[40]), .ZN(cell_1754_a_HPC2_and_n9)
         );
  AND2_X1 cell_1754_a_HPC2_and_U7 ( .A1(cell_1754_and_in[1]), .A2(n412), .ZN(
        cell_1754_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1754_a_HPC2_and_U6 ( .A1(cell_1754_and_in[0]), .A2(n395), .ZN(
        cell_1754_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1754_a_HPC2_and_U5 ( .A(cell_1754_a_HPC2_and_n8), .B(
        cell_1754_a_HPC2_and_z_1__1_), .ZN(cell_1754_and_out[1]) );
  XNOR2_X1 cell_1754_a_HPC2_and_U4 ( .A(
        cell_1754_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1754_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1754_a_HPC2_and_n8) );
  XNOR2_X1 cell_1754_a_HPC2_and_U3 ( .A(cell_1754_a_HPC2_and_n7), .B(
        cell_1754_a_HPC2_and_z_0__0_), .ZN(cell_1754_and_out[0]) );
  XNOR2_X1 cell_1754_a_HPC2_and_U2 ( .A(
        cell_1754_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1754_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1754_a_HPC2_and_n7) );
  DFF_X1 cell_1754_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1754_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1754_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1754_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1754_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1754_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1754_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1754_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1754_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1754_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1755_U4 ( .A(1'b0), .B(cell_1755_and_out[1]), .Z(signal_3461)
         );
  XOR2_X1 cell_1755_U3 ( .A(1'b0), .B(cell_1755_and_out[0]), .Z(signal_2023)
         );
  XOR2_X1 cell_1755_U2 ( .A(1'b0), .B(n365), .Z(cell_1755_and_in[1]) );
  XOR2_X1 cell_1755_U1 ( .A(1'b0), .B(n363), .Z(cell_1755_and_in[0]) );
  XOR2_X1 cell_1755_a_HPC2_and_U14 ( .A(Fresh[41]), .B(cell_1755_and_in[0]), 
        .Z(cell_1755_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1755_a_HPC2_and_U13 ( .A(Fresh[41]), .B(cell_1755_and_in[1]), 
        .Z(cell_1755_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1755_a_HPC2_and_U12 ( .A1(cell_1755_a_HPC2_and_a_reg[1]), .A2(
        cell_1755_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1755_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1755_a_HPC2_and_U11 ( .A1(cell_1755_a_HPC2_and_a_reg[0]), .A2(
        cell_1755_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1755_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1755_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1755_a_HPC2_and_n9), 
        .ZN(cell_1755_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1755_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1755_a_HPC2_and_n9), 
        .ZN(cell_1755_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1755_a_HPC2_and_U8 ( .A(Fresh[41]), .ZN(cell_1755_a_HPC2_and_n9)
         );
  AND2_X1 cell_1755_a_HPC2_and_U7 ( .A1(cell_1755_and_in[1]), .A2(n411), .ZN(
        cell_1755_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1755_a_HPC2_and_U6 ( .A1(cell_1755_and_in[0]), .A2(n394), .ZN(
        cell_1755_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1755_a_HPC2_and_U5 ( .A(cell_1755_a_HPC2_and_n8), .B(
        cell_1755_a_HPC2_and_z_1__1_), .ZN(cell_1755_and_out[1]) );
  XNOR2_X1 cell_1755_a_HPC2_and_U4 ( .A(
        cell_1755_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1755_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1755_a_HPC2_and_n8) );
  XNOR2_X1 cell_1755_a_HPC2_and_U3 ( .A(cell_1755_a_HPC2_and_n7), .B(
        cell_1755_a_HPC2_and_z_0__0_), .ZN(cell_1755_and_out[0]) );
  XNOR2_X1 cell_1755_a_HPC2_and_U2 ( .A(
        cell_1755_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1755_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1755_a_HPC2_and_n7) );
  DFF_X1 cell_1755_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1755_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1755_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1755_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1755_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1755_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1755_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1755_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1755_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1755_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1756_U4 ( .A(n383), .B(cell_1756_and_out[1]), .Z(signal_3462)
         );
  XOR2_X1 cell_1756_U3 ( .A(n382), .B(cell_1756_and_out[0]), .Z(signal_2024)
         );
  XOR2_X1 cell_1756_U2 ( .A(n383), .B(n371), .Z(cell_1756_and_in[1]) );
  XOR2_X1 cell_1756_U1 ( .A(n382), .B(n369), .Z(cell_1756_and_in[0]) );
  XOR2_X1 cell_1756_a_HPC2_and_U14 ( .A(Fresh[42]), .B(cell_1756_and_in[0]), 
        .Z(cell_1756_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1756_a_HPC2_and_U13 ( .A(Fresh[42]), .B(cell_1756_and_in[1]), 
        .Z(cell_1756_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1756_a_HPC2_and_U12 ( .A1(cell_1756_a_HPC2_and_a_reg[1]), .A2(
        cell_1756_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1756_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1756_a_HPC2_and_U11 ( .A1(cell_1756_a_HPC2_and_a_reg[0]), .A2(
        cell_1756_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1756_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1756_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1756_a_HPC2_and_n9), 
        .ZN(cell_1756_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1756_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1756_a_HPC2_and_n9), 
        .ZN(cell_1756_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1756_a_HPC2_and_U8 ( .A(Fresh[42]), .ZN(cell_1756_a_HPC2_and_n9)
         );
  AND2_X1 cell_1756_a_HPC2_and_U7 ( .A1(cell_1756_and_in[1]), .A2(n412), .ZN(
        cell_1756_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1756_a_HPC2_and_U6 ( .A1(cell_1756_and_in[0]), .A2(n395), .ZN(
        cell_1756_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1756_a_HPC2_and_U5 ( .A(cell_1756_a_HPC2_and_n8), .B(
        cell_1756_a_HPC2_and_z_1__1_), .ZN(cell_1756_and_out[1]) );
  XNOR2_X1 cell_1756_a_HPC2_and_U4 ( .A(
        cell_1756_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1756_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1756_a_HPC2_and_n8) );
  XNOR2_X1 cell_1756_a_HPC2_and_U3 ( .A(cell_1756_a_HPC2_and_n7), .B(
        cell_1756_a_HPC2_and_z_0__0_), .ZN(cell_1756_and_out[0]) );
  XNOR2_X1 cell_1756_a_HPC2_and_U2 ( .A(
        cell_1756_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1756_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1756_a_HPC2_and_n7) );
  DFF_X1 cell_1756_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1756_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1756_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1756_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1756_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1756_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1756_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1756_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1756_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1756_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1757_U4 ( .A(n365), .B(cell_1757_and_out[1]), .Z(signal_3463)
         );
  XOR2_X1 cell_1757_U3 ( .A(n363), .B(cell_1757_and_out[0]), .Z(signal_2025)
         );
  XOR2_X1 cell_1757_U2 ( .A(n365), .B(n381), .Z(cell_1757_and_in[1]) );
  XOR2_X1 cell_1757_U1 ( .A(n363), .B(n380), .Z(cell_1757_and_in[0]) );
  XOR2_X1 cell_1757_a_HPC2_and_U14 ( .A(Fresh[43]), .B(cell_1757_and_in[0]), 
        .Z(cell_1757_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1757_a_HPC2_and_U13 ( .A(Fresh[43]), .B(cell_1757_and_in[1]), 
        .Z(cell_1757_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1757_a_HPC2_and_U12 ( .A1(cell_1757_a_HPC2_and_a_reg[1]), .A2(
        cell_1757_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1757_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1757_a_HPC2_and_U11 ( .A1(cell_1757_a_HPC2_and_a_reg[0]), .A2(
        cell_1757_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1757_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1757_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1757_a_HPC2_and_n9), 
        .ZN(cell_1757_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1757_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1757_a_HPC2_and_n9), 
        .ZN(cell_1757_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1757_a_HPC2_and_U8 ( .A(Fresh[43]), .ZN(cell_1757_a_HPC2_and_n9)
         );
  AND2_X1 cell_1757_a_HPC2_and_U7 ( .A1(cell_1757_and_in[1]), .A2(n413), .ZN(
        cell_1757_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1757_a_HPC2_and_U6 ( .A1(cell_1757_and_in[0]), .A2(n396), .ZN(
        cell_1757_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1757_a_HPC2_and_U5 ( .A(cell_1757_a_HPC2_and_n8), .B(
        cell_1757_a_HPC2_and_z_1__1_), .ZN(cell_1757_and_out[1]) );
  XNOR2_X1 cell_1757_a_HPC2_and_U4 ( .A(
        cell_1757_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1757_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1757_a_HPC2_and_n8) );
  XNOR2_X1 cell_1757_a_HPC2_and_U3 ( .A(cell_1757_a_HPC2_and_n7), .B(
        cell_1757_a_HPC2_and_z_0__0_), .ZN(cell_1757_and_out[0]) );
  XNOR2_X1 cell_1757_a_HPC2_and_U2 ( .A(
        cell_1757_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1757_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1757_a_HPC2_and_n7) );
  DFF_X1 cell_1757_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1757_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1757_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1757_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1757_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1757_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1757_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1757_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1757_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1757_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1758_U4 ( .A(1'b0), .B(cell_1758_and_out[1]), .Z(signal_3464)
         );
  XOR2_X1 cell_1758_U3 ( .A(1'b0), .B(cell_1758_and_out[0]), .Z(signal_2026)
         );
  XOR2_X1 cell_1758_U2 ( .A(1'b0), .B(n375), .Z(cell_1758_and_in[1]) );
  XOR2_X1 cell_1758_U1 ( .A(1'b0), .B(n373), .Z(cell_1758_and_in[0]) );
  XOR2_X1 cell_1758_a_HPC2_and_U14 ( .A(Fresh[44]), .B(cell_1758_and_in[0]), 
        .Z(cell_1758_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1758_a_HPC2_and_U13 ( .A(Fresh[44]), .B(cell_1758_and_in[1]), 
        .Z(cell_1758_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1758_a_HPC2_and_U12 ( .A1(cell_1758_a_HPC2_and_a_reg[1]), .A2(
        cell_1758_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1758_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1758_a_HPC2_and_U11 ( .A1(cell_1758_a_HPC2_and_a_reg[0]), .A2(
        cell_1758_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1758_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1758_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1758_a_HPC2_and_n9), 
        .ZN(cell_1758_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1758_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1758_a_HPC2_and_n9), 
        .ZN(cell_1758_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1758_a_HPC2_and_U8 ( .A(Fresh[44]), .ZN(cell_1758_a_HPC2_and_n9)
         );
  AND2_X1 cell_1758_a_HPC2_and_U7 ( .A1(cell_1758_and_in[1]), .A2(n426), .ZN(
        cell_1758_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1758_a_HPC2_and_U6 ( .A1(cell_1758_and_in[0]), .A2(n409), .ZN(
        cell_1758_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1758_a_HPC2_and_U5 ( .A(cell_1758_a_HPC2_and_n8), .B(
        cell_1758_a_HPC2_and_z_1__1_), .ZN(cell_1758_and_out[1]) );
  XNOR2_X1 cell_1758_a_HPC2_and_U4 ( .A(
        cell_1758_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1758_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1758_a_HPC2_and_n8) );
  XNOR2_X1 cell_1758_a_HPC2_and_U3 ( .A(cell_1758_a_HPC2_and_n7), .B(
        cell_1758_a_HPC2_and_z_0__0_), .ZN(cell_1758_and_out[0]) );
  XNOR2_X1 cell_1758_a_HPC2_and_U2 ( .A(
        cell_1758_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1758_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1758_a_HPC2_and_n7) );
  DFF_X1 cell_1758_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1758_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1758_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1758_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1758_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1758_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1758_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1758_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1758_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1758_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1759_U4 ( .A(n357), .B(cell_1759_and_out[1]), .Z(signal_3465)
         );
  XOR2_X1 cell_1759_U3 ( .A(n356), .B(cell_1759_and_out[0]), .Z(signal_2027)
         );
  XOR2_X1 cell_1759_U2 ( .A(n357), .B(signal_3406), .Z(cell_1759_and_in[1]) );
  XOR2_X1 cell_1759_U1 ( .A(n356), .B(signal_1992), .Z(cell_1759_and_in[0]) );
  XOR2_X1 cell_1759_a_HPC2_and_U14 ( .A(Fresh[45]), .B(cell_1759_and_in[0]), 
        .Z(cell_1759_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1759_a_HPC2_and_U13 ( .A(Fresh[45]), .B(cell_1759_and_in[1]), 
        .Z(cell_1759_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1759_a_HPC2_and_U12 ( .A1(cell_1759_a_HPC2_and_a_reg[1]), .A2(
        cell_1759_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1759_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1759_a_HPC2_and_U11 ( .A1(cell_1759_a_HPC2_and_a_reg[0]), .A2(
        cell_1759_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1759_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1759_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1759_a_HPC2_and_n9), 
        .ZN(cell_1759_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1759_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1759_a_HPC2_and_n9), 
        .ZN(cell_1759_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1759_a_HPC2_and_U8 ( .A(Fresh[45]), .ZN(cell_1759_a_HPC2_and_n9)
         );
  AND2_X1 cell_1759_a_HPC2_and_U7 ( .A1(cell_1759_and_in[1]), .A2(n413), .ZN(
        cell_1759_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1759_a_HPC2_and_U6 ( .A1(cell_1759_and_in[0]), .A2(n396), .ZN(
        cell_1759_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1759_a_HPC2_and_U5 ( .A(cell_1759_a_HPC2_and_n8), .B(
        cell_1759_a_HPC2_and_z_1__1_), .ZN(cell_1759_and_out[1]) );
  XNOR2_X1 cell_1759_a_HPC2_and_U4 ( .A(
        cell_1759_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1759_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1759_a_HPC2_and_n8) );
  XNOR2_X1 cell_1759_a_HPC2_and_U3 ( .A(cell_1759_a_HPC2_and_n7), .B(
        cell_1759_a_HPC2_and_z_0__0_), .ZN(cell_1759_and_out[0]) );
  XNOR2_X1 cell_1759_a_HPC2_and_U2 ( .A(
        cell_1759_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1759_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1759_a_HPC2_and_n7) );
  DFF_X1 cell_1759_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1759_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1759_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1759_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1759_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1759_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1759_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1759_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1759_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1759_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1760_U6 ( .A(cell_1760_n4), .B(cell_1760_and_out[1]), .Z(
        signal_3466) );
  XOR2_X1 cell_1760_U5 ( .A(cell_1760_n3), .B(cell_1760_and_out[0]), .Z(
        signal_2028) );
  XOR2_X1 cell_1760_U4 ( .A(cell_1760_n4), .B(n375), .Z(cell_1760_and_in[1])
         );
  XOR2_X1 cell_1760_U3 ( .A(cell_1760_n3), .B(n373), .Z(cell_1760_and_in[0])
         );
  BUF_X1 cell_1760_U2 ( .A(signal_3426), .Z(cell_1760_n4) );
  BUF_X1 cell_1760_U1 ( .A(signal_2012), .Z(cell_1760_n3) );
  XOR2_X1 cell_1760_a_HPC2_and_U14 ( .A(Fresh[46]), .B(cell_1760_and_in[0]), 
        .Z(cell_1760_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1760_a_HPC2_and_U13 ( .A(Fresh[46]), .B(cell_1760_and_in[1]), 
        .Z(cell_1760_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1760_a_HPC2_and_U12 ( .A1(cell_1760_a_HPC2_and_a_reg[1]), .A2(
        cell_1760_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1760_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1760_a_HPC2_and_U11 ( .A1(cell_1760_a_HPC2_and_a_reg[0]), .A2(
        cell_1760_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1760_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1760_a_HPC2_and_U10 ( .A1(signal_3237), .A2(
        cell_1760_a_HPC2_and_n9), .ZN(cell_1760_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1760_a_HPC2_and_U9 ( .A1(signal_1512), .A2(
        cell_1760_a_HPC2_and_n9), .ZN(cell_1760_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1760_a_HPC2_and_U8 ( .A(Fresh[46]), .ZN(cell_1760_a_HPC2_and_n9)
         );
  AND2_X1 cell_1760_a_HPC2_and_U7 ( .A1(cell_1760_and_in[1]), .A2(signal_3237), 
        .ZN(cell_1760_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1760_a_HPC2_and_U6 ( .A1(cell_1760_and_in[0]), .A2(signal_1512), 
        .ZN(cell_1760_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1760_a_HPC2_and_U5 ( .A(cell_1760_a_HPC2_and_n8), .B(
        cell_1760_a_HPC2_and_z_1__1_), .ZN(cell_1760_and_out[1]) );
  XNOR2_X1 cell_1760_a_HPC2_and_U4 ( .A(
        cell_1760_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1760_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1760_a_HPC2_and_n8) );
  XNOR2_X1 cell_1760_a_HPC2_and_U3 ( .A(cell_1760_a_HPC2_and_n7), .B(
        cell_1760_a_HPC2_and_z_0__0_), .ZN(cell_1760_and_out[0]) );
  XNOR2_X1 cell_1760_a_HPC2_and_U2 ( .A(
        cell_1760_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1760_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1760_a_HPC2_and_n7) );
  DFF_X1 cell_1760_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1760_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1760_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1512), 
        .CK(clk), .Q(cell_1760_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1760_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1760_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3237), 
        .CK(clk), .Q(cell_1760_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1760_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1760_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1760_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1761_U4 ( .A(n374), .B(cell_1761_and_out[1]), .Z(signal_3467)
         );
  XOR2_X1 cell_1761_U3 ( .A(n372), .B(cell_1761_and_out[0]), .Z(signal_2029)
         );
  XOR2_X1 cell_1761_U2 ( .A(n374), .B(signal_3426), .Z(cell_1761_and_in[1]) );
  XOR2_X1 cell_1761_U1 ( .A(n372), .B(signal_2012), .Z(cell_1761_and_in[0]) );
  XOR2_X1 cell_1761_a_HPC2_and_U14 ( .A(Fresh[47]), .B(cell_1761_and_in[0]), 
        .Z(cell_1761_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1761_a_HPC2_and_U13 ( .A(Fresh[47]), .B(cell_1761_and_in[1]), 
        .Z(cell_1761_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1761_a_HPC2_and_U12 ( .A1(cell_1761_a_HPC2_and_a_reg[1]), .A2(
        cell_1761_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1761_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1761_a_HPC2_and_U11 ( .A1(cell_1761_a_HPC2_and_a_reg[0]), .A2(
        cell_1761_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1761_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1761_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1761_a_HPC2_and_n9), 
        .ZN(cell_1761_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1761_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1761_a_HPC2_and_n9), 
        .ZN(cell_1761_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1761_a_HPC2_and_U8 ( .A(Fresh[47]), .ZN(cell_1761_a_HPC2_and_n9)
         );
  AND2_X1 cell_1761_a_HPC2_and_U7 ( .A1(cell_1761_and_in[1]), .A2(n413), .ZN(
        cell_1761_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1761_a_HPC2_and_U6 ( .A1(cell_1761_and_in[0]), .A2(n396), .ZN(
        cell_1761_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1761_a_HPC2_and_U5 ( .A(cell_1761_a_HPC2_and_n8), .B(
        cell_1761_a_HPC2_and_z_1__1_), .ZN(cell_1761_and_out[1]) );
  XNOR2_X1 cell_1761_a_HPC2_and_U4 ( .A(
        cell_1761_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1761_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1761_a_HPC2_and_n8) );
  XNOR2_X1 cell_1761_a_HPC2_and_U3 ( .A(cell_1761_a_HPC2_and_n7), .B(
        cell_1761_a_HPC2_and_z_0__0_), .ZN(cell_1761_and_out[0]) );
  XNOR2_X1 cell_1761_a_HPC2_and_U2 ( .A(
        cell_1761_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1761_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1761_a_HPC2_and_n7) );
  DFF_X1 cell_1761_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1761_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1761_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1761_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1761_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1761_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1761_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1761_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1761_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1761_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1762_U4 ( .A(n354), .B(cell_1762_and_out[1]), .Z(signal_3468)
         );
  XOR2_X1 cell_1762_U3 ( .A(n352), .B(cell_1762_and_out[0]), .Z(signal_2030)
         );
  XOR2_X1 cell_1762_U2 ( .A(n354), .B(n360), .Z(cell_1762_and_in[1]) );
  XOR2_X1 cell_1762_U1 ( .A(n352), .B(n358), .Z(cell_1762_and_in[0]) );
  XOR2_X1 cell_1762_a_HPC2_and_U14 ( .A(Fresh[48]), .B(cell_1762_and_in[0]), 
        .Z(cell_1762_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1762_a_HPC2_and_U13 ( .A(Fresh[48]), .B(cell_1762_and_in[1]), 
        .Z(cell_1762_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1762_a_HPC2_and_U12 ( .A1(cell_1762_a_HPC2_and_a_reg[1]), .A2(
        cell_1762_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1762_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1762_a_HPC2_and_U11 ( .A1(cell_1762_a_HPC2_and_a_reg[0]), .A2(
        cell_1762_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1762_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1762_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1762_a_HPC2_and_n9), 
        .ZN(cell_1762_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1762_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1762_a_HPC2_and_n9), 
        .ZN(cell_1762_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1762_a_HPC2_and_U8 ( .A(Fresh[48]), .ZN(cell_1762_a_HPC2_and_n9)
         );
  AND2_X1 cell_1762_a_HPC2_and_U7 ( .A1(cell_1762_and_in[1]), .A2(n413), .ZN(
        cell_1762_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1762_a_HPC2_and_U6 ( .A1(cell_1762_and_in[0]), .A2(n396), .ZN(
        cell_1762_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1762_a_HPC2_and_U5 ( .A(cell_1762_a_HPC2_and_n8), .B(
        cell_1762_a_HPC2_and_z_1__1_), .ZN(cell_1762_and_out[1]) );
  XNOR2_X1 cell_1762_a_HPC2_and_U4 ( .A(
        cell_1762_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1762_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1762_a_HPC2_and_n8) );
  XNOR2_X1 cell_1762_a_HPC2_and_U3 ( .A(cell_1762_a_HPC2_and_n7), .B(
        cell_1762_a_HPC2_and_z_0__0_), .ZN(cell_1762_and_out[0]) );
  XNOR2_X1 cell_1762_a_HPC2_and_U2 ( .A(
        cell_1762_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1762_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1762_a_HPC2_and_n7) );
  DFF_X1 cell_1762_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1762_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1762_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1762_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1762_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1762_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1762_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1762_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1762_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1762_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1763_U4 ( .A(n389), .B(cell_1763_and_out[1]), .Z(signal_3469)
         );
  XOR2_X1 cell_1763_U3 ( .A(n388), .B(cell_1763_and_out[0]), .Z(signal_2031)
         );
  XOR2_X1 cell_1763_U2 ( .A(n389), .B(n367), .Z(cell_1763_and_in[1]) );
  XOR2_X1 cell_1763_U1 ( .A(n388), .B(n366), .Z(cell_1763_and_in[0]) );
  XOR2_X1 cell_1763_a_HPC2_and_U14 ( .A(Fresh[49]), .B(cell_1763_and_in[0]), 
        .Z(cell_1763_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1763_a_HPC2_and_U13 ( .A(Fresh[49]), .B(cell_1763_and_in[1]), 
        .Z(cell_1763_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1763_a_HPC2_and_U12 ( .A1(cell_1763_a_HPC2_and_a_reg[1]), .A2(
        cell_1763_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1763_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1763_a_HPC2_and_U11 ( .A1(cell_1763_a_HPC2_and_a_reg[0]), .A2(
        cell_1763_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1763_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1763_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1763_a_HPC2_and_n9), 
        .ZN(cell_1763_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1763_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1763_a_HPC2_and_n9), 
        .ZN(cell_1763_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1763_a_HPC2_and_U8 ( .A(Fresh[49]), .ZN(cell_1763_a_HPC2_and_n9)
         );
  AND2_X1 cell_1763_a_HPC2_and_U7 ( .A1(cell_1763_and_in[1]), .A2(n413), .ZN(
        cell_1763_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1763_a_HPC2_and_U6 ( .A1(cell_1763_and_in[0]), .A2(n396), .ZN(
        cell_1763_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1763_a_HPC2_and_U5 ( .A(cell_1763_a_HPC2_and_n8), .B(
        cell_1763_a_HPC2_and_z_1__1_), .ZN(cell_1763_and_out[1]) );
  XNOR2_X1 cell_1763_a_HPC2_and_U4 ( .A(
        cell_1763_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1763_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1763_a_HPC2_and_n8) );
  XNOR2_X1 cell_1763_a_HPC2_and_U3 ( .A(cell_1763_a_HPC2_and_n7), .B(
        cell_1763_a_HPC2_and_z_0__0_), .ZN(cell_1763_and_out[0]) );
  XNOR2_X1 cell_1763_a_HPC2_and_U2 ( .A(
        cell_1763_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1763_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1763_a_HPC2_and_n7) );
  DFF_X1 cell_1763_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1763_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1763_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1763_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1763_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1763_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1763_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1763_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1763_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1763_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1764_U4 ( .A(n387), .B(cell_1764_and_out[1]), .Z(signal_3470)
         );
  XOR2_X1 cell_1764_U3 ( .A(n385), .B(cell_1764_and_out[0]), .Z(signal_2032)
         );
  XOR2_X1 cell_1764_U2 ( .A(n387), .B(n355), .Z(cell_1764_and_in[1]) );
  XOR2_X1 cell_1764_U1 ( .A(n385), .B(n353), .Z(cell_1764_and_in[0]) );
  XOR2_X1 cell_1764_a_HPC2_and_U14 ( .A(Fresh[50]), .B(cell_1764_and_in[0]), 
        .Z(cell_1764_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1764_a_HPC2_and_U13 ( .A(Fresh[50]), .B(cell_1764_and_in[1]), 
        .Z(cell_1764_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1764_a_HPC2_and_U12 ( .A1(cell_1764_a_HPC2_and_a_reg[1]), .A2(
        cell_1764_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1764_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1764_a_HPC2_and_U11 ( .A1(cell_1764_a_HPC2_and_a_reg[0]), .A2(
        cell_1764_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1764_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1764_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1764_a_HPC2_and_n9), 
        .ZN(cell_1764_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1764_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1764_a_HPC2_and_n9), 
        .ZN(cell_1764_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1764_a_HPC2_and_U8 ( .A(Fresh[50]), .ZN(cell_1764_a_HPC2_and_n9)
         );
  AND2_X1 cell_1764_a_HPC2_and_U7 ( .A1(cell_1764_and_in[1]), .A2(n413), .ZN(
        cell_1764_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1764_a_HPC2_and_U6 ( .A1(cell_1764_and_in[0]), .A2(n396), .ZN(
        cell_1764_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1764_a_HPC2_and_U5 ( .A(cell_1764_a_HPC2_and_n8), .B(
        cell_1764_a_HPC2_and_z_1__1_), .ZN(cell_1764_and_out[1]) );
  XNOR2_X1 cell_1764_a_HPC2_and_U4 ( .A(
        cell_1764_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1764_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1764_a_HPC2_and_n8) );
  XNOR2_X1 cell_1764_a_HPC2_and_U3 ( .A(cell_1764_a_HPC2_and_n7), .B(
        cell_1764_a_HPC2_and_z_0__0_), .ZN(cell_1764_and_out[0]) );
  XNOR2_X1 cell_1764_a_HPC2_and_U2 ( .A(
        cell_1764_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1764_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1764_a_HPC2_and_n7) );
  DFF_X1 cell_1764_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1764_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1764_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1764_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1764_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1764_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1764_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1764_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1764_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1764_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1765_U4 ( .A(n361), .B(cell_1765_and_out[1]), .Z(signal_3471)
         );
  XOR2_X1 cell_1765_U3 ( .A(n359), .B(cell_1765_and_out[0]), .Z(signal_2033)
         );
  XOR2_X1 cell_1765_U2 ( .A(n361), .B(signal_3418), .Z(cell_1765_and_in[1]) );
  XOR2_X1 cell_1765_U1 ( .A(n359), .B(signal_2004), .Z(cell_1765_and_in[0]) );
  XOR2_X1 cell_1765_a_HPC2_and_U14 ( .A(Fresh[51]), .B(cell_1765_and_in[0]), 
        .Z(cell_1765_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1765_a_HPC2_and_U13 ( .A(Fresh[51]), .B(cell_1765_and_in[1]), 
        .Z(cell_1765_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1765_a_HPC2_and_U12 ( .A1(cell_1765_a_HPC2_and_a_reg[1]), .A2(
        cell_1765_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1765_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1765_a_HPC2_and_U11 ( .A1(cell_1765_a_HPC2_and_a_reg[0]), .A2(
        cell_1765_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1765_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1765_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1765_a_HPC2_and_n9), 
        .ZN(cell_1765_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1765_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1765_a_HPC2_and_n9), 
        .ZN(cell_1765_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1765_a_HPC2_and_U8 ( .A(Fresh[51]), .ZN(cell_1765_a_HPC2_and_n9)
         );
  AND2_X1 cell_1765_a_HPC2_and_U7 ( .A1(cell_1765_and_in[1]), .A2(n442), .ZN(
        cell_1765_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1765_a_HPC2_and_U6 ( .A1(cell_1765_and_in[0]), .A2(n428), .ZN(
        cell_1765_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1765_a_HPC2_and_U5 ( .A(cell_1765_a_HPC2_and_n8), .B(
        cell_1765_a_HPC2_and_z_1__1_), .ZN(cell_1765_and_out[1]) );
  XNOR2_X1 cell_1765_a_HPC2_and_U4 ( .A(
        cell_1765_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1765_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1765_a_HPC2_and_n8) );
  XNOR2_X1 cell_1765_a_HPC2_and_U3 ( .A(cell_1765_a_HPC2_and_n7), .B(
        cell_1765_a_HPC2_and_z_0__0_), .ZN(cell_1765_and_out[0]) );
  XNOR2_X1 cell_1765_a_HPC2_and_U2 ( .A(
        cell_1765_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1765_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1765_a_HPC2_and_n7) );
  DFF_X1 cell_1765_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1765_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1765_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1765_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1765_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1765_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1765_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1765_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1765_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1765_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1766_U4 ( .A(n383), .B(cell_1766_and_out[1]), .Z(signal_3472)
         );
  XOR2_X1 cell_1766_U3 ( .A(n382), .B(cell_1766_and_out[0]), .Z(signal_2034)
         );
  XOR2_X1 cell_1766_U2 ( .A(n383), .B(n357), .Z(cell_1766_and_in[1]) );
  XOR2_X1 cell_1766_U1 ( .A(n382), .B(n356), .Z(cell_1766_and_in[0]) );
  XOR2_X1 cell_1766_a_HPC2_and_U14 ( .A(Fresh[52]), .B(cell_1766_and_in[0]), 
        .Z(cell_1766_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1766_a_HPC2_and_U13 ( .A(Fresh[52]), .B(cell_1766_and_in[1]), 
        .Z(cell_1766_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1766_a_HPC2_and_U12 ( .A1(cell_1766_a_HPC2_and_a_reg[1]), .A2(
        cell_1766_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1766_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1766_a_HPC2_and_U11 ( .A1(cell_1766_a_HPC2_and_a_reg[0]), .A2(
        cell_1766_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1766_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1766_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1766_a_HPC2_and_n9), 
        .ZN(cell_1766_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1766_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1766_a_HPC2_and_n9), 
        .ZN(cell_1766_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1766_a_HPC2_and_U8 ( .A(Fresh[52]), .ZN(cell_1766_a_HPC2_and_n9)
         );
  AND2_X1 cell_1766_a_HPC2_and_U7 ( .A1(cell_1766_and_in[1]), .A2(n413), .ZN(
        cell_1766_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1766_a_HPC2_and_U6 ( .A1(cell_1766_and_in[0]), .A2(n396), .ZN(
        cell_1766_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1766_a_HPC2_and_U5 ( .A(cell_1766_a_HPC2_and_n8), .B(
        cell_1766_a_HPC2_and_z_1__1_), .ZN(cell_1766_and_out[1]) );
  XNOR2_X1 cell_1766_a_HPC2_and_U4 ( .A(
        cell_1766_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1766_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1766_a_HPC2_and_n8) );
  XNOR2_X1 cell_1766_a_HPC2_and_U3 ( .A(cell_1766_a_HPC2_and_n7), .B(
        cell_1766_a_HPC2_and_z_0__0_), .ZN(cell_1766_and_out[0]) );
  XNOR2_X1 cell_1766_a_HPC2_and_U2 ( .A(
        cell_1766_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1766_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1766_a_HPC2_and_n7) );
  DFF_X1 cell_1766_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1766_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1766_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1766_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1766_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1766_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1766_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1766_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1766_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1766_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1767_U4 ( .A(signal_3427), .B(cell_1767_and_out[1]), .Z(
        signal_3473) );
  XOR2_X1 cell_1767_U3 ( .A(n356), .B(cell_1767_and_out[0]), .Z(signal_2035)
         );
  XOR2_X1 cell_1767_U2 ( .A(signal_3427), .B(n367), .Z(cell_1767_and_in[1]) );
  XOR2_X1 cell_1767_U1 ( .A(n356), .B(n366), .Z(cell_1767_and_in[0]) );
  XOR2_X1 cell_1767_a_HPC2_and_U14 ( .A(Fresh[53]), .B(cell_1767_and_in[0]), 
        .Z(cell_1767_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1767_a_HPC2_and_U13 ( .A(Fresh[53]), .B(cell_1767_and_in[1]), 
        .Z(cell_1767_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1767_a_HPC2_and_U12 ( .A1(cell_1767_a_HPC2_and_a_reg[1]), .A2(
        cell_1767_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1767_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1767_a_HPC2_and_U11 ( .A1(cell_1767_a_HPC2_and_a_reg[0]), .A2(
        cell_1767_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1767_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1767_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1767_a_HPC2_and_n9), 
        .ZN(cell_1767_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1767_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1767_a_HPC2_and_n9), 
        .ZN(cell_1767_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1767_a_HPC2_and_U8 ( .A(Fresh[53]), .ZN(cell_1767_a_HPC2_and_n9)
         );
  AND2_X1 cell_1767_a_HPC2_and_U7 ( .A1(cell_1767_and_in[1]), .A2(n414), .ZN(
        cell_1767_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1767_a_HPC2_and_U6 ( .A1(cell_1767_and_in[0]), .A2(n397), .ZN(
        cell_1767_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1767_a_HPC2_and_U5 ( .A(cell_1767_a_HPC2_and_n8), .B(
        cell_1767_a_HPC2_and_z_1__1_), .ZN(cell_1767_and_out[1]) );
  XNOR2_X1 cell_1767_a_HPC2_and_U4 ( .A(
        cell_1767_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1767_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1767_a_HPC2_and_n8) );
  XNOR2_X1 cell_1767_a_HPC2_and_U3 ( .A(cell_1767_a_HPC2_and_n7), .B(
        cell_1767_a_HPC2_and_z_0__0_), .ZN(cell_1767_and_out[0]) );
  XNOR2_X1 cell_1767_a_HPC2_and_U2 ( .A(
        cell_1767_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1767_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1767_a_HPC2_and_n7) );
  DFF_X1 cell_1767_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1767_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1767_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1767_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1767_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1767_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1767_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1767_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1767_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1767_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1768_U4 ( .A(n370), .B(cell_1768_and_out[1]), .Z(signal_3474)
         );
  XOR2_X1 cell_1768_U3 ( .A(n368), .B(cell_1768_and_out[0]), .Z(signal_2036)
         );
  XOR2_X1 cell_1768_U2 ( .A(n370), .B(signal_3261), .Z(cell_1768_and_in[1]) );
  XOR2_X1 cell_1768_U1 ( .A(n368), .B(signal_1987), .Z(cell_1768_and_in[0]) );
  XOR2_X1 cell_1768_a_HPC2_and_U14 ( .A(Fresh[54]), .B(cell_1768_and_in[0]), 
        .Z(cell_1768_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1768_a_HPC2_and_U13 ( .A(Fresh[54]), .B(cell_1768_and_in[1]), 
        .Z(cell_1768_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1768_a_HPC2_and_U12 ( .A1(cell_1768_a_HPC2_and_a_reg[1]), .A2(
        cell_1768_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1768_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1768_a_HPC2_and_U11 ( .A1(cell_1768_a_HPC2_and_a_reg[0]), .A2(
        cell_1768_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1768_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1768_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1768_a_HPC2_and_n9), 
        .ZN(cell_1768_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1768_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1768_a_HPC2_and_n9), 
        .ZN(cell_1768_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1768_a_HPC2_and_U8 ( .A(Fresh[54]), .ZN(cell_1768_a_HPC2_and_n9)
         );
  AND2_X1 cell_1768_a_HPC2_and_U7 ( .A1(cell_1768_and_in[1]), .A2(n414), .ZN(
        cell_1768_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1768_a_HPC2_and_U6 ( .A1(cell_1768_and_in[0]), .A2(n397), .ZN(
        cell_1768_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1768_a_HPC2_and_U5 ( .A(cell_1768_a_HPC2_and_n8), .B(
        cell_1768_a_HPC2_and_z_1__1_), .ZN(cell_1768_and_out[1]) );
  XNOR2_X1 cell_1768_a_HPC2_and_U4 ( .A(
        cell_1768_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1768_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1768_a_HPC2_and_n8) );
  XNOR2_X1 cell_1768_a_HPC2_and_U3 ( .A(cell_1768_a_HPC2_and_n7), .B(
        cell_1768_a_HPC2_and_z_0__0_), .ZN(cell_1768_and_out[0]) );
  XNOR2_X1 cell_1768_a_HPC2_and_U2 ( .A(
        cell_1768_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1768_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1768_a_HPC2_and_n7) );
  DFF_X1 cell_1768_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1768_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1768_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1768_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1768_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1768_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1768_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1768_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1768_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1768_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1769_U4 ( .A(n374), .B(cell_1769_and_out[1]), .Z(signal_3475)
         );
  XOR2_X1 cell_1769_U3 ( .A(n372), .B(cell_1769_and_out[0]), .Z(signal_2037)
         );
  XOR2_X1 cell_1769_U2 ( .A(n374), .B(n360), .Z(cell_1769_and_in[1]) );
  XOR2_X1 cell_1769_U1 ( .A(n372), .B(n358), .Z(cell_1769_and_in[0]) );
  XOR2_X1 cell_1769_a_HPC2_and_U14 ( .A(Fresh[55]), .B(cell_1769_and_in[0]), 
        .Z(cell_1769_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1769_a_HPC2_and_U13 ( .A(Fresh[55]), .B(cell_1769_and_in[1]), 
        .Z(cell_1769_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1769_a_HPC2_and_U12 ( .A1(cell_1769_a_HPC2_and_a_reg[1]), .A2(
        cell_1769_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1769_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1769_a_HPC2_and_U11 ( .A1(cell_1769_a_HPC2_and_a_reg[0]), .A2(
        cell_1769_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1769_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1769_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1769_a_HPC2_and_n9), 
        .ZN(cell_1769_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1769_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1769_a_HPC2_and_n9), 
        .ZN(cell_1769_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1769_a_HPC2_and_U8 ( .A(Fresh[55]), .ZN(cell_1769_a_HPC2_and_n9)
         );
  AND2_X1 cell_1769_a_HPC2_and_U7 ( .A1(cell_1769_and_in[1]), .A2(n414), .ZN(
        cell_1769_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1769_a_HPC2_and_U6 ( .A1(cell_1769_and_in[0]), .A2(n397), .ZN(
        cell_1769_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1769_a_HPC2_and_U5 ( .A(cell_1769_a_HPC2_and_n8), .B(
        cell_1769_a_HPC2_and_z_1__1_), .ZN(cell_1769_and_out[1]) );
  XNOR2_X1 cell_1769_a_HPC2_and_U4 ( .A(
        cell_1769_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1769_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1769_a_HPC2_and_n8) );
  XNOR2_X1 cell_1769_a_HPC2_and_U3 ( .A(cell_1769_a_HPC2_and_n7), .B(
        cell_1769_a_HPC2_and_z_0__0_), .ZN(cell_1769_and_out[0]) );
  XNOR2_X1 cell_1769_a_HPC2_and_U2 ( .A(
        cell_1769_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1769_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1769_a_HPC2_and_n7) );
  DFF_X1 cell_1769_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1769_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1769_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1769_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1769_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1769_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1769_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1769_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1769_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1769_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1770_U4 ( .A(n354), .B(cell_1770_and_out[1]), .Z(signal_3476)
         );
  XOR2_X1 cell_1770_U3 ( .A(n352), .B(cell_1770_and_out[0]), .Z(signal_2038)
         );
  XOR2_X1 cell_1770_U2 ( .A(n354), .B(n357), .Z(cell_1770_and_in[1]) );
  XOR2_X1 cell_1770_U1 ( .A(n352), .B(n356), .Z(cell_1770_and_in[0]) );
  XOR2_X1 cell_1770_a_HPC2_and_U14 ( .A(Fresh[56]), .B(cell_1770_and_in[0]), 
        .Z(cell_1770_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1770_a_HPC2_and_U13 ( .A(Fresh[56]), .B(cell_1770_and_in[1]), 
        .Z(cell_1770_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1770_a_HPC2_and_U12 ( .A1(cell_1770_a_HPC2_and_a_reg[1]), .A2(
        cell_1770_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1770_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1770_a_HPC2_and_U11 ( .A1(cell_1770_a_HPC2_and_a_reg[0]), .A2(
        cell_1770_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1770_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1770_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1770_a_HPC2_and_n9), 
        .ZN(cell_1770_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1770_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1770_a_HPC2_and_n9), 
        .ZN(cell_1770_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1770_a_HPC2_and_U8 ( .A(Fresh[56]), .ZN(cell_1770_a_HPC2_and_n9)
         );
  AND2_X1 cell_1770_a_HPC2_and_U7 ( .A1(cell_1770_and_in[1]), .A2(n414), .ZN(
        cell_1770_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1770_a_HPC2_and_U6 ( .A1(cell_1770_and_in[0]), .A2(n397), .ZN(
        cell_1770_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1770_a_HPC2_and_U5 ( .A(cell_1770_a_HPC2_and_n8), .B(
        cell_1770_a_HPC2_and_z_1__1_), .ZN(cell_1770_and_out[1]) );
  XNOR2_X1 cell_1770_a_HPC2_and_U4 ( .A(
        cell_1770_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1770_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1770_a_HPC2_and_n8) );
  XNOR2_X1 cell_1770_a_HPC2_and_U3 ( .A(cell_1770_a_HPC2_and_n7), .B(
        cell_1770_a_HPC2_and_z_0__0_), .ZN(cell_1770_and_out[0]) );
  XNOR2_X1 cell_1770_a_HPC2_and_U2 ( .A(
        cell_1770_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1770_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1770_a_HPC2_and_n7) );
  DFF_X1 cell_1770_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1770_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1770_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1770_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1770_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1770_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1770_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1770_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1770_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1770_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1771_U4 ( .A(n365), .B(cell_1771_and_out[1]), .Z(signal_3477)
         );
  XOR2_X1 cell_1771_U3 ( .A(n363), .B(cell_1771_and_out[0]), .Z(signal_2039)
         );
  XOR2_X1 cell_1771_U2 ( .A(n365), .B(signal_3407), .Z(cell_1771_and_in[1]) );
  XOR2_X1 cell_1771_U1 ( .A(n363), .B(signal_1993), .Z(cell_1771_and_in[0]) );
  XOR2_X1 cell_1771_a_HPC2_and_U14 ( .A(Fresh[57]), .B(cell_1771_and_in[0]), 
        .Z(cell_1771_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1771_a_HPC2_and_U13 ( .A(Fresh[57]), .B(cell_1771_and_in[1]), 
        .Z(cell_1771_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1771_a_HPC2_and_U12 ( .A1(cell_1771_a_HPC2_and_a_reg[1]), .A2(
        cell_1771_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1771_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1771_a_HPC2_and_U11 ( .A1(cell_1771_a_HPC2_and_a_reg[0]), .A2(
        cell_1771_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1771_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1771_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1771_a_HPC2_and_n9), 
        .ZN(cell_1771_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1771_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1771_a_HPC2_and_n9), 
        .ZN(cell_1771_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1771_a_HPC2_and_U8 ( .A(Fresh[57]), .ZN(cell_1771_a_HPC2_and_n9)
         );
  AND2_X1 cell_1771_a_HPC2_and_U7 ( .A1(cell_1771_and_in[1]), .A2(n414), .ZN(
        cell_1771_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1771_a_HPC2_and_U6 ( .A1(cell_1771_and_in[0]), .A2(n397), .ZN(
        cell_1771_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1771_a_HPC2_and_U5 ( .A(cell_1771_a_HPC2_and_n8), .B(
        cell_1771_a_HPC2_and_z_1__1_), .ZN(cell_1771_and_out[1]) );
  XNOR2_X1 cell_1771_a_HPC2_and_U4 ( .A(
        cell_1771_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1771_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1771_a_HPC2_and_n8) );
  XNOR2_X1 cell_1771_a_HPC2_and_U3 ( .A(cell_1771_a_HPC2_and_n7), .B(
        cell_1771_a_HPC2_and_z_0__0_), .ZN(cell_1771_and_out[0]) );
  XNOR2_X1 cell_1771_a_HPC2_and_U2 ( .A(
        cell_1771_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1771_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1771_a_HPC2_and_n7) );
  DFF_X1 cell_1771_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1771_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1771_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1771_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1771_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1771_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1771_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1771_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1771_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1771_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1772_U4 ( .A(1'b0), .B(cell_1772_and_out[1]), .Z(signal_3478)
         );
  XOR2_X1 cell_1772_U3 ( .A(1'b0), .B(cell_1772_and_out[0]), .Z(signal_2040)
         );
  XOR2_X1 cell_1772_U2 ( .A(1'b0), .B(n367), .Z(cell_1772_and_in[1]) );
  XOR2_X1 cell_1772_U1 ( .A(1'b0), .B(n366), .Z(cell_1772_and_in[0]) );
  XOR2_X1 cell_1772_a_HPC2_and_U14 ( .A(Fresh[58]), .B(cell_1772_and_in[0]), 
        .Z(cell_1772_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1772_a_HPC2_and_U13 ( .A(Fresh[58]), .B(cell_1772_and_in[1]), 
        .Z(cell_1772_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1772_a_HPC2_and_U12 ( .A1(cell_1772_a_HPC2_and_a_reg[1]), .A2(
        cell_1772_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1772_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1772_a_HPC2_and_U11 ( .A1(cell_1772_a_HPC2_and_a_reg[0]), .A2(
        cell_1772_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1772_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1772_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1772_a_HPC2_and_n9), 
        .ZN(cell_1772_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1772_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1772_a_HPC2_and_n9), 
        .ZN(cell_1772_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1772_a_HPC2_and_U8 ( .A(Fresh[58]), .ZN(cell_1772_a_HPC2_and_n9)
         );
  AND2_X1 cell_1772_a_HPC2_and_U7 ( .A1(cell_1772_and_in[1]), .A2(n425), .ZN(
        cell_1772_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1772_a_HPC2_and_U6 ( .A1(cell_1772_and_in[0]), .A2(n408), .ZN(
        cell_1772_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1772_a_HPC2_and_U5 ( .A(cell_1772_a_HPC2_and_n8), .B(
        cell_1772_a_HPC2_and_z_1__1_), .ZN(cell_1772_and_out[1]) );
  XNOR2_X1 cell_1772_a_HPC2_and_U4 ( .A(
        cell_1772_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1772_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1772_a_HPC2_and_n8) );
  XNOR2_X1 cell_1772_a_HPC2_and_U3 ( .A(cell_1772_a_HPC2_and_n7), .B(
        cell_1772_a_HPC2_and_z_0__0_), .ZN(cell_1772_and_out[0]) );
  XNOR2_X1 cell_1772_a_HPC2_and_U2 ( .A(
        cell_1772_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1772_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1772_a_HPC2_and_n7) );
  DFF_X1 cell_1772_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1772_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1772_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1772_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1772_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1772_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1772_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1772_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1772_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1772_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1773_U4 ( .A(n389), .B(cell_1773_and_out[1]), .Z(signal_3479)
         );
  XOR2_X1 cell_1773_U3 ( .A(n388), .B(cell_1773_and_out[0]), .Z(signal_2041)
         );
  XOR2_X1 cell_1773_U2 ( .A(n389), .B(n357), .Z(cell_1773_and_in[1]) );
  XOR2_X1 cell_1773_U1 ( .A(n388), .B(n356), .Z(cell_1773_and_in[0]) );
  XOR2_X1 cell_1773_a_HPC2_and_U14 ( .A(Fresh[59]), .B(cell_1773_and_in[0]), 
        .Z(cell_1773_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1773_a_HPC2_and_U13 ( .A(Fresh[59]), .B(cell_1773_and_in[1]), 
        .Z(cell_1773_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1773_a_HPC2_and_U12 ( .A1(cell_1773_a_HPC2_and_a_reg[1]), .A2(
        cell_1773_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1773_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1773_a_HPC2_and_U11 ( .A1(cell_1773_a_HPC2_and_a_reg[0]), .A2(
        cell_1773_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1773_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1773_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1773_a_HPC2_and_n9), 
        .ZN(cell_1773_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1773_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1773_a_HPC2_and_n9), 
        .ZN(cell_1773_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1773_a_HPC2_and_U8 ( .A(Fresh[59]), .ZN(cell_1773_a_HPC2_and_n9)
         );
  AND2_X1 cell_1773_a_HPC2_and_U7 ( .A1(cell_1773_and_in[1]), .A2(n414), .ZN(
        cell_1773_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1773_a_HPC2_and_U6 ( .A1(cell_1773_and_in[0]), .A2(n397), .ZN(
        cell_1773_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1773_a_HPC2_and_U5 ( .A(cell_1773_a_HPC2_and_n8), .B(
        cell_1773_a_HPC2_and_z_1__1_), .ZN(cell_1773_and_out[1]) );
  XNOR2_X1 cell_1773_a_HPC2_and_U4 ( .A(
        cell_1773_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1773_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1773_a_HPC2_and_n8) );
  XNOR2_X1 cell_1773_a_HPC2_and_U3 ( .A(cell_1773_a_HPC2_and_n7), .B(
        cell_1773_a_HPC2_and_z_0__0_), .ZN(cell_1773_and_out[0]) );
  XNOR2_X1 cell_1773_a_HPC2_and_U2 ( .A(
        cell_1773_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1773_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1773_a_HPC2_and_n7) );
  DFF_X1 cell_1773_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1773_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1773_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1773_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1773_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1773_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1773_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1773_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1773_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1773_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1774_U4 ( .A(n355), .B(1'b0), .Z(cell_1774_and_in[1]) );
  XOR2_X1 cell_1774_U3 ( .A(n353), .B(1'b0), .Z(cell_1774_and_in[0]) );
  XOR2_X2 cell_1774_U2 ( .A(n355), .B(cell_1774_and_out[1]), .Z(signal_3480)
         );
  XOR2_X2 cell_1774_U1 ( .A(n353), .B(cell_1774_and_out[0]), .Z(signal_2042)
         );
  XOR2_X1 cell_1774_a_HPC2_and_U14 ( .A(Fresh[60]), .B(cell_1774_and_in[0]), 
        .Z(cell_1774_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1774_a_HPC2_and_U13 ( .A(Fresh[60]), .B(cell_1774_and_in[1]), 
        .Z(cell_1774_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1774_a_HPC2_and_U12 ( .A1(cell_1774_a_HPC2_and_a_reg[1]), .A2(
        cell_1774_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1774_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1774_a_HPC2_and_U11 ( .A1(cell_1774_a_HPC2_and_a_reg[0]), .A2(
        cell_1774_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1774_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1774_a_HPC2_and_U10 ( .A1(signal_3237), .A2(
        cell_1774_a_HPC2_and_n9), .ZN(cell_1774_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1774_a_HPC2_and_U9 ( .A1(signal_1512), .A2(
        cell_1774_a_HPC2_and_n9), .ZN(cell_1774_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1774_a_HPC2_and_U8 ( .A(Fresh[60]), .ZN(cell_1774_a_HPC2_and_n9)
         );
  AND2_X1 cell_1774_a_HPC2_and_U7 ( .A1(cell_1774_and_in[1]), .A2(signal_3237), 
        .ZN(cell_1774_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1774_a_HPC2_and_U6 ( .A1(cell_1774_and_in[0]), .A2(signal_1512), 
        .ZN(cell_1774_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1774_a_HPC2_and_U5 ( .A(cell_1774_a_HPC2_and_n8), .B(
        cell_1774_a_HPC2_and_z_1__1_), .ZN(cell_1774_and_out[1]) );
  XNOR2_X1 cell_1774_a_HPC2_and_U4 ( .A(
        cell_1774_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1774_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1774_a_HPC2_and_n8) );
  XNOR2_X1 cell_1774_a_HPC2_and_U3 ( .A(cell_1774_a_HPC2_and_n7), .B(
        cell_1774_a_HPC2_and_z_0__0_), .ZN(cell_1774_and_out[0]) );
  XNOR2_X1 cell_1774_a_HPC2_and_U2 ( .A(
        cell_1774_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1774_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1774_a_HPC2_and_n7) );
  DFF_X1 cell_1774_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1774_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1774_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1512), 
        .CK(clk), .Q(cell_1774_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1774_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1774_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3237), 
        .CK(clk), .Q(cell_1774_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1774_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1774_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1774_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1775_U4 ( .A(n370), .B(cell_1775_and_out[1]), .Z(signal_3481)
         );
  XOR2_X1 cell_1775_U3 ( .A(n368), .B(cell_1775_and_out[0]), .Z(signal_2043)
         );
  XOR2_X1 cell_1775_U2 ( .A(n370), .B(n387), .Z(cell_1775_and_in[1]) );
  XOR2_X1 cell_1775_U1 ( .A(n368), .B(n385), .Z(cell_1775_and_in[0]) );
  XOR2_X1 cell_1775_a_HPC2_and_U14 ( .A(Fresh[61]), .B(cell_1775_and_in[0]), 
        .Z(cell_1775_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1775_a_HPC2_and_U13 ( .A(Fresh[61]), .B(cell_1775_and_in[1]), 
        .Z(cell_1775_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1775_a_HPC2_and_U12 ( .A1(cell_1775_a_HPC2_and_a_reg[1]), .A2(
        cell_1775_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1775_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1775_a_HPC2_and_U11 ( .A1(cell_1775_a_HPC2_and_a_reg[0]), .A2(
        cell_1775_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1775_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1775_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1775_a_HPC2_and_n9), 
        .ZN(cell_1775_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1775_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1775_a_HPC2_and_n9), 
        .ZN(cell_1775_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1775_a_HPC2_and_U8 ( .A(Fresh[61]), .ZN(cell_1775_a_HPC2_and_n9)
         );
  AND2_X1 cell_1775_a_HPC2_and_U7 ( .A1(cell_1775_and_in[1]), .A2(n414), .ZN(
        cell_1775_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1775_a_HPC2_and_U6 ( .A1(cell_1775_and_in[0]), .A2(n397), .ZN(
        cell_1775_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1775_a_HPC2_and_U5 ( .A(cell_1775_a_HPC2_and_n8), .B(
        cell_1775_a_HPC2_and_z_1__1_), .ZN(cell_1775_and_out[1]) );
  XNOR2_X1 cell_1775_a_HPC2_and_U4 ( .A(
        cell_1775_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1775_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1775_a_HPC2_and_n8) );
  XNOR2_X1 cell_1775_a_HPC2_and_U3 ( .A(cell_1775_a_HPC2_and_n7), .B(
        cell_1775_a_HPC2_and_z_0__0_), .ZN(cell_1775_and_out[0]) );
  XNOR2_X1 cell_1775_a_HPC2_and_U2 ( .A(
        cell_1775_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1775_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1775_a_HPC2_and_n7) );
  DFF_X1 cell_1775_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1775_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1775_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1775_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1775_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1775_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1775_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1775_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1775_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1775_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1776_U4 ( .A(n381), .B(cell_1776_and_out[1]), .Z(signal_3482)
         );
  XOR2_X1 cell_1776_U3 ( .A(n380), .B(cell_1776_and_out[0]), .Z(signal_2044)
         );
  XOR2_X1 cell_1776_U2 ( .A(n381), .B(n379), .Z(cell_1776_and_in[1]) );
  XOR2_X1 cell_1776_U1 ( .A(n380), .B(n377), .Z(cell_1776_and_in[0]) );
  XOR2_X1 cell_1776_a_HPC2_and_U14 ( .A(Fresh[62]), .B(cell_1776_and_in[0]), 
        .Z(cell_1776_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1776_a_HPC2_and_U13 ( .A(Fresh[62]), .B(cell_1776_and_in[1]), 
        .Z(cell_1776_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1776_a_HPC2_and_U12 ( .A1(cell_1776_a_HPC2_and_a_reg[1]), .A2(
        cell_1776_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1776_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1776_a_HPC2_and_U11 ( .A1(cell_1776_a_HPC2_and_a_reg[0]), .A2(
        cell_1776_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1776_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1776_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1776_a_HPC2_and_n9), 
        .ZN(cell_1776_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1776_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1776_a_HPC2_and_n9), 
        .ZN(cell_1776_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1776_a_HPC2_and_U8 ( .A(Fresh[62]), .ZN(cell_1776_a_HPC2_and_n9)
         );
  AND2_X1 cell_1776_a_HPC2_and_U7 ( .A1(cell_1776_and_in[1]), .A2(n415), .ZN(
        cell_1776_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1776_a_HPC2_and_U6 ( .A1(cell_1776_and_in[0]), .A2(n398), .ZN(
        cell_1776_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1776_a_HPC2_and_U5 ( .A(cell_1776_a_HPC2_and_n8), .B(
        cell_1776_a_HPC2_and_z_1__1_), .ZN(cell_1776_and_out[1]) );
  XNOR2_X1 cell_1776_a_HPC2_and_U4 ( .A(
        cell_1776_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1776_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1776_a_HPC2_and_n8) );
  XNOR2_X1 cell_1776_a_HPC2_and_U3 ( .A(cell_1776_a_HPC2_and_n7), .B(
        cell_1776_a_HPC2_and_z_0__0_), .ZN(cell_1776_and_out[0]) );
  XNOR2_X1 cell_1776_a_HPC2_and_U2 ( .A(
        cell_1776_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1776_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1776_a_HPC2_and_n7) );
  DFF_X1 cell_1776_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1776_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1776_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1776_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1776_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1776_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1776_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1776_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1776_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1776_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1777_U4 ( .A(n374), .B(cell_1777_and_out[1]), .Z(signal_3483)
         );
  XOR2_X1 cell_1777_U3 ( .A(n372), .B(cell_1777_and_out[0]), .Z(signal_2045)
         );
  XOR2_X1 cell_1777_U2 ( .A(n374), .B(signal_3256), .Z(cell_1777_and_in[1]) );
  XOR2_X1 cell_1777_U1 ( .A(n372), .B(signal_1982), .Z(cell_1777_and_in[0]) );
  XOR2_X1 cell_1777_a_HPC2_and_U14 ( .A(Fresh[63]), .B(cell_1777_and_in[0]), 
        .Z(cell_1777_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1777_a_HPC2_and_U13 ( .A(Fresh[63]), .B(cell_1777_and_in[1]), 
        .Z(cell_1777_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1777_a_HPC2_and_U12 ( .A1(cell_1777_a_HPC2_and_a_reg[1]), .A2(
        cell_1777_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1777_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1777_a_HPC2_and_U11 ( .A1(cell_1777_a_HPC2_and_a_reg[0]), .A2(
        cell_1777_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1777_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1777_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1777_a_HPC2_and_n9), 
        .ZN(cell_1777_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1777_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1777_a_HPC2_and_n9), 
        .ZN(cell_1777_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1777_a_HPC2_and_U8 ( .A(Fresh[63]), .ZN(cell_1777_a_HPC2_and_n9)
         );
  AND2_X1 cell_1777_a_HPC2_and_U7 ( .A1(cell_1777_and_in[1]), .A2(n415), .ZN(
        cell_1777_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1777_a_HPC2_and_U6 ( .A1(cell_1777_and_in[0]), .A2(n398), .ZN(
        cell_1777_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1777_a_HPC2_and_U5 ( .A(cell_1777_a_HPC2_and_n8), .B(
        cell_1777_a_HPC2_and_z_1__1_), .ZN(cell_1777_and_out[1]) );
  XNOR2_X1 cell_1777_a_HPC2_and_U4 ( .A(
        cell_1777_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1777_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1777_a_HPC2_and_n8) );
  XNOR2_X1 cell_1777_a_HPC2_and_U3 ( .A(cell_1777_a_HPC2_and_n7), .B(
        cell_1777_a_HPC2_and_z_0__0_), .ZN(cell_1777_and_out[0]) );
  XNOR2_X1 cell_1777_a_HPC2_and_U2 ( .A(
        cell_1777_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1777_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1777_a_HPC2_and_n7) );
  DFF_X1 cell_1777_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1777_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1777_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1777_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1777_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1777_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1777_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1777_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1777_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1777_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1778_U4 ( .A(signal_3406), .B(cell_1778_and_out[1]), .Z(
        signal_3484) );
  XOR2_X1 cell_1778_U3 ( .A(signal_1992), .B(cell_1778_and_out[0]), .Z(
        signal_2046) );
  XOR2_X1 cell_1778_U2 ( .A(signal_3406), .B(n357), .Z(cell_1778_and_in[1]) );
  XOR2_X1 cell_1778_U1 ( .A(signal_1992), .B(n356), .Z(cell_1778_and_in[0]) );
  XOR2_X1 cell_1778_a_HPC2_and_U14 ( .A(Fresh[64]), .B(cell_1778_and_in[0]), 
        .Z(cell_1778_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1778_a_HPC2_and_U13 ( .A(Fresh[64]), .B(cell_1778_and_in[1]), 
        .Z(cell_1778_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1778_a_HPC2_and_U12 ( .A1(cell_1778_a_HPC2_and_a_reg[1]), .A2(
        cell_1778_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1778_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1778_a_HPC2_and_U11 ( .A1(cell_1778_a_HPC2_and_a_reg[0]), .A2(
        cell_1778_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1778_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1778_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1778_a_HPC2_and_n9), 
        .ZN(cell_1778_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1778_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1778_a_HPC2_and_n9), 
        .ZN(cell_1778_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1778_a_HPC2_and_U8 ( .A(Fresh[64]), .ZN(cell_1778_a_HPC2_and_n9)
         );
  AND2_X1 cell_1778_a_HPC2_and_U7 ( .A1(cell_1778_and_in[1]), .A2(n423), .ZN(
        cell_1778_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1778_a_HPC2_and_U6 ( .A1(cell_1778_and_in[0]), .A2(n406), .ZN(
        cell_1778_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1778_a_HPC2_and_U5 ( .A(cell_1778_a_HPC2_and_n8), .B(
        cell_1778_a_HPC2_and_z_1__1_), .ZN(cell_1778_and_out[1]) );
  XNOR2_X1 cell_1778_a_HPC2_and_U4 ( .A(
        cell_1778_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1778_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1778_a_HPC2_and_n8) );
  XNOR2_X1 cell_1778_a_HPC2_and_U3 ( .A(cell_1778_a_HPC2_and_n7), .B(
        cell_1778_a_HPC2_and_z_0__0_), .ZN(cell_1778_and_out[0]) );
  XNOR2_X1 cell_1778_a_HPC2_and_U2 ( .A(
        cell_1778_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1778_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1778_a_HPC2_and_n7) );
  DFF_X1 cell_1778_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1778_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1778_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1778_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1778_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1778_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1778_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1778_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1778_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1778_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1779_U4 ( .A(1'b0), .B(cell_1779_and_out[1]), .Z(signal_3485)
         );
  XOR2_X1 cell_1779_U3 ( .A(1'b0), .B(cell_1779_and_out[0]), .Z(signal_2047)
         );
  XOR2_X1 cell_1779_U2 ( .A(1'b0), .B(n379), .Z(cell_1779_and_in[1]) );
  XOR2_X1 cell_1779_U1 ( .A(1'b0), .B(n377), .Z(cell_1779_and_in[0]) );
  XOR2_X1 cell_1779_a_HPC2_and_U14 ( .A(Fresh[65]), .B(cell_1779_and_in[0]), 
        .Z(cell_1779_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1779_a_HPC2_and_U13 ( .A(Fresh[65]), .B(cell_1779_and_in[1]), 
        .Z(cell_1779_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1779_a_HPC2_and_U12 ( .A1(cell_1779_a_HPC2_and_a_reg[1]), .A2(
        cell_1779_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1779_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1779_a_HPC2_and_U11 ( .A1(cell_1779_a_HPC2_and_a_reg[0]), .A2(
        cell_1779_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1779_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1779_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1779_a_HPC2_and_n9), 
        .ZN(cell_1779_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1779_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1779_a_HPC2_and_n9), 
        .ZN(cell_1779_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1779_a_HPC2_and_U8 ( .A(Fresh[65]), .ZN(cell_1779_a_HPC2_and_n9)
         );
  AND2_X1 cell_1779_a_HPC2_and_U7 ( .A1(cell_1779_and_in[1]), .A2(n424), .ZN(
        cell_1779_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1779_a_HPC2_and_U6 ( .A1(cell_1779_and_in[0]), .A2(n407), .ZN(
        cell_1779_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1779_a_HPC2_and_U5 ( .A(cell_1779_a_HPC2_and_n8), .B(
        cell_1779_a_HPC2_and_z_1__1_), .ZN(cell_1779_and_out[1]) );
  XNOR2_X1 cell_1779_a_HPC2_and_U4 ( .A(
        cell_1779_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1779_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1779_a_HPC2_and_n8) );
  XNOR2_X1 cell_1779_a_HPC2_and_U3 ( .A(cell_1779_a_HPC2_and_n7), .B(
        cell_1779_a_HPC2_and_z_0__0_), .ZN(cell_1779_and_out[0]) );
  XNOR2_X1 cell_1779_a_HPC2_and_U2 ( .A(
        cell_1779_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1779_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1779_a_HPC2_and_n7) );
  DFF_X1 cell_1779_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1779_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1779_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1779_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1779_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1779_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1779_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1779_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1779_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1779_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1780_U4 ( .A(n389), .B(cell_1780_and_out[1]), .Z(signal_3486)
         );
  XOR2_X1 cell_1780_U3 ( .A(n388), .B(cell_1780_and_out[0]), .Z(signal_2048)
         );
  XOR2_X1 cell_1780_U2 ( .A(n389), .B(signal_3406), .Z(cell_1780_and_in[1]) );
  XOR2_X1 cell_1780_U1 ( .A(n388), .B(signal_1992), .Z(cell_1780_and_in[0]) );
  XOR2_X1 cell_1780_a_HPC2_and_U14 ( .A(Fresh[66]), .B(cell_1780_and_in[0]), 
        .Z(cell_1780_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1780_a_HPC2_and_U13 ( .A(Fresh[66]), .B(cell_1780_and_in[1]), 
        .Z(cell_1780_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1780_a_HPC2_and_U12 ( .A1(cell_1780_a_HPC2_and_a_reg[1]), .A2(
        cell_1780_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1780_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1780_a_HPC2_and_U11 ( .A1(cell_1780_a_HPC2_and_a_reg[0]), .A2(
        cell_1780_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1780_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1780_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1780_a_HPC2_and_n9), 
        .ZN(cell_1780_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1780_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1780_a_HPC2_and_n9), 
        .ZN(cell_1780_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1780_a_HPC2_and_U8 ( .A(Fresh[66]), .ZN(cell_1780_a_HPC2_and_n9)
         );
  AND2_X1 cell_1780_a_HPC2_and_U7 ( .A1(cell_1780_and_in[1]), .A2(n415), .ZN(
        cell_1780_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1780_a_HPC2_and_U6 ( .A1(cell_1780_and_in[0]), .A2(n398), .ZN(
        cell_1780_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1780_a_HPC2_and_U5 ( .A(cell_1780_a_HPC2_and_n8), .B(
        cell_1780_a_HPC2_and_z_1__1_), .ZN(cell_1780_and_out[1]) );
  XNOR2_X1 cell_1780_a_HPC2_and_U4 ( .A(
        cell_1780_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1780_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1780_a_HPC2_and_n8) );
  XNOR2_X1 cell_1780_a_HPC2_and_U3 ( .A(cell_1780_a_HPC2_and_n7), .B(
        cell_1780_a_HPC2_and_z_0__0_), .ZN(cell_1780_and_out[0]) );
  XNOR2_X1 cell_1780_a_HPC2_and_U2 ( .A(
        cell_1780_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1780_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1780_a_HPC2_and_n7) );
  DFF_X1 cell_1780_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1780_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1780_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1780_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1780_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1780_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1780_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1780_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1780_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1780_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1781_U4 ( .A(n374), .B(cell_1781_and_out[1]), .Z(signal_3487)
         );
  XOR2_X1 cell_1781_U3 ( .A(n372), .B(cell_1781_and_out[0]), .Z(signal_2049)
         );
  XOR2_X1 cell_1781_U2 ( .A(n374), .B(signal_3406), .Z(cell_1781_and_in[1]) );
  XOR2_X1 cell_1781_U1 ( .A(n372), .B(signal_1992), .Z(cell_1781_and_in[0]) );
  XOR2_X1 cell_1781_a_HPC2_and_U14 ( .A(Fresh[67]), .B(cell_1781_and_in[0]), 
        .Z(cell_1781_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1781_a_HPC2_and_U13 ( .A(Fresh[67]), .B(cell_1781_and_in[1]), 
        .Z(cell_1781_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1781_a_HPC2_and_U12 ( .A1(cell_1781_a_HPC2_and_a_reg[1]), .A2(
        cell_1781_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1781_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1781_a_HPC2_and_U11 ( .A1(cell_1781_a_HPC2_and_a_reg[0]), .A2(
        cell_1781_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1781_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1781_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1781_a_HPC2_and_n9), 
        .ZN(cell_1781_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1781_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1781_a_HPC2_and_n9), 
        .ZN(cell_1781_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1781_a_HPC2_and_U8 ( .A(Fresh[67]), .ZN(cell_1781_a_HPC2_and_n9)
         );
  AND2_X1 cell_1781_a_HPC2_and_U7 ( .A1(cell_1781_and_in[1]), .A2(n415), .ZN(
        cell_1781_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1781_a_HPC2_and_U6 ( .A1(cell_1781_and_in[0]), .A2(n398), .ZN(
        cell_1781_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1781_a_HPC2_and_U5 ( .A(cell_1781_a_HPC2_and_n8), .B(
        cell_1781_a_HPC2_and_z_1__1_), .ZN(cell_1781_and_out[1]) );
  XNOR2_X1 cell_1781_a_HPC2_and_U4 ( .A(
        cell_1781_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1781_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1781_a_HPC2_and_n8) );
  XNOR2_X1 cell_1781_a_HPC2_and_U3 ( .A(cell_1781_a_HPC2_and_n7), .B(
        cell_1781_a_HPC2_and_z_0__0_), .ZN(cell_1781_and_out[0]) );
  XNOR2_X1 cell_1781_a_HPC2_and_U2 ( .A(
        cell_1781_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1781_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1781_a_HPC2_and_n7) );
  DFF_X1 cell_1781_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1781_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1781_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1781_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1781_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1781_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1781_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1781_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1781_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1781_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1782_U4 ( .A(n365), .B(cell_1782_and_out[1]), .Z(signal_3488)
         );
  XOR2_X1 cell_1782_U3 ( .A(n363), .B(cell_1782_and_out[0]), .Z(signal_2050)
         );
  XOR2_X1 cell_1782_U2 ( .A(n365), .B(signal_3256), .Z(cell_1782_and_in[1]) );
  XOR2_X1 cell_1782_U1 ( .A(n363), .B(signal_1982), .Z(cell_1782_and_in[0]) );
  XOR2_X1 cell_1782_a_HPC2_and_U14 ( .A(Fresh[68]), .B(cell_1782_and_in[0]), 
        .Z(cell_1782_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1782_a_HPC2_and_U13 ( .A(Fresh[68]), .B(cell_1782_and_in[1]), 
        .Z(cell_1782_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1782_a_HPC2_and_U12 ( .A1(cell_1782_a_HPC2_and_a_reg[1]), .A2(
        cell_1782_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1782_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1782_a_HPC2_and_U11 ( .A1(cell_1782_a_HPC2_and_a_reg[0]), .A2(
        cell_1782_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1782_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1782_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1782_a_HPC2_and_n9), 
        .ZN(cell_1782_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1782_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1782_a_HPC2_and_n9), 
        .ZN(cell_1782_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1782_a_HPC2_and_U8 ( .A(Fresh[68]), .ZN(cell_1782_a_HPC2_and_n9)
         );
  AND2_X1 cell_1782_a_HPC2_and_U7 ( .A1(cell_1782_and_in[1]), .A2(n415), .ZN(
        cell_1782_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1782_a_HPC2_and_U6 ( .A1(cell_1782_and_in[0]), .A2(n398), .ZN(
        cell_1782_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1782_a_HPC2_and_U5 ( .A(cell_1782_a_HPC2_and_n8), .B(
        cell_1782_a_HPC2_and_z_1__1_), .ZN(cell_1782_and_out[1]) );
  XNOR2_X1 cell_1782_a_HPC2_and_U4 ( .A(
        cell_1782_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1782_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1782_a_HPC2_and_n8) );
  XNOR2_X1 cell_1782_a_HPC2_and_U3 ( .A(cell_1782_a_HPC2_and_n7), .B(
        cell_1782_a_HPC2_and_z_0__0_), .ZN(cell_1782_and_out[0]) );
  XNOR2_X1 cell_1782_a_HPC2_and_U2 ( .A(
        cell_1782_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1782_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1782_a_HPC2_and_n7) );
  DFF_X1 cell_1782_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1782_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1782_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1782_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1782_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1782_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1782_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1782_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1782_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1782_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1783_U4 ( .A(1'b0), .B(cell_1783_and_out[1]), .Z(signal_3489)
         );
  XOR2_X1 cell_1783_U3 ( .A(1'b0), .B(cell_1783_and_out[0]), .Z(signal_2051)
         );
  XOR2_X1 cell_1783_U2 ( .A(1'b0), .B(n355), .Z(cell_1783_and_in[1]) );
  XOR2_X1 cell_1783_U1 ( .A(1'b0), .B(n353), .Z(cell_1783_and_in[0]) );
  XOR2_X1 cell_1783_a_HPC2_and_U14 ( .A(Fresh[69]), .B(cell_1783_and_in[0]), 
        .Z(cell_1783_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1783_a_HPC2_and_U13 ( .A(Fresh[69]), .B(cell_1783_and_in[1]), 
        .Z(cell_1783_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1783_a_HPC2_and_U12 ( .A1(cell_1783_a_HPC2_and_a_reg[1]), .A2(
        cell_1783_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1783_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1783_a_HPC2_and_U11 ( .A1(cell_1783_a_HPC2_and_a_reg[0]), .A2(
        cell_1783_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1783_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1783_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1783_a_HPC2_and_n9), 
        .ZN(cell_1783_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1783_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1783_a_HPC2_and_n9), 
        .ZN(cell_1783_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1783_a_HPC2_and_U8 ( .A(Fresh[69]), .ZN(cell_1783_a_HPC2_and_n9)
         );
  AND2_X1 cell_1783_a_HPC2_and_U7 ( .A1(cell_1783_and_in[1]), .A2(n427), .ZN(
        cell_1783_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1783_a_HPC2_and_U6 ( .A1(cell_1783_and_in[0]), .A2(n410), .ZN(
        cell_1783_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1783_a_HPC2_and_U5 ( .A(cell_1783_a_HPC2_and_n8), .B(
        cell_1783_a_HPC2_and_z_1__1_), .ZN(cell_1783_and_out[1]) );
  XNOR2_X1 cell_1783_a_HPC2_and_U4 ( .A(
        cell_1783_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1783_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1783_a_HPC2_and_n8) );
  XNOR2_X1 cell_1783_a_HPC2_and_U3 ( .A(cell_1783_a_HPC2_and_n7), .B(
        cell_1783_a_HPC2_and_z_0__0_), .ZN(cell_1783_and_out[0]) );
  XNOR2_X1 cell_1783_a_HPC2_and_U2 ( .A(
        cell_1783_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1783_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1783_a_HPC2_and_n7) );
  DFF_X1 cell_1783_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1783_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1783_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1783_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1783_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1783_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1783_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1783_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1783_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1783_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1784_U4 ( .A(n389), .B(cell_1784_and_out[1]), .Z(signal_3490)
         );
  XOR2_X1 cell_1784_U3 ( .A(n388), .B(cell_1784_and_out[0]), .Z(signal_2052)
         );
  XOR2_X1 cell_1784_U2 ( .A(n389), .B(n365), .Z(cell_1784_and_in[1]) );
  XOR2_X1 cell_1784_U1 ( .A(n388), .B(n363), .Z(cell_1784_and_in[0]) );
  XOR2_X1 cell_1784_a_HPC2_and_U14 ( .A(Fresh[70]), .B(cell_1784_and_in[0]), 
        .Z(cell_1784_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1784_a_HPC2_and_U13 ( .A(Fresh[70]), .B(cell_1784_and_in[1]), 
        .Z(cell_1784_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1784_a_HPC2_and_U12 ( .A1(cell_1784_a_HPC2_and_a_reg[1]), .A2(
        cell_1784_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1784_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1784_a_HPC2_and_U11 ( .A1(cell_1784_a_HPC2_and_a_reg[0]), .A2(
        cell_1784_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1784_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1784_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1784_a_HPC2_and_n9), 
        .ZN(cell_1784_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1784_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1784_a_HPC2_and_n9), 
        .ZN(cell_1784_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1784_a_HPC2_and_U8 ( .A(Fresh[70]), .ZN(cell_1784_a_HPC2_and_n9)
         );
  AND2_X1 cell_1784_a_HPC2_and_U7 ( .A1(cell_1784_and_in[1]), .A2(n415), .ZN(
        cell_1784_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1784_a_HPC2_and_U6 ( .A1(cell_1784_and_in[0]), .A2(n398), .ZN(
        cell_1784_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1784_a_HPC2_and_U5 ( .A(cell_1784_a_HPC2_and_n8), .B(
        cell_1784_a_HPC2_and_z_1__1_), .ZN(cell_1784_and_out[1]) );
  XNOR2_X1 cell_1784_a_HPC2_and_U4 ( .A(
        cell_1784_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1784_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1784_a_HPC2_and_n8) );
  XNOR2_X1 cell_1784_a_HPC2_and_U3 ( .A(cell_1784_a_HPC2_and_n7), .B(
        cell_1784_a_HPC2_and_z_0__0_), .ZN(cell_1784_and_out[0]) );
  XNOR2_X1 cell_1784_a_HPC2_and_U2 ( .A(
        cell_1784_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1784_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1784_a_HPC2_and_n7) );
  DFF_X1 cell_1784_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1784_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1784_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1784_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1784_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1784_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1784_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1784_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1784_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1784_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1785_U4 ( .A(1'b0), .B(cell_1785_and_out[1]), .Z(signal_3491)
         );
  XOR2_X1 cell_1785_U3 ( .A(1'b0), .B(cell_1785_and_out[0]), .Z(signal_2053)
         );
  XOR2_X1 cell_1785_U2 ( .A(1'b0), .B(signal_3406), .Z(cell_1785_and_in[1]) );
  XOR2_X1 cell_1785_U1 ( .A(1'b0), .B(signal_1992), .Z(cell_1785_and_in[0]) );
  XOR2_X1 cell_1785_a_HPC2_and_U14 ( .A(Fresh[71]), .B(cell_1785_and_in[0]), 
        .Z(cell_1785_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1785_a_HPC2_and_U13 ( .A(Fresh[71]), .B(cell_1785_and_in[1]), 
        .Z(cell_1785_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1785_a_HPC2_and_U12 ( .A1(cell_1785_a_HPC2_and_a_reg[1]), .A2(
        cell_1785_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1785_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1785_a_HPC2_and_U11 ( .A1(cell_1785_a_HPC2_and_a_reg[0]), .A2(
        cell_1785_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1785_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1785_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1785_a_HPC2_and_n9), 
        .ZN(cell_1785_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1785_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1785_a_HPC2_and_n9), 
        .ZN(cell_1785_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1785_a_HPC2_and_U8 ( .A(Fresh[71]), .ZN(cell_1785_a_HPC2_and_n9)
         );
  AND2_X1 cell_1785_a_HPC2_and_U7 ( .A1(cell_1785_and_in[1]), .A2(n413), .ZN(
        cell_1785_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1785_a_HPC2_and_U6 ( .A1(cell_1785_and_in[0]), .A2(n396), .ZN(
        cell_1785_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1785_a_HPC2_and_U5 ( .A(cell_1785_a_HPC2_and_n8), .B(
        cell_1785_a_HPC2_and_z_1__1_), .ZN(cell_1785_and_out[1]) );
  XNOR2_X1 cell_1785_a_HPC2_and_U4 ( .A(
        cell_1785_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1785_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1785_a_HPC2_and_n8) );
  XNOR2_X1 cell_1785_a_HPC2_and_U3 ( .A(cell_1785_a_HPC2_and_n7), .B(
        cell_1785_a_HPC2_and_z_0__0_), .ZN(cell_1785_and_out[0]) );
  XNOR2_X1 cell_1785_a_HPC2_and_U2 ( .A(
        cell_1785_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1785_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1785_a_HPC2_and_n7) );
  DFF_X1 cell_1785_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1785_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1785_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1785_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1785_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1785_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1785_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1785_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1785_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1785_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1786_U4 ( .A(n381), .B(cell_1786_and_out[1]), .Z(signal_3492)
         );
  XOR2_X1 cell_1786_U3 ( .A(n380), .B(cell_1786_and_out[0]), .Z(signal_2054)
         );
  XOR2_X1 cell_1786_U2 ( .A(n381), .B(signal_3406), .Z(cell_1786_and_in[1]) );
  XOR2_X1 cell_1786_U1 ( .A(n380), .B(signal_1992), .Z(cell_1786_and_in[0]) );
  XOR2_X1 cell_1786_a_HPC2_and_U14 ( .A(Fresh[72]), .B(cell_1786_and_in[0]), 
        .Z(cell_1786_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1786_a_HPC2_and_U13 ( .A(Fresh[72]), .B(cell_1786_and_in[1]), 
        .Z(cell_1786_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1786_a_HPC2_and_U12 ( .A1(cell_1786_a_HPC2_and_a_reg[1]), .A2(
        cell_1786_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1786_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1786_a_HPC2_and_U11 ( .A1(cell_1786_a_HPC2_and_a_reg[0]), .A2(
        cell_1786_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1786_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1786_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1786_a_HPC2_and_n9), 
        .ZN(cell_1786_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1786_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1786_a_HPC2_and_n9), 
        .ZN(cell_1786_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1786_a_HPC2_and_U8 ( .A(Fresh[72]), .ZN(cell_1786_a_HPC2_and_n9)
         );
  AND2_X1 cell_1786_a_HPC2_and_U7 ( .A1(cell_1786_and_in[1]), .A2(n415), .ZN(
        cell_1786_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1786_a_HPC2_and_U6 ( .A1(cell_1786_and_in[0]), .A2(n398), .ZN(
        cell_1786_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1786_a_HPC2_and_U5 ( .A(cell_1786_a_HPC2_and_n8), .B(
        cell_1786_a_HPC2_and_z_1__1_), .ZN(cell_1786_and_out[1]) );
  XNOR2_X1 cell_1786_a_HPC2_and_U4 ( .A(
        cell_1786_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1786_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1786_a_HPC2_and_n8) );
  XNOR2_X1 cell_1786_a_HPC2_and_U3 ( .A(cell_1786_a_HPC2_and_n7), .B(
        cell_1786_a_HPC2_and_z_0__0_), .ZN(cell_1786_and_out[0]) );
  XNOR2_X1 cell_1786_a_HPC2_and_U2 ( .A(
        cell_1786_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1786_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1786_a_HPC2_and_n7) );
  DFF_X1 cell_1786_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1786_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1786_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1786_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1786_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1786_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1786_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1786_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1786_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1786_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1787_U4 ( .A(n357), .B(cell_1787_and_out[1]), .Z(signal_3493)
         );
  XOR2_X1 cell_1787_U3 ( .A(signal_2013), .B(cell_1787_and_out[0]), .Z(
        signal_2055) );
  XOR2_X1 cell_1787_U2 ( .A(n357), .B(n383), .Z(cell_1787_and_in[1]) );
  XOR2_X1 cell_1787_U1 ( .A(signal_2013), .B(n382), .Z(cell_1787_and_in[0]) );
  XOR2_X1 cell_1787_a_HPC2_and_U14 ( .A(Fresh[73]), .B(cell_1787_and_in[0]), 
        .Z(cell_1787_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1787_a_HPC2_and_U13 ( .A(Fresh[73]), .B(cell_1787_and_in[1]), 
        .Z(cell_1787_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1787_a_HPC2_and_U12 ( .A1(cell_1787_a_HPC2_and_a_reg[1]), .A2(
        cell_1787_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1787_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1787_a_HPC2_and_U11 ( .A1(cell_1787_a_HPC2_and_a_reg[0]), .A2(
        cell_1787_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1787_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1787_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1787_a_HPC2_and_n9), 
        .ZN(cell_1787_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1787_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1787_a_HPC2_and_n9), 
        .ZN(cell_1787_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1787_a_HPC2_and_U8 ( .A(Fresh[73]), .ZN(cell_1787_a_HPC2_and_n9)
         );
  AND2_X1 cell_1787_a_HPC2_and_U7 ( .A1(cell_1787_and_in[1]), .A2(n416), .ZN(
        cell_1787_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1787_a_HPC2_and_U6 ( .A1(cell_1787_and_in[0]), .A2(n399), .ZN(
        cell_1787_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1787_a_HPC2_and_U5 ( .A(cell_1787_a_HPC2_and_n8), .B(
        cell_1787_a_HPC2_and_z_1__1_), .ZN(cell_1787_and_out[1]) );
  XNOR2_X1 cell_1787_a_HPC2_and_U4 ( .A(
        cell_1787_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1787_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1787_a_HPC2_and_n8) );
  XNOR2_X1 cell_1787_a_HPC2_and_U3 ( .A(cell_1787_a_HPC2_and_n7), .B(
        cell_1787_a_HPC2_and_z_0__0_), .ZN(cell_1787_and_out[0]) );
  XNOR2_X1 cell_1787_a_HPC2_and_U2 ( .A(
        cell_1787_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1787_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1787_a_HPC2_and_n7) );
  DFF_X1 cell_1787_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1787_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1787_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1787_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1787_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1787_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1787_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1787_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1787_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1787_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1788_U4 ( .A(n357), .B(cell_1788_and_out[1]), .Z(signal_3494)
         );
  XOR2_X1 cell_1788_U3 ( .A(n356), .B(cell_1788_and_out[0]), .Z(signal_2056)
         );
  XOR2_X1 cell_1788_U2 ( .A(n357), .B(n387), .Z(cell_1788_and_in[1]) );
  XOR2_X1 cell_1788_U1 ( .A(n356), .B(n385), .Z(cell_1788_and_in[0]) );
  XOR2_X1 cell_1788_a_HPC2_and_U14 ( .A(Fresh[74]), .B(cell_1788_and_in[0]), 
        .Z(cell_1788_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1788_a_HPC2_and_U13 ( .A(Fresh[74]), .B(cell_1788_and_in[1]), 
        .Z(cell_1788_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1788_a_HPC2_and_U12 ( .A1(cell_1788_a_HPC2_and_a_reg[1]), .A2(
        cell_1788_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1788_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1788_a_HPC2_and_U11 ( .A1(cell_1788_a_HPC2_and_a_reg[0]), .A2(
        cell_1788_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1788_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1788_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1788_a_HPC2_and_n9), 
        .ZN(cell_1788_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1788_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1788_a_HPC2_and_n9), 
        .ZN(cell_1788_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1788_a_HPC2_and_U8 ( .A(Fresh[74]), .ZN(cell_1788_a_HPC2_and_n9)
         );
  AND2_X1 cell_1788_a_HPC2_and_U7 ( .A1(cell_1788_and_in[1]), .A2(n416), .ZN(
        cell_1788_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1788_a_HPC2_and_U6 ( .A1(cell_1788_and_in[0]), .A2(n399), .ZN(
        cell_1788_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1788_a_HPC2_and_U5 ( .A(cell_1788_a_HPC2_and_n8), .B(
        cell_1788_a_HPC2_and_z_1__1_), .ZN(cell_1788_and_out[1]) );
  XNOR2_X1 cell_1788_a_HPC2_and_U4 ( .A(
        cell_1788_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1788_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1788_a_HPC2_and_n8) );
  XNOR2_X1 cell_1788_a_HPC2_and_U3 ( .A(cell_1788_a_HPC2_and_n7), .B(
        cell_1788_a_HPC2_and_z_0__0_), .ZN(cell_1788_and_out[0]) );
  XNOR2_X1 cell_1788_a_HPC2_and_U2 ( .A(
        cell_1788_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1788_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1788_a_HPC2_and_n7) );
  DFF_X1 cell_1788_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1788_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1788_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1788_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1788_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1788_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1788_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1788_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1788_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1788_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1789_U4 ( .A(n365), .B(cell_1789_and_out[1]), .Z(signal_3495)
         );
  XOR2_X1 cell_1789_U3 ( .A(n363), .B(cell_1789_and_out[0]), .Z(signal_2057)
         );
  XOR2_X1 cell_1789_U2 ( .A(n365), .B(signal_3426), .Z(cell_1789_and_in[1]) );
  XOR2_X1 cell_1789_U1 ( .A(n363), .B(signal_2012), .Z(cell_1789_and_in[0]) );
  XOR2_X1 cell_1789_a_HPC2_and_U14 ( .A(Fresh[75]), .B(cell_1789_and_in[0]), 
        .Z(cell_1789_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1789_a_HPC2_and_U13 ( .A(Fresh[75]), .B(cell_1789_and_in[1]), 
        .Z(cell_1789_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1789_a_HPC2_and_U12 ( .A1(cell_1789_a_HPC2_and_a_reg[1]), .A2(
        cell_1789_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1789_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1789_a_HPC2_and_U11 ( .A1(cell_1789_a_HPC2_and_a_reg[0]), .A2(
        cell_1789_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1789_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1789_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1789_a_HPC2_and_n9), 
        .ZN(cell_1789_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1789_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1789_a_HPC2_and_n9), 
        .ZN(cell_1789_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1789_a_HPC2_and_U8 ( .A(Fresh[75]), .ZN(cell_1789_a_HPC2_and_n9)
         );
  AND2_X1 cell_1789_a_HPC2_and_U7 ( .A1(cell_1789_and_in[1]), .A2(n416), .ZN(
        cell_1789_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1789_a_HPC2_and_U6 ( .A1(cell_1789_and_in[0]), .A2(n399), .ZN(
        cell_1789_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1789_a_HPC2_and_U5 ( .A(cell_1789_a_HPC2_and_n8), .B(
        cell_1789_a_HPC2_and_z_1__1_), .ZN(cell_1789_and_out[1]) );
  XNOR2_X1 cell_1789_a_HPC2_and_U4 ( .A(
        cell_1789_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1789_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1789_a_HPC2_and_n8) );
  XNOR2_X1 cell_1789_a_HPC2_and_U3 ( .A(cell_1789_a_HPC2_and_n7), .B(
        cell_1789_a_HPC2_and_z_0__0_), .ZN(cell_1789_and_out[0]) );
  XNOR2_X1 cell_1789_a_HPC2_and_U2 ( .A(
        cell_1789_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1789_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1789_a_HPC2_and_n7) );
  DFF_X1 cell_1789_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1789_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1789_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1789_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1789_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1789_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1789_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1789_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1789_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1789_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1790_U4 ( .A(n367), .B(cell_1790_and_out[1]), .Z(signal_3496)
         );
  XOR2_X1 cell_1790_U3 ( .A(n366), .B(cell_1790_and_out[0]), .Z(signal_2058)
         );
  XOR2_X1 cell_1790_U2 ( .A(n367), .B(n361), .Z(cell_1790_and_in[1]) );
  XOR2_X1 cell_1790_U1 ( .A(n366), .B(n359), .Z(cell_1790_and_in[0]) );
  XOR2_X1 cell_1790_a_HPC2_and_U14 ( .A(Fresh[76]), .B(cell_1790_and_in[0]), 
        .Z(cell_1790_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1790_a_HPC2_and_U13 ( .A(Fresh[76]), .B(cell_1790_and_in[1]), 
        .Z(cell_1790_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1790_a_HPC2_and_U12 ( .A1(cell_1790_a_HPC2_and_a_reg[1]), .A2(
        cell_1790_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1790_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1790_a_HPC2_and_U11 ( .A1(cell_1790_a_HPC2_and_a_reg[0]), .A2(
        cell_1790_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1790_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1790_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1790_a_HPC2_and_n9), 
        .ZN(cell_1790_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1790_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1790_a_HPC2_and_n9), 
        .ZN(cell_1790_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1790_a_HPC2_and_U8 ( .A(Fresh[76]), .ZN(cell_1790_a_HPC2_and_n9)
         );
  AND2_X1 cell_1790_a_HPC2_and_U7 ( .A1(cell_1790_and_in[1]), .A2(n416), .ZN(
        cell_1790_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1790_a_HPC2_and_U6 ( .A1(cell_1790_and_in[0]), .A2(n399), .ZN(
        cell_1790_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1790_a_HPC2_and_U5 ( .A(cell_1790_a_HPC2_and_n8), .B(
        cell_1790_a_HPC2_and_z_1__1_), .ZN(cell_1790_and_out[1]) );
  XNOR2_X1 cell_1790_a_HPC2_and_U4 ( .A(
        cell_1790_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1790_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1790_a_HPC2_and_n8) );
  XNOR2_X1 cell_1790_a_HPC2_and_U3 ( .A(cell_1790_a_HPC2_and_n7), .B(
        cell_1790_a_HPC2_and_z_0__0_), .ZN(cell_1790_and_out[0]) );
  XNOR2_X1 cell_1790_a_HPC2_and_U2 ( .A(
        cell_1790_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1790_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1790_a_HPC2_and_n7) );
  DFF_X1 cell_1790_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1790_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1790_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1790_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1790_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1790_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1790_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1790_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1790_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1790_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1791_U6 ( .A(cell_1791_n4), .B(cell_1791_and_out[1]), .Z(
        signal_3497) );
  XOR2_X1 cell_1791_U5 ( .A(cell_1791_n3), .B(cell_1791_and_out[0]), .Z(
        signal_2059) );
  XOR2_X1 cell_1791_U4 ( .A(cell_1791_n4), .B(signal_3406), .Z(
        cell_1791_and_in[1]) );
  XOR2_X1 cell_1791_U3 ( .A(cell_1791_n3), .B(signal_1992), .Z(
        cell_1791_and_in[0]) );
  BUF_X1 cell_1791_U2 ( .A(signal_3426), .Z(cell_1791_n4) );
  BUF_X1 cell_1791_U1 ( .A(signal_2012), .Z(cell_1791_n3) );
  XOR2_X1 cell_1791_a_HPC2_and_U14 ( .A(Fresh[77]), .B(cell_1791_and_in[0]), 
        .Z(cell_1791_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1791_a_HPC2_and_U13 ( .A(Fresh[77]), .B(cell_1791_and_in[1]), 
        .Z(cell_1791_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1791_a_HPC2_and_U12 ( .A1(cell_1791_a_HPC2_and_a_reg[1]), .A2(
        cell_1791_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1791_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1791_a_HPC2_and_U11 ( .A1(cell_1791_a_HPC2_and_a_reg[0]), .A2(
        cell_1791_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1791_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1791_a_HPC2_and_U10 ( .A1(n414), .A2(cell_1791_a_HPC2_and_n9), 
        .ZN(cell_1791_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1791_a_HPC2_and_U9 ( .A1(n397), .A2(cell_1791_a_HPC2_and_n9), 
        .ZN(cell_1791_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1791_a_HPC2_and_U8 ( .A(Fresh[77]), .ZN(cell_1791_a_HPC2_and_n9)
         );
  AND2_X1 cell_1791_a_HPC2_and_U7 ( .A1(cell_1791_and_in[1]), .A2(n414), .ZN(
        cell_1791_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1791_a_HPC2_and_U6 ( .A1(cell_1791_and_in[0]), .A2(n397), .ZN(
        cell_1791_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1791_a_HPC2_and_U5 ( .A(cell_1791_a_HPC2_and_n8), .B(
        cell_1791_a_HPC2_and_z_1__1_), .ZN(cell_1791_and_out[1]) );
  XNOR2_X1 cell_1791_a_HPC2_and_U4 ( .A(
        cell_1791_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1791_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1791_a_HPC2_and_n8) );
  XNOR2_X1 cell_1791_a_HPC2_and_U3 ( .A(cell_1791_a_HPC2_and_n7), .B(
        cell_1791_a_HPC2_and_z_0__0_), .ZN(cell_1791_and_out[0]) );
  XNOR2_X1 cell_1791_a_HPC2_and_U2 ( .A(
        cell_1791_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1791_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1791_a_HPC2_and_n7) );
  DFF_X1 cell_1791_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1791_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1791_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n397), .CK(clk), 
        .Q(cell_1791_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1791_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1791_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n414), .CK(clk), 
        .Q(cell_1791_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1791_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1791_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1791_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1792_U4 ( .A(n355), .B(cell_1792_and_out[1]), .Z(signal_3498)
         );
  XOR2_X1 cell_1792_U3 ( .A(n353), .B(cell_1792_and_out[0]), .Z(signal_2060)
         );
  XOR2_X1 cell_1792_U2 ( .A(n355), .B(n371), .Z(cell_1792_and_in[1]) );
  XOR2_X1 cell_1792_U1 ( .A(n353), .B(n369), .Z(cell_1792_and_in[0]) );
  XOR2_X1 cell_1792_a_HPC2_and_U14 ( .A(Fresh[78]), .B(cell_1792_and_in[0]), 
        .Z(cell_1792_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1792_a_HPC2_and_U13 ( .A(Fresh[78]), .B(cell_1792_and_in[1]), 
        .Z(cell_1792_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1792_a_HPC2_and_U12 ( .A1(cell_1792_a_HPC2_and_a_reg[1]), .A2(
        cell_1792_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1792_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1792_a_HPC2_and_U11 ( .A1(cell_1792_a_HPC2_and_a_reg[0]), .A2(
        cell_1792_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1792_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1792_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1792_a_HPC2_and_n9), 
        .ZN(cell_1792_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1792_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1792_a_HPC2_and_n9), 
        .ZN(cell_1792_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1792_a_HPC2_and_U8 ( .A(Fresh[78]), .ZN(cell_1792_a_HPC2_and_n9)
         );
  AND2_X1 cell_1792_a_HPC2_and_U7 ( .A1(cell_1792_and_in[1]), .A2(n416), .ZN(
        cell_1792_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1792_a_HPC2_and_U6 ( .A1(cell_1792_and_in[0]), .A2(n399), .ZN(
        cell_1792_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1792_a_HPC2_and_U5 ( .A(cell_1792_a_HPC2_and_n8), .B(
        cell_1792_a_HPC2_and_z_1__1_), .ZN(cell_1792_and_out[1]) );
  XNOR2_X1 cell_1792_a_HPC2_and_U4 ( .A(
        cell_1792_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1792_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1792_a_HPC2_and_n8) );
  XNOR2_X1 cell_1792_a_HPC2_and_U3 ( .A(cell_1792_a_HPC2_and_n7), .B(
        cell_1792_a_HPC2_and_z_0__0_), .ZN(cell_1792_and_out[0]) );
  XNOR2_X1 cell_1792_a_HPC2_and_U2 ( .A(
        cell_1792_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1792_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1792_a_HPC2_and_n7) );
  DFF_X1 cell_1792_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1792_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1792_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1792_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1792_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1792_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1792_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1792_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1792_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1792_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1793_U4 ( .A(n378), .B(cell_1793_and_out[1]), .Z(signal_3499)
         );
  XOR2_X1 cell_1793_U3 ( .A(n376), .B(cell_1793_and_out[0]), .Z(signal_2061)
         );
  XOR2_X1 cell_1793_U2 ( .A(n378), .B(signal_3261), .Z(cell_1793_and_in[1]) );
  XOR2_X1 cell_1793_U1 ( .A(n376), .B(signal_1987), .Z(cell_1793_and_in[0]) );
  XOR2_X1 cell_1793_a_HPC2_and_U14 ( .A(Fresh[79]), .B(cell_1793_and_in[0]), 
        .Z(cell_1793_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1793_a_HPC2_and_U13 ( .A(Fresh[79]), .B(cell_1793_and_in[1]), 
        .Z(cell_1793_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1793_a_HPC2_and_U12 ( .A1(cell_1793_a_HPC2_and_a_reg[1]), .A2(
        cell_1793_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1793_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1793_a_HPC2_and_U11 ( .A1(cell_1793_a_HPC2_and_a_reg[0]), .A2(
        cell_1793_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1793_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1793_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1793_a_HPC2_and_n9), 
        .ZN(cell_1793_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1793_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1793_a_HPC2_and_n9), 
        .ZN(cell_1793_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1793_a_HPC2_and_U8 ( .A(Fresh[79]), .ZN(cell_1793_a_HPC2_and_n9)
         );
  AND2_X1 cell_1793_a_HPC2_and_U7 ( .A1(cell_1793_and_in[1]), .A2(n416), .ZN(
        cell_1793_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1793_a_HPC2_and_U6 ( .A1(cell_1793_and_in[0]), .A2(n399), .ZN(
        cell_1793_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1793_a_HPC2_and_U5 ( .A(cell_1793_a_HPC2_and_n8), .B(
        cell_1793_a_HPC2_and_z_1__1_), .ZN(cell_1793_and_out[1]) );
  XNOR2_X1 cell_1793_a_HPC2_and_U4 ( .A(
        cell_1793_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1793_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1793_a_HPC2_and_n8) );
  XNOR2_X1 cell_1793_a_HPC2_and_U3 ( .A(cell_1793_a_HPC2_and_n7), .B(
        cell_1793_a_HPC2_and_z_0__0_), .ZN(cell_1793_and_out[0]) );
  XNOR2_X1 cell_1793_a_HPC2_and_U2 ( .A(
        cell_1793_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1793_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1793_a_HPC2_and_n7) );
  DFF_X1 cell_1793_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1793_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1793_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1793_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1793_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1793_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1793_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1793_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1793_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1793_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1794_U4 ( .A(signal_3406), .B(cell_1794_and_out[1]), .Z(
        signal_3500) );
  XOR2_X1 cell_1794_U3 ( .A(signal_1992), .B(cell_1794_and_out[0]), .Z(
        signal_2062) );
  XOR2_X1 cell_1794_U2 ( .A(signal_3406), .B(n375), .Z(cell_1794_and_in[1]) );
  XOR2_X1 cell_1794_U1 ( .A(signal_1992), .B(n373), .Z(cell_1794_and_in[0]) );
  XOR2_X1 cell_1794_a_HPC2_and_U14 ( .A(Fresh[80]), .B(cell_1794_and_in[0]), 
        .Z(cell_1794_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1794_a_HPC2_and_U13 ( .A(Fresh[80]), .B(cell_1794_and_in[1]), 
        .Z(cell_1794_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1794_a_HPC2_and_U12 ( .A1(cell_1794_a_HPC2_and_a_reg[1]), .A2(
        cell_1794_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1794_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1794_a_HPC2_and_U11 ( .A1(cell_1794_a_HPC2_and_a_reg[0]), .A2(
        cell_1794_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1794_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1794_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1794_a_HPC2_and_n9), 
        .ZN(cell_1794_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1794_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1794_a_HPC2_and_n9), 
        .ZN(cell_1794_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1794_a_HPC2_and_U8 ( .A(Fresh[80]), .ZN(cell_1794_a_HPC2_and_n9)
         );
  AND2_X1 cell_1794_a_HPC2_and_U7 ( .A1(cell_1794_and_in[1]), .A2(n419), .ZN(
        cell_1794_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1794_a_HPC2_and_U6 ( .A1(cell_1794_and_in[0]), .A2(n402), .ZN(
        cell_1794_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1794_a_HPC2_and_U5 ( .A(cell_1794_a_HPC2_and_n8), .B(
        cell_1794_a_HPC2_and_z_1__1_), .ZN(cell_1794_and_out[1]) );
  XNOR2_X1 cell_1794_a_HPC2_and_U4 ( .A(
        cell_1794_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1794_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1794_a_HPC2_and_n8) );
  XNOR2_X1 cell_1794_a_HPC2_and_U3 ( .A(cell_1794_a_HPC2_and_n7), .B(
        cell_1794_a_HPC2_and_z_0__0_), .ZN(cell_1794_and_out[0]) );
  XNOR2_X1 cell_1794_a_HPC2_and_U2 ( .A(
        cell_1794_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1794_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1794_a_HPC2_and_n7) );
  DFF_X1 cell_1794_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1794_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1794_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1794_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1794_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1794_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1794_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1794_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1794_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1794_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1795_U4 ( .A(signal_3427), .B(cell_1795_and_out[1]), .Z(
        signal_3501) );
  XOR2_X1 cell_1795_U3 ( .A(signal_2013), .B(cell_1795_and_out[0]), .Z(
        signal_2063) );
  XOR2_X1 cell_1795_U2 ( .A(signal_3427), .B(signal_3422), .Z(
        cell_1795_and_in[1]) );
  XOR2_X1 cell_1795_U1 ( .A(signal_2013), .B(signal_2008), .Z(
        cell_1795_and_in[0]) );
  XOR2_X1 cell_1795_a_HPC2_and_U14 ( .A(Fresh[81]), .B(cell_1795_and_in[0]), 
        .Z(cell_1795_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1795_a_HPC2_and_U13 ( .A(Fresh[81]), .B(cell_1795_and_in[1]), 
        .Z(cell_1795_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1795_a_HPC2_and_U12 ( .A1(cell_1795_a_HPC2_and_a_reg[1]), .A2(
        cell_1795_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1795_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1795_a_HPC2_and_U11 ( .A1(cell_1795_a_HPC2_and_a_reg[0]), .A2(
        cell_1795_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1795_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1795_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1795_a_HPC2_and_n9), 
        .ZN(cell_1795_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1795_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1795_a_HPC2_and_n9), 
        .ZN(cell_1795_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1795_a_HPC2_and_U8 ( .A(Fresh[81]), .ZN(cell_1795_a_HPC2_and_n9)
         );
  AND2_X1 cell_1795_a_HPC2_and_U7 ( .A1(cell_1795_and_in[1]), .A2(n442), .ZN(
        cell_1795_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1795_a_HPC2_and_U6 ( .A1(cell_1795_and_in[0]), .A2(n428), .ZN(
        cell_1795_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1795_a_HPC2_and_U5 ( .A(cell_1795_a_HPC2_and_n8), .B(
        cell_1795_a_HPC2_and_z_1__1_), .ZN(cell_1795_and_out[1]) );
  XNOR2_X1 cell_1795_a_HPC2_and_U4 ( .A(
        cell_1795_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1795_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1795_a_HPC2_and_n8) );
  XNOR2_X1 cell_1795_a_HPC2_and_U3 ( .A(cell_1795_a_HPC2_and_n7), .B(
        cell_1795_a_HPC2_and_z_0__0_), .ZN(cell_1795_and_out[0]) );
  XNOR2_X1 cell_1795_a_HPC2_and_U2 ( .A(
        cell_1795_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1795_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1795_a_HPC2_and_n7) );
  DFF_X1 cell_1795_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1795_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1795_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1795_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1795_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1795_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1795_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1795_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1795_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1795_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1796_U6 ( .A(cell_1796_n4), .B(cell_1796_and_out[1]), .Z(
        signal_3502) );
  XOR2_X1 cell_1796_U5 ( .A(cell_1796_n3), .B(cell_1796_and_out[0]), .Z(
        signal_2064) );
  XOR2_X1 cell_1796_U4 ( .A(cell_1796_n4), .B(n383), .Z(cell_1796_and_in[1])
         );
  XOR2_X1 cell_1796_U3 ( .A(cell_1796_n3), .B(n382), .Z(cell_1796_and_in[0])
         );
  BUF_X1 cell_1796_U2 ( .A(signal_3426), .Z(cell_1796_n4) );
  BUF_X1 cell_1796_U1 ( .A(signal_2012), .Z(cell_1796_n3) );
  XOR2_X1 cell_1796_a_HPC2_and_U14 ( .A(Fresh[82]), .B(cell_1796_and_in[0]), 
        .Z(cell_1796_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1796_a_HPC2_and_U13 ( .A(Fresh[82]), .B(cell_1796_and_in[1]), 
        .Z(cell_1796_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1796_a_HPC2_and_U12 ( .A1(cell_1796_a_HPC2_and_a_reg[1]), .A2(
        cell_1796_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1796_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1796_a_HPC2_and_U11 ( .A1(cell_1796_a_HPC2_and_a_reg[0]), .A2(
        cell_1796_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1796_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1796_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1796_a_HPC2_and_n9), 
        .ZN(cell_1796_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1796_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1796_a_HPC2_and_n9), 
        .ZN(cell_1796_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1796_a_HPC2_and_U8 ( .A(Fresh[82]), .ZN(cell_1796_a_HPC2_and_n9)
         );
  AND2_X1 cell_1796_a_HPC2_and_U7 ( .A1(cell_1796_and_in[1]), .A2(n420), .ZN(
        cell_1796_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1796_a_HPC2_and_U6 ( .A1(cell_1796_and_in[0]), .A2(n403), .ZN(
        cell_1796_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1796_a_HPC2_and_U5 ( .A(cell_1796_a_HPC2_and_n8), .B(
        cell_1796_a_HPC2_and_z_1__1_), .ZN(cell_1796_and_out[1]) );
  XNOR2_X1 cell_1796_a_HPC2_and_U4 ( .A(
        cell_1796_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1796_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1796_a_HPC2_and_n8) );
  XNOR2_X1 cell_1796_a_HPC2_and_U3 ( .A(cell_1796_a_HPC2_and_n7), .B(
        cell_1796_a_HPC2_and_z_0__0_), .ZN(cell_1796_and_out[0]) );
  XNOR2_X1 cell_1796_a_HPC2_and_U2 ( .A(
        cell_1796_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1796_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1796_a_HPC2_and_n7) );
  DFF_X1 cell_1796_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1796_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1796_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1796_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1796_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1796_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1796_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1796_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1796_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1796_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1797_U4 ( .A(n387), .B(cell_1797_and_out[1]), .Z(signal_3503)
         );
  XOR2_X1 cell_1797_U3 ( .A(n385), .B(cell_1797_and_out[0]), .Z(signal_2065)
         );
  XOR2_X1 cell_1797_U2 ( .A(n387), .B(n364), .Z(cell_1797_and_in[1]) );
  XOR2_X1 cell_1797_U1 ( .A(n385), .B(n362), .Z(cell_1797_and_in[0]) );
  XOR2_X1 cell_1797_a_HPC2_and_U14 ( .A(Fresh[83]), .B(cell_1797_and_in[0]), 
        .Z(cell_1797_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1797_a_HPC2_and_U13 ( .A(Fresh[83]), .B(cell_1797_and_in[1]), 
        .Z(cell_1797_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1797_a_HPC2_and_U12 ( .A1(cell_1797_a_HPC2_and_a_reg[1]), .A2(
        cell_1797_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1797_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1797_a_HPC2_and_U11 ( .A1(cell_1797_a_HPC2_and_a_reg[0]), .A2(
        cell_1797_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1797_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1797_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1797_a_HPC2_and_n9), 
        .ZN(cell_1797_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1797_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1797_a_HPC2_and_n9), 
        .ZN(cell_1797_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1797_a_HPC2_and_U8 ( .A(Fresh[83]), .ZN(cell_1797_a_HPC2_and_n9)
         );
  AND2_X1 cell_1797_a_HPC2_and_U7 ( .A1(cell_1797_and_in[1]), .A2(n416), .ZN(
        cell_1797_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1797_a_HPC2_and_U6 ( .A1(cell_1797_and_in[0]), .A2(n399), .ZN(
        cell_1797_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1797_a_HPC2_and_U5 ( .A(cell_1797_a_HPC2_and_n8), .B(
        cell_1797_a_HPC2_and_z_1__1_), .ZN(cell_1797_and_out[1]) );
  XNOR2_X1 cell_1797_a_HPC2_and_U4 ( .A(
        cell_1797_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1797_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1797_a_HPC2_and_n8) );
  XNOR2_X1 cell_1797_a_HPC2_and_U3 ( .A(cell_1797_a_HPC2_and_n7), .B(
        cell_1797_a_HPC2_and_z_0__0_), .ZN(cell_1797_and_out[0]) );
  XNOR2_X1 cell_1797_a_HPC2_and_U2 ( .A(
        cell_1797_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1797_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1797_a_HPC2_and_n7) );
  DFF_X1 cell_1797_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1797_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1797_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1797_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1797_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1797_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1797_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1797_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1797_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1797_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1798_U4 ( .A(n378), .B(cell_1798_and_out[1]), .Z(signal_3504)
         );
  XOR2_X1 cell_1798_U3 ( .A(n376), .B(cell_1798_and_out[0]), .Z(signal_2066)
         );
  XOR2_X1 cell_1798_U2 ( .A(n378), .B(n387), .Z(cell_1798_and_in[1]) );
  XOR2_X1 cell_1798_U1 ( .A(n376), .B(n385), .Z(cell_1798_and_in[0]) );
  XOR2_X1 cell_1798_a_HPC2_and_U14 ( .A(Fresh[84]), .B(cell_1798_and_in[0]), 
        .Z(cell_1798_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1798_a_HPC2_and_U13 ( .A(Fresh[84]), .B(cell_1798_and_in[1]), 
        .Z(cell_1798_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1798_a_HPC2_and_U12 ( .A1(cell_1798_a_HPC2_and_a_reg[1]), .A2(
        cell_1798_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1798_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1798_a_HPC2_and_U11 ( .A1(cell_1798_a_HPC2_and_a_reg[0]), .A2(
        cell_1798_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1798_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1798_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1798_a_HPC2_and_n9), 
        .ZN(cell_1798_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1798_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1798_a_HPC2_and_n9), 
        .ZN(cell_1798_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1798_a_HPC2_and_U8 ( .A(Fresh[84]), .ZN(cell_1798_a_HPC2_and_n9)
         );
  AND2_X1 cell_1798_a_HPC2_and_U7 ( .A1(cell_1798_and_in[1]), .A2(n417), .ZN(
        cell_1798_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1798_a_HPC2_and_U6 ( .A1(cell_1798_and_in[0]), .A2(n400), .ZN(
        cell_1798_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1798_a_HPC2_and_U5 ( .A(cell_1798_a_HPC2_and_n8), .B(
        cell_1798_a_HPC2_and_z_1__1_), .ZN(cell_1798_and_out[1]) );
  XNOR2_X1 cell_1798_a_HPC2_and_U4 ( .A(
        cell_1798_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1798_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1798_a_HPC2_and_n8) );
  XNOR2_X1 cell_1798_a_HPC2_and_U3 ( .A(cell_1798_a_HPC2_and_n7), .B(
        cell_1798_a_HPC2_and_z_0__0_), .ZN(cell_1798_and_out[0]) );
  XNOR2_X1 cell_1798_a_HPC2_and_U2 ( .A(
        cell_1798_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1798_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1798_a_HPC2_and_n7) );
  DFF_X1 cell_1798_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1798_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1798_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1798_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1798_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1798_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1798_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1798_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1798_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1798_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1799_U4 ( .A(n386), .B(cell_1799_and_out[1]), .Z(signal_3505)
         );
  XOR2_X1 cell_1799_U3 ( .A(n384), .B(cell_1799_and_out[0]), .Z(signal_2067)
         );
  XOR2_X1 cell_1799_U2 ( .A(n386), .B(signal_3413), .Z(cell_1799_and_in[1]) );
  XOR2_X1 cell_1799_U1 ( .A(n384), .B(signal_1999), .Z(cell_1799_and_in[0]) );
  XOR2_X1 cell_1799_a_HPC2_and_U14 ( .A(Fresh[85]), .B(cell_1799_and_in[0]), 
        .Z(cell_1799_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1799_a_HPC2_and_U13 ( .A(Fresh[85]), .B(cell_1799_and_in[1]), 
        .Z(cell_1799_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1799_a_HPC2_and_U12 ( .A1(cell_1799_a_HPC2_and_a_reg[1]), .A2(
        cell_1799_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1799_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1799_a_HPC2_and_U11 ( .A1(cell_1799_a_HPC2_and_a_reg[0]), .A2(
        cell_1799_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1799_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1799_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1799_a_HPC2_and_n9), 
        .ZN(cell_1799_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1799_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1799_a_HPC2_and_n9), 
        .ZN(cell_1799_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1799_a_HPC2_and_U8 ( .A(Fresh[85]), .ZN(cell_1799_a_HPC2_and_n9)
         );
  AND2_X1 cell_1799_a_HPC2_and_U7 ( .A1(cell_1799_and_in[1]), .A2(n417), .ZN(
        cell_1799_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1799_a_HPC2_and_U6 ( .A1(cell_1799_and_in[0]), .A2(n400), .ZN(
        cell_1799_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1799_a_HPC2_and_U5 ( .A(cell_1799_a_HPC2_and_n8), .B(
        cell_1799_a_HPC2_and_z_1__1_), .ZN(cell_1799_and_out[1]) );
  XNOR2_X1 cell_1799_a_HPC2_and_U4 ( .A(
        cell_1799_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1799_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1799_a_HPC2_and_n8) );
  XNOR2_X1 cell_1799_a_HPC2_and_U3 ( .A(cell_1799_a_HPC2_and_n7), .B(
        cell_1799_a_HPC2_and_z_0__0_), .ZN(cell_1799_and_out[0]) );
  XNOR2_X1 cell_1799_a_HPC2_and_U2 ( .A(
        cell_1799_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1799_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1799_a_HPC2_and_n7) );
  DFF_X1 cell_1799_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1799_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1799_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1799_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1799_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1799_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1799_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1799_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1799_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1799_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1800_U4 ( .A(1'b0), .B(cell_1800_and_out[1]), .Z(signal_3506)
         );
  XOR2_X1 cell_1800_U3 ( .A(1'b1), .B(cell_1800_and_out[0]), .Z(signal_2068)
         );
  XOR2_X1 cell_1800_U2 ( .A(1'b0), .B(signal_3407), .Z(cell_1800_and_in[1]) );
  XOR2_X1 cell_1800_U1 ( .A(1'b1), .B(signal_1993), .Z(cell_1800_and_in[0]) );
  XOR2_X1 cell_1800_a_HPC2_and_U14 ( .A(Fresh[86]), .B(cell_1800_and_in[0]), 
        .Z(cell_1800_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1800_a_HPC2_and_U13 ( .A(Fresh[86]), .B(cell_1800_and_in[1]), 
        .Z(cell_1800_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1800_a_HPC2_and_U12 ( .A1(cell_1800_a_HPC2_and_a_reg[1]), .A2(
        cell_1800_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1800_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1800_a_HPC2_and_U11 ( .A1(cell_1800_a_HPC2_and_a_reg[0]), .A2(
        cell_1800_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1800_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1800_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1800_a_HPC2_and_n9), 
        .ZN(cell_1800_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1800_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1800_a_HPC2_and_n9), 
        .ZN(cell_1800_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1800_a_HPC2_and_U8 ( .A(Fresh[86]), .ZN(cell_1800_a_HPC2_and_n9)
         );
  AND2_X1 cell_1800_a_HPC2_and_U7 ( .A1(cell_1800_and_in[1]), .A2(n422), .ZN(
        cell_1800_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1800_a_HPC2_and_U6 ( .A1(cell_1800_and_in[0]), .A2(n398), .ZN(
        cell_1800_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1800_a_HPC2_and_U5 ( .A(cell_1800_a_HPC2_and_n8), .B(
        cell_1800_a_HPC2_and_z_1__1_), .ZN(cell_1800_and_out[1]) );
  XNOR2_X1 cell_1800_a_HPC2_and_U4 ( .A(
        cell_1800_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1800_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1800_a_HPC2_and_n8) );
  XNOR2_X1 cell_1800_a_HPC2_and_U3 ( .A(cell_1800_a_HPC2_and_n7), .B(
        cell_1800_a_HPC2_and_z_0__0_), .ZN(cell_1800_and_out[0]) );
  XNOR2_X1 cell_1800_a_HPC2_and_U2 ( .A(
        cell_1800_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1800_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1800_a_HPC2_and_n7) );
  DFF_X1 cell_1800_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1800_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1800_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1800_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1800_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1800_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1800_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1800_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1800_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1800_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1801_U4 ( .A(n367), .B(cell_1801_and_out[1]), .Z(signal_3507)
         );
  XOR2_X1 cell_1801_U3 ( .A(n366), .B(cell_1801_and_out[0]), .Z(signal_2069)
         );
  XOR2_X1 cell_1801_U2 ( .A(n367), .B(n357), .Z(cell_1801_and_in[1]) );
  XOR2_X1 cell_1801_U1 ( .A(n366), .B(n356), .Z(cell_1801_and_in[0]) );
  XOR2_X1 cell_1801_a_HPC2_and_U14 ( .A(Fresh[87]), .B(cell_1801_and_in[0]), 
        .Z(cell_1801_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1801_a_HPC2_and_U13 ( .A(Fresh[87]), .B(cell_1801_and_in[1]), 
        .Z(cell_1801_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1801_a_HPC2_and_U12 ( .A1(cell_1801_a_HPC2_and_a_reg[1]), .A2(
        cell_1801_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1801_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1801_a_HPC2_and_U11 ( .A1(cell_1801_a_HPC2_and_a_reg[0]), .A2(
        cell_1801_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1801_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1801_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1801_a_HPC2_and_n9), 
        .ZN(cell_1801_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1801_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1801_a_HPC2_and_n9), 
        .ZN(cell_1801_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1801_a_HPC2_and_U8 ( .A(Fresh[87]), .ZN(cell_1801_a_HPC2_and_n9)
         );
  AND2_X1 cell_1801_a_HPC2_and_U7 ( .A1(cell_1801_and_in[1]), .A2(n417), .ZN(
        cell_1801_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1801_a_HPC2_and_U6 ( .A1(cell_1801_and_in[0]), .A2(n400), .ZN(
        cell_1801_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1801_a_HPC2_and_U5 ( .A(cell_1801_a_HPC2_and_n8), .B(
        cell_1801_a_HPC2_and_z_1__1_), .ZN(cell_1801_and_out[1]) );
  XNOR2_X1 cell_1801_a_HPC2_and_U4 ( .A(
        cell_1801_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1801_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1801_a_HPC2_and_n8) );
  XNOR2_X1 cell_1801_a_HPC2_and_U3 ( .A(cell_1801_a_HPC2_and_n7), .B(
        cell_1801_a_HPC2_and_z_0__0_), .ZN(cell_1801_and_out[0]) );
  XNOR2_X1 cell_1801_a_HPC2_and_U2 ( .A(
        cell_1801_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1801_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1801_a_HPC2_and_n7) );
  DFF_X1 cell_1801_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1801_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1801_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1801_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1801_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1801_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1801_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1801_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1801_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1801_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1802_U4 ( .A(n367), .B(cell_1802_and_out[1]), .Z(signal_3508)
         );
  XOR2_X1 cell_1802_U3 ( .A(n366), .B(cell_1802_and_out[0]), .Z(signal_2070)
         );
  XOR2_X1 cell_1802_U2 ( .A(n367), .B(signal_3258), .Z(cell_1802_and_in[1]) );
  XOR2_X1 cell_1802_U1 ( .A(n366), .B(signal_1984), .Z(cell_1802_and_in[0]) );
  XOR2_X1 cell_1802_a_HPC2_and_U14 ( .A(Fresh[88]), .B(cell_1802_and_in[0]), 
        .Z(cell_1802_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1802_a_HPC2_and_U13 ( .A(Fresh[88]), .B(cell_1802_and_in[1]), 
        .Z(cell_1802_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1802_a_HPC2_and_U12 ( .A1(cell_1802_a_HPC2_and_a_reg[1]), .A2(
        cell_1802_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1802_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1802_a_HPC2_and_U11 ( .A1(cell_1802_a_HPC2_and_a_reg[0]), .A2(
        cell_1802_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1802_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1802_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1802_a_HPC2_and_n9), 
        .ZN(cell_1802_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1802_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1802_a_HPC2_and_n9), 
        .ZN(cell_1802_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1802_a_HPC2_and_U8 ( .A(Fresh[88]), .ZN(cell_1802_a_HPC2_and_n9)
         );
  AND2_X1 cell_1802_a_HPC2_and_U7 ( .A1(cell_1802_and_in[1]), .A2(n417), .ZN(
        cell_1802_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1802_a_HPC2_and_U6 ( .A1(cell_1802_and_in[0]), .A2(n400), .ZN(
        cell_1802_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1802_a_HPC2_and_U5 ( .A(cell_1802_a_HPC2_and_n8), .B(
        cell_1802_a_HPC2_and_z_1__1_), .ZN(cell_1802_and_out[1]) );
  XNOR2_X1 cell_1802_a_HPC2_and_U4 ( .A(
        cell_1802_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1802_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1802_a_HPC2_and_n8) );
  XNOR2_X1 cell_1802_a_HPC2_and_U3 ( .A(cell_1802_a_HPC2_and_n7), .B(
        cell_1802_a_HPC2_and_z_0__0_), .ZN(cell_1802_and_out[0]) );
  XNOR2_X1 cell_1802_a_HPC2_and_U2 ( .A(
        cell_1802_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1802_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1802_a_HPC2_and_n7) );
  DFF_X1 cell_1802_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1802_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1802_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1802_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1802_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1802_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1802_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1802_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1802_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1802_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1803_U4 ( .A(signal_3406), .B(cell_1803_and_out[1]), .Z(
        signal_3509) );
  XOR2_X1 cell_1803_U3 ( .A(signal_1992), .B(cell_1803_and_out[0]), .Z(
        signal_2071) );
  XOR2_X1 cell_1803_U2 ( .A(signal_3406), .B(n371), .Z(cell_1803_and_in[1]) );
  XOR2_X1 cell_1803_U1 ( .A(signal_1992), .B(n369), .Z(cell_1803_and_in[0]) );
  XOR2_X1 cell_1803_a_HPC2_and_U14 ( .A(Fresh[89]), .B(cell_1803_and_in[0]), 
        .Z(cell_1803_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1803_a_HPC2_and_U13 ( .A(Fresh[89]), .B(cell_1803_and_in[1]), 
        .Z(cell_1803_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1803_a_HPC2_and_U12 ( .A1(cell_1803_a_HPC2_and_a_reg[1]), .A2(
        cell_1803_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1803_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1803_a_HPC2_and_U11 ( .A1(cell_1803_a_HPC2_and_a_reg[0]), .A2(
        cell_1803_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1803_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1803_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1803_a_HPC2_and_n9), 
        .ZN(cell_1803_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1803_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1803_a_HPC2_and_n9), 
        .ZN(cell_1803_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1803_a_HPC2_and_U8 ( .A(Fresh[89]), .ZN(cell_1803_a_HPC2_and_n9)
         );
  AND2_X1 cell_1803_a_HPC2_and_U7 ( .A1(cell_1803_and_in[1]), .A2(n418), .ZN(
        cell_1803_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1803_a_HPC2_and_U6 ( .A1(cell_1803_and_in[0]), .A2(n401), .ZN(
        cell_1803_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1803_a_HPC2_and_U5 ( .A(cell_1803_a_HPC2_and_n8), .B(
        cell_1803_a_HPC2_and_z_1__1_), .ZN(cell_1803_and_out[1]) );
  XNOR2_X1 cell_1803_a_HPC2_and_U4 ( .A(
        cell_1803_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1803_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1803_a_HPC2_and_n8) );
  XNOR2_X1 cell_1803_a_HPC2_and_U3 ( .A(cell_1803_a_HPC2_and_n7), .B(
        cell_1803_a_HPC2_and_z_0__0_), .ZN(cell_1803_and_out[0]) );
  XNOR2_X1 cell_1803_a_HPC2_and_U2 ( .A(
        cell_1803_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1803_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1803_a_HPC2_and_n7) );
  DFF_X1 cell_1803_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1803_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1803_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1803_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1803_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1803_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1803_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1803_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1803_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1803_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1804_U4 ( .A(n381), .B(cell_1804_and_out[1]), .Z(signal_3510)
         );
  XOR2_X1 cell_1804_U3 ( .A(n380), .B(cell_1804_and_out[0]), .Z(signal_2072)
         );
  XOR2_X1 cell_1804_U2 ( .A(n381), .B(n367), .Z(cell_1804_and_in[1]) );
  XOR2_X1 cell_1804_U1 ( .A(n380), .B(n366), .Z(cell_1804_and_in[0]) );
  XOR2_X1 cell_1804_a_HPC2_and_U14 ( .A(Fresh[90]), .B(cell_1804_and_in[0]), 
        .Z(cell_1804_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1804_a_HPC2_and_U13 ( .A(Fresh[90]), .B(cell_1804_and_in[1]), 
        .Z(cell_1804_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1804_a_HPC2_and_U12 ( .A1(cell_1804_a_HPC2_and_a_reg[1]), .A2(
        cell_1804_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1804_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1804_a_HPC2_and_U11 ( .A1(cell_1804_a_HPC2_and_a_reg[0]), .A2(
        cell_1804_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1804_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1804_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1804_a_HPC2_and_n9), 
        .ZN(cell_1804_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1804_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1804_a_HPC2_and_n9), 
        .ZN(cell_1804_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1804_a_HPC2_and_U8 ( .A(Fresh[90]), .ZN(cell_1804_a_HPC2_and_n9)
         );
  AND2_X1 cell_1804_a_HPC2_and_U7 ( .A1(cell_1804_and_in[1]), .A2(n417), .ZN(
        cell_1804_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1804_a_HPC2_and_U6 ( .A1(cell_1804_and_in[0]), .A2(n400), .ZN(
        cell_1804_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1804_a_HPC2_and_U5 ( .A(cell_1804_a_HPC2_and_n8), .B(
        cell_1804_a_HPC2_and_z_1__1_), .ZN(cell_1804_and_out[1]) );
  XNOR2_X1 cell_1804_a_HPC2_and_U4 ( .A(
        cell_1804_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1804_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1804_a_HPC2_and_n8) );
  XNOR2_X1 cell_1804_a_HPC2_and_U3 ( .A(cell_1804_a_HPC2_and_n7), .B(
        cell_1804_a_HPC2_and_z_0__0_), .ZN(cell_1804_and_out[0]) );
  XNOR2_X1 cell_1804_a_HPC2_and_U2 ( .A(
        cell_1804_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1804_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1804_a_HPC2_and_n7) );
  DFF_X1 cell_1804_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1804_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1804_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1804_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1804_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1804_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1804_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1804_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1804_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1804_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1805_U4 ( .A(signal_3427), .B(cell_1805_and_out[1]), .Z(
        signal_3511) );
  XOR2_X1 cell_1805_U3 ( .A(signal_2013), .B(cell_1805_and_out[0]), .Z(
        signal_2073) );
  XOR2_X1 cell_1805_U2 ( .A(signal_3427), .B(signal_3256), .Z(
        cell_1805_and_in[1]) );
  XOR2_X1 cell_1805_U1 ( .A(signal_2013), .B(signal_1982), .Z(
        cell_1805_and_in[0]) );
  XOR2_X1 cell_1805_a_HPC2_and_U14 ( .A(Fresh[91]), .B(cell_1805_and_in[0]), 
        .Z(cell_1805_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1805_a_HPC2_and_U13 ( .A(Fresh[91]), .B(cell_1805_and_in[1]), 
        .Z(cell_1805_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1805_a_HPC2_and_U12 ( .A1(cell_1805_a_HPC2_and_a_reg[1]), .A2(
        cell_1805_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1805_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1805_a_HPC2_and_U11 ( .A1(cell_1805_a_HPC2_and_a_reg[0]), .A2(
        cell_1805_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1805_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1805_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1805_a_HPC2_and_n9), 
        .ZN(cell_1805_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1805_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1805_a_HPC2_and_n9), 
        .ZN(cell_1805_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1805_a_HPC2_and_U8 ( .A(Fresh[91]), .ZN(cell_1805_a_HPC2_and_n9)
         );
  AND2_X1 cell_1805_a_HPC2_and_U7 ( .A1(cell_1805_and_in[1]), .A2(n417), .ZN(
        cell_1805_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1805_a_HPC2_and_U6 ( .A1(cell_1805_and_in[0]), .A2(n400), .ZN(
        cell_1805_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1805_a_HPC2_and_U5 ( .A(cell_1805_a_HPC2_and_n8), .B(
        cell_1805_a_HPC2_and_z_1__1_), .ZN(cell_1805_and_out[1]) );
  XNOR2_X1 cell_1805_a_HPC2_and_U4 ( .A(
        cell_1805_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1805_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1805_a_HPC2_and_n8) );
  XNOR2_X1 cell_1805_a_HPC2_and_U3 ( .A(cell_1805_a_HPC2_and_n7), .B(
        cell_1805_a_HPC2_and_z_0__0_), .ZN(cell_1805_and_out[0]) );
  XNOR2_X1 cell_1805_a_HPC2_and_U2 ( .A(
        cell_1805_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1805_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1805_a_HPC2_and_n7) );
  DFF_X1 cell_1805_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1805_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1805_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1805_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1805_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1805_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1805_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1805_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1805_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1805_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1806_U4 ( .A(n378), .B(cell_1806_and_out[1]), .Z(signal_3512)
         );
  XOR2_X1 cell_1806_U3 ( .A(n376), .B(cell_1806_and_out[0]), .Z(signal_2074)
         );
  XOR2_X1 cell_1806_U2 ( .A(n378), .B(n371), .Z(cell_1806_and_in[1]) );
  XOR2_X1 cell_1806_U1 ( .A(n376), .B(n369), .Z(cell_1806_and_in[0]) );
  XOR2_X1 cell_1806_a_HPC2_and_U14 ( .A(Fresh[92]), .B(cell_1806_and_in[0]), 
        .Z(cell_1806_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1806_a_HPC2_and_U13 ( .A(Fresh[92]), .B(cell_1806_and_in[1]), 
        .Z(cell_1806_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1806_a_HPC2_and_U12 ( .A1(cell_1806_a_HPC2_and_a_reg[1]), .A2(
        cell_1806_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1806_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1806_a_HPC2_and_U11 ( .A1(cell_1806_a_HPC2_and_a_reg[0]), .A2(
        cell_1806_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1806_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1806_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1806_a_HPC2_and_n9), 
        .ZN(cell_1806_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1806_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1806_a_HPC2_and_n9), 
        .ZN(cell_1806_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1806_a_HPC2_and_U8 ( .A(Fresh[92]), .ZN(cell_1806_a_HPC2_and_n9)
         );
  AND2_X1 cell_1806_a_HPC2_and_U7 ( .A1(cell_1806_and_in[1]), .A2(n417), .ZN(
        cell_1806_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1806_a_HPC2_and_U6 ( .A1(cell_1806_and_in[0]), .A2(n400), .ZN(
        cell_1806_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1806_a_HPC2_and_U5 ( .A(cell_1806_a_HPC2_and_n8), .B(
        cell_1806_a_HPC2_and_z_1__1_), .ZN(cell_1806_and_out[1]) );
  XNOR2_X1 cell_1806_a_HPC2_and_U4 ( .A(
        cell_1806_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1806_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1806_a_HPC2_and_n8) );
  XNOR2_X1 cell_1806_a_HPC2_and_U3 ( .A(cell_1806_a_HPC2_and_n7), .B(
        cell_1806_a_HPC2_and_z_0__0_), .ZN(cell_1806_and_out[0]) );
  XNOR2_X1 cell_1806_a_HPC2_and_U2 ( .A(
        cell_1806_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1806_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1806_a_HPC2_and_n7) );
  DFF_X1 cell_1806_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1806_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1806_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1806_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1806_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1806_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1806_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1806_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1806_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1806_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1807_U6 ( .A(cell_1807_n4), .B(cell_1807_and_out[1]), .Z(
        signal_3513) );
  XOR2_X1 cell_1807_U5 ( .A(cell_1807_n3), .B(cell_1807_and_out[0]), .Z(
        signal_2075) );
  XOR2_X1 cell_1807_U4 ( .A(cell_1807_n4), .B(n357), .Z(cell_1807_and_in[1])
         );
  XOR2_X1 cell_1807_U3 ( .A(cell_1807_n3), .B(n356), .Z(cell_1807_and_in[0])
         );
  BUF_X1 cell_1807_U2 ( .A(signal_3426), .Z(cell_1807_n4) );
  BUF_X1 cell_1807_U1 ( .A(signal_2012), .Z(cell_1807_n3) );
  XOR2_X1 cell_1807_a_HPC2_and_U14 ( .A(Fresh[93]), .B(cell_1807_and_in[0]), 
        .Z(cell_1807_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1807_a_HPC2_and_U13 ( .A(Fresh[93]), .B(cell_1807_and_in[1]), 
        .Z(cell_1807_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1807_a_HPC2_and_U12 ( .A1(cell_1807_a_HPC2_and_a_reg[1]), .A2(
        cell_1807_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1807_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1807_a_HPC2_and_U11 ( .A1(cell_1807_a_HPC2_and_a_reg[0]), .A2(
        cell_1807_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1807_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1807_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1807_a_HPC2_and_n9), 
        .ZN(cell_1807_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1807_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1807_a_HPC2_and_n9), 
        .ZN(cell_1807_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1807_a_HPC2_and_U8 ( .A(Fresh[93]), .ZN(cell_1807_a_HPC2_and_n9)
         );
  AND2_X1 cell_1807_a_HPC2_and_U7 ( .A1(cell_1807_and_in[1]), .A2(n421), .ZN(
        cell_1807_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1807_a_HPC2_and_U6 ( .A1(cell_1807_and_in[0]), .A2(n404), .ZN(
        cell_1807_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1807_a_HPC2_and_U5 ( .A(cell_1807_a_HPC2_and_n8), .B(
        cell_1807_a_HPC2_and_z_1__1_), .ZN(cell_1807_and_out[1]) );
  XNOR2_X1 cell_1807_a_HPC2_and_U4 ( .A(
        cell_1807_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1807_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1807_a_HPC2_and_n8) );
  XNOR2_X1 cell_1807_a_HPC2_and_U3 ( .A(cell_1807_a_HPC2_and_n7), .B(
        cell_1807_a_HPC2_and_z_0__0_), .ZN(cell_1807_and_out[0]) );
  XNOR2_X1 cell_1807_a_HPC2_and_U2 ( .A(
        cell_1807_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1807_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1807_a_HPC2_and_n7) );
  DFF_X1 cell_1807_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1807_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1807_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1807_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1807_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1807_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1807_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1807_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1807_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1807_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1808_U4 ( .A(n383), .B(cell_1808_and_out[1]), .Z(signal_3514)
         );
  XOR2_X1 cell_1808_U3 ( .A(n382), .B(cell_1808_and_out[0]), .Z(signal_2076)
         );
  XOR2_X1 cell_1808_U2 ( .A(n383), .B(n367), .Z(cell_1808_and_in[1]) );
  XOR2_X1 cell_1808_U1 ( .A(n382), .B(n366), .Z(cell_1808_and_in[0]) );
  XOR2_X1 cell_1808_a_HPC2_and_U14 ( .A(Fresh[94]), .B(cell_1808_and_in[0]), 
        .Z(cell_1808_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1808_a_HPC2_and_U13 ( .A(Fresh[94]), .B(cell_1808_and_in[1]), 
        .Z(cell_1808_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1808_a_HPC2_and_U12 ( .A1(cell_1808_a_HPC2_and_a_reg[1]), .A2(
        cell_1808_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1808_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1808_a_HPC2_and_U11 ( .A1(cell_1808_a_HPC2_and_a_reg[0]), .A2(
        cell_1808_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1808_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1808_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1808_a_HPC2_and_n9), 
        .ZN(cell_1808_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1808_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1808_a_HPC2_and_n9), 
        .ZN(cell_1808_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1808_a_HPC2_and_U8 ( .A(Fresh[94]), .ZN(cell_1808_a_HPC2_and_n9)
         );
  AND2_X1 cell_1808_a_HPC2_and_U7 ( .A1(cell_1808_and_in[1]), .A2(n418), .ZN(
        cell_1808_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1808_a_HPC2_and_U6 ( .A1(cell_1808_and_in[0]), .A2(n401), .ZN(
        cell_1808_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1808_a_HPC2_and_U5 ( .A(cell_1808_a_HPC2_and_n8), .B(
        cell_1808_a_HPC2_and_z_1__1_), .ZN(cell_1808_and_out[1]) );
  XNOR2_X1 cell_1808_a_HPC2_and_U4 ( .A(
        cell_1808_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1808_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1808_a_HPC2_and_n8) );
  XNOR2_X1 cell_1808_a_HPC2_and_U3 ( .A(cell_1808_a_HPC2_and_n7), .B(
        cell_1808_a_HPC2_and_z_0__0_), .ZN(cell_1808_and_out[0]) );
  XNOR2_X1 cell_1808_a_HPC2_and_U2 ( .A(
        cell_1808_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1808_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1808_a_HPC2_and_n7) );
  DFF_X1 cell_1808_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1808_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1808_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1808_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1808_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1808_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1808_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1808_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1808_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1808_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1809_U4 ( .A(1'b0), .B(cell_1809_and_out[1]), .Z(signal_3515)
         );
  XOR2_X1 cell_1809_U3 ( .A(1'b1), .B(cell_1809_and_out[0]), .Z(signal_2077)
         );
  XOR2_X1 cell_1809_U2 ( .A(1'b0), .B(n355), .Z(cell_1809_and_in[1]) );
  XOR2_X1 cell_1809_U1 ( .A(1'b1), .B(n353), .Z(cell_1809_and_in[0]) );
  XOR2_X1 cell_1809_a_HPC2_and_U14 ( .A(Fresh[95]), .B(cell_1809_and_in[0]), 
        .Z(cell_1809_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1809_a_HPC2_and_U13 ( .A(Fresh[95]), .B(cell_1809_and_in[1]), 
        .Z(cell_1809_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1809_a_HPC2_and_U12 ( .A1(cell_1809_a_HPC2_and_a_reg[1]), .A2(
        cell_1809_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1809_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1809_a_HPC2_and_U11 ( .A1(cell_1809_a_HPC2_and_a_reg[0]), .A2(
        cell_1809_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1809_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1809_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1809_a_HPC2_and_n9), 
        .ZN(cell_1809_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1809_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1809_a_HPC2_and_n9), 
        .ZN(cell_1809_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1809_a_HPC2_and_U8 ( .A(Fresh[95]), .ZN(cell_1809_a_HPC2_and_n9)
         );
  AND2_X1 cell_1809_a_HPC2_and_U7 ( .A1(cell_1809_and_in[1]), .A2(n415), .ZN(
        cell_1809_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1809_a_HPC2_and_U6 ( .A1(cell_1809_and_in[0]), .A2(n405), .ZN(
        cell_1809_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1809_a_HPC2_and_U5 ( .A(cell_1809_a_HPC2_and_n8), .B(
        cell_1809_a_HPC2_and_z_1__1_), .ZN(cell_1809_and_out[1]) );
  XNOR2_X1 cell_1809_a_HPC2_and_U4 ( .A(
        cell_1809_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1809_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1809_a_HPC2_and_n8) );
  XNOR2_X1 cell_1809_a_HPC2_and_U3 ( .A(cell_1809_a_HPC2_and_n7), .B(
        cell_1809_a_HPC2_and_z_0__0_), .ZN(cell_1809_and_out[0]) );
  XNOR2_X1 cell_1809_a_HPC2_and_U2 ( .A(
        cell_1809_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1809_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1809_a_HPC2_and_n7) );
  DFF_X1 cell_1809_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1809_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1809_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1809_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1809_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1809_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1809_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1809_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1809_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1809_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1810_U4 ( .A(n367), .B(cell_1810_and_out[1]), .Z(signal_3516)
         );
  XOR2_X1 cell_1810_U3 ( .A(n366), .B(cell_1810_and_out[0]), .Z(signal_2078)
         );
  XOR2_X1 cell_1810_U2 ( .A(n367), .B(n387), .Z(cell_1810_and_in[1]) );
  XOR2_X1 cell_1810_U1 ( .A(n366), .B(n385), .Z(cell_1810_and_in[0]) );
  XOR2_X1 cell_1810_a_HPC2_and_U14 ( .A(Fresh[96]), .B(cell_1810_and_in[0]), 
        .Z(cell_1810_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1810_a_HPC2_and_U13 ( .A(Fresh[96]), .B(cell_1810_and_in[1]), 
        .Z(cell_1810_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1810_a_HPC2_and_U12 ( .A1(cell_1810_a_HPC2_and_a_reg[1]), .A2(
        cell_1810_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1810_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1810_a_HPC2_and_U11 ( .A1(cell_1810_a_HPC2_and_a_reg[0]), .A2(
        cell_1810_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1810_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1810_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1810_a_HPC2_and_n9), 
        .ZN(cell_1810_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1810_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1810_a_HPC2_and_n9), 
        .ZN(cell_1810_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1810_a_HPC2_and_U8 ( .A(Fresh[96]), .ZN(cell_1810_a_HPC2_and_n9)
         );
  AND2_X1 cell_1810_a_HPC2_and_U7 ( .A1(cell_1810_and_in[1]), .A2(n418), .ZN(
        cell_1810_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1810_a_HPC2_and_U6 ( .A1(cell_1810_and_in[0]), .A2(n401), .ZN(
        cell_1810_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1810_a_HPC2_and_U5 ( .A(cell_1810_a_HPC2_and_n8), .B(
        cell_1810_a_HPC2_and_z_1__1_), .ZN(cell_1810_and_out[1]) );
  XNOR2_X1 cell_1810_a_HPC2_and_U4 ( .A(
        cell_1810_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1810_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1810_a_HPC2_and_n8) );
  XNOR2_X1 cell_1810_a_HPC2_and_U3 ( .A(cell_1810_a_HPC2_and_n7), .B(
        cell_1810_a_HPC2_and_z_0__0_), .ZN(cell_1810_and_out[0]) );
  XNOR2_X1 cell_1810_a_HPC2_and_U2 ( .A(
        cell_1810_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1810_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1810_a_HPC2_and_n7) );
  DFF_X1 cell_1810_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1810_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1810_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1810_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1810_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1810_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1810_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1810_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1810_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1810_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1811_U4 ( .A(n378), .B(cell_1811_and_out[1]), .Z(signal_3517)
         );
  XOR2_X1 cell_1811_U3 ( .A(n376), .B(cell_1811_and_out[0]), .Z(signal_2079)
         );
  XOR2_X1 cell_1811_U2 ( .A(n378), .B(n365), .Z(cell_1811_and_in[1]) );
  XOR2_X1 cell_1811_U1 ( .A(n376), .B(n363), .Z(cell_1811_and_in[0]) );
  XOR2_X1 cell_1811_a_HPC2_and_U14 ( .A(Fresh[97]), .B(cell_1811_and_in[0]), 
        .Z(cell_1811_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1811_a_HPC2_and_U13 ( .A(Fresh[97]), .B(cell_1811_and_in[1]), 
        .Z(cell_1811_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1811_a_HPC2_and_U12 ( .A1(cell_1811_a_HPC2_and_a_reg[1]), .A2(
        cell_1811_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1811_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1811_a_HPC2_and_U11 ( .A1(cell_1811_a_HPC2_and_a_reg[0]), .A2(
        cell_1811_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1811_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1811_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1811_a_HPC2_and_n9), 
        .ZN(cell_1811_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1811_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1811_a_HPC2_and_n9), 
        .ZN(cell_1811_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1811_a_HPC2_and_U8 ( .A(Fresh[97]), .ZN(cell_1811_a_HPC2_and_n9)
         );
  AND2_X1 cell_1811_a_HPC2_and_U7 ( .A1(cell_1811_and_in[1]), .A2(n418), .ZN(
        cell_1811_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1811_a_HPC2_and_U6 ( .A1(cell_1811_and_in[0]), .A2(n401), .ZN(
        cell_1811_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1811_a_HPC2_and_U5 ( .A(cell_1811_a_HPC2_and_n8), .B(
        cell_1811_a_HPC2_and_z_1__1_), .ZN(cell_1811_and_out[1]) );
  XNOR2_X1 cell_1811_a_HPC2_and_U4 ( .A(
        cell_1811_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1811_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1811_a_HPC2_and_n8) );
  XNOR2_X1 cell_1811_a_HPC2_and_U3 ( .A(cell_1811_a_HPC2_and_n7), .B(
        cell_1811_a_HPC2_and_z_0__0_), .ZN(cell_1811_and_out[0]) );
  XNOR2_X1 cell_1811_a_HPC2_and_U2 ( .A(
        cell_1811_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1811_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1811_a_HPC2_and_n7) );
  DFF_X1 cell_1811_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1811_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1811_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1811_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1811_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1811_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1811_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1811_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1811_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1811_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1812_U4 ( .A(signal_3404), .B(cell_1812_and_out[1]), .Z(
        signal_3518) );
  XOR2_X1 cell_1812_U3 ( .A(signal_1990), .B(cell_1812_and_out[0]), .Z(
        signal_2080) );
  XOR2_X1 cell_1812_U2 ( .A(signal_3404), .B(signal_3432), .Z(
        cell_1812_and_in[1]) );
  XOR2_X1 cell_1812_U1 ( .A(signal_1990), .B(signal_2018), .Z(
        cell_1812_and_in[0]) );
  XOR2_X1 cell_1812_a_HPC2_and_U14 ( .A(Fresh[98]), .B(cell_1812_and_in[0]), 
        .Z(cell_1812_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1812_a_HPC2_and_U13 ( .A(Fresh[98]), .B(cell_1812_and_in[1]), 
        .Z(cell_1812_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1812_a_HPC2_and_U12 ( .A1(cell_1812_a_HPC2_and_a_reg[1]), .A2(
        cell_1812_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1812_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1812_a_HPC2_and_U11 ( .A1(cell_1812_a_HPC2_and_a_reg[0]), .A2(
        cell_1812_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1812_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1812_a_HPC2_and_U10 ( .A1(n450), .A2(cell_1812_a_HPC2_and_n9), 
        .ZN(cell_1812_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1812_a_HPC2_and_U9 ( .A1(n436), .A2(cell_1812_a_HPC2_and_n9), 
        .ZN(cell_1812_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1812_a_HPC2_and_U8 ( .A(Fresh[98]), .ZN(cell_1812_a_HPC2_and_n9)
         );
  AND2_X1 cell_1812_a_HPC2_and_U7 ( .A1(cell_1812_and_in[1]), .A2(n450), .ZN(
        cell_1812_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1812_a_HPC2_and_U6 ( .A1(cell_1812_and_in[0]), .A2(n436), .ZN(
        cell_1812_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1812_a_HPC2_and_U5 ( .A(cell_1812_a_HPC2_and_n8), .B(
        cell_1812_a_HPC2_and_z_1__1_), .ZN(cell_1812_and_out[1]) );
  XNOR2_X1 cell_1812_a_HPC2_and_U4 ( .A(
        cell_1812_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1812_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1812_a_HPC2_and_n8) );
  XNOR2_X1 cell_1812_a_HPC2_and_U3 ( .A(cell_1812_a_HPC2_and_n7), .B(
        cell_1812_a_HPC2_and_z_0__0_), .ZN(cell_1812_and_out[0]) );
  XNOR2_X1 cell_1812_a_HPC2_and_U2 ( .A(
        cell_1812_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1812_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1812_a_HPC2_and_n7) );
  DFF_X1 cell_1812_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1812_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1812_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_1812_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1812_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1812_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_1812_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1812_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1812_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1812_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1813_U4 ( .A(n364), .B(cell_1813_and_out[1]), .Z(signal_3519)
         );
  XOR2_X1 cell_1813_U3 ( .A(n362), .B(cell_1813_and_out[0]), .Z(signal_2081)
         );
  XOR2_X1 cell_1813_U2 ( .A(n364), .B(1'b0), .Z(cell_1813_and_in[1]) );
  XOR2_X1 cell_1813_U1 ( .A(n362), .B(1'b1), .Z(cell_1813_and_in[0]) );
  XOR2_X1 cell_1813_a_HPC2_and_U14 ( .A(Fresh[99]), .B(cell_1813_and_in[0]), 
        .Z(cell_1813_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1813_a_HPC2_and_U13 ( .A(Fresh[99]), .B(cell_1813_and_in[1]), 
        .Z(cell_1813_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1813_a_HPC2_and_U12 ( .A1(cell_1813_a_HPC2_and_a_reg[1]), .A2(
        cell_1813_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1813_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1813_a_HPC2_and_U11 ( .A1(cell_1813_a_HPC2_and_a_reg[0]), .A2(
        cell_1813_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1813_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1813_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1813_a_HPC2_and_n9), 
        .ZN(cell_1813_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1813_a_HPC2_and_U9 ( .A1(n398), .A2(cell_1813_a_HPC2_and_n9), 
        .ZN(cell_1813_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1813_a_HPC2_and_U8 ( .A(Fresh[99]), .ZN(cell_1813_a_HPC2_and_n9)
         );
  AND2_X1 cell_1813_a_HPC2_and_U7 ( .A1(cell_1813_and_in[1]), .A2(n422), .ZN(
        cell_1813_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1813_a_HPC2_and_U6 ( .A1(cell_1813_and_in[0]), .A2(n398), .ZN(
        cell_1813_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1813_a_HPC2_and_U5 ( .A(cell_1813_a_HPC2_and_n8), .B(
        cell_1813_a_HPC2_and_z_1__1_), .ZN(cell_1813_and_out[1]) );
  XNOR2_X1 cell_1813_a_HPC2_and_U4 ( .A(
        cell_1813_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1813_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1813_a_HPC2_and_n8) );
  XNOR2_X1 cell_1813_a_HPC2_and_U3 ( .A(cell_1813_a_HPC2_and_n7), .B(
        cell_1813_a_HPC2_and_z_0__0_), .ZN(cell_1813_and_out[0]) );
  XNOR2_X1 cell_1813_a_HPC2_and_U2 ( .A(
        cell_1813_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1813_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1813_a_HPC2_and_n7) );
  DFF_X1 cell_1813_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1813_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1813_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n398), .CK(clk), 
        .Q(cell_1813_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1813_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1813_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1813_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1813_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1813_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1813_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1814_U4 ( .A(1'b0), .B(cell_1814_and_out[1]), .Z(signal_3520)
         );
  XOR2_X1 cell_1814_U3 ( .A(1'b1), .B(cell_1814_and_out[0]), .Z(signal_2082)
         );
  XOR2_X1 cell_1814_U2 ( .A(1'b0), .B(signal_3424), .Z(cell_1814_and_in[1]) );
  XOR2_X1 cell_1814_U1 ( .A(1'b1), .B(signal_2010), .Z(cell_1814_and_in[0]) );
  XOR2_X1 cell_1814_a_HPC2_and_U14 ( .A(Fresh[100]), .B(cell_1814_and_in[0]), 
        .Z(cell_1814_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1814_a_HPC2_and_U13 ( .A(Fresh[100]), .B(cell_1814_and_in[1]), 
        .Z(cell_1814_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1814_a_HPC2_and_U12 ( .A1(cell_1814_a_HPC2_and_a_reg[1]), .A2(
        cell_1814_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1814_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1814_a_HPC2_and_U11 ( .A1(cell_1814_a_HPC2_and_a_reg[0]), .A2(
        cell_1814_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1814_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1814_a_HPC2_and_U10 ( .A1(n415), .A2(cell_1814_a_HPC2_and_n9), 
        .ZN(cell_1814_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1814_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1814_a_HPC2_and_n9), 
        .ZN(cell_1814_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1814_a_HPC2_and_U8 ( .A(Fresh[100]), .ZN(cell_1814_a_HPC2_and_n9) );
  AND2_X1 cell_1814_a_HPC2_and_U7 ( .A1(cell_1814_and_in[1]), .A2(n415), .ZN(
        cell_1814_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1814_a_HPC2_and_U6 ( .A1(cell_1814_and_in[0]), .A2(n405), .ZN(
        cell_1814_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1814_a_HPC2_and_U5 ( .A(cell_1814_a_HPC2_and_n8), .B(
        cell_1814_a_HPC2_and_z_1__1_), .ZN(cell_1814_and_out[1]) );
  XNOR2_X1 cell_1814_a_HPC2_and_U4 ( .A(
        cell_1814_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1814_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1814_a_HPC2_and_n8) );
  XNOR2_X1 cell_1814_a_HPC2_and_U3 ( .A(cell_1814_a_HPC2_and_n7), .B(
        cell_1814_a_HPC2_and_z_0__0_), .ZN(cell_1814_and_out[0]) );
  XNOR2_X1 cell_1814_a_HPC2_and_U2 ( .A(
        cell_1814_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1814_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1814_a_HPC2_and_n7) );
  DFF_X1 cell_1814_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1814_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1814_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1814_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1814_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1814_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n415), .CK(clk), 
        .Q(cell_1814_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1814_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1814_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1814_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1815_U4 ( .A(n381), .B(cell_1815_and_out[1]), .Z(signal_3521)
         );
  XOR2_X1 cell_1815_U3 ( .A(n380), .B(cell_1815_and_out[0]), .Z(signal_2083)
         );
  XOR2_X1 cell_1815_U2 ( .A(n381), .B(signal_3426), .Z(cell_1815_and_in[1]) );
  XOR2_X1 cell_1815_U1 ( .A(n380), .B(signal_2012), .Z(cell_1815_and_in[0]) );
  XOR2_X1 cell_1815_a_HPC2_and_U14 ( .A(Fresh[101]), .B(cell_1815_and_in[0]), 
        .Z(cell_1815_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1815_a_HPC2_and_U13 ( .A(Fresh[101]), .B(cell_1815_and_in[1]), 
        .Z(cell_1815_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1815_a_HPC2_and_U12 ( .A1(cell_1815_a_HPC2_and_a_reg[1]), .A2(
        cell_1815_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1815_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1815_a_HPC2_and_U11 ( .A1(cell_1815_a_HPC2_and_a_reg[0]), .A2(
        cell_1815_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1815_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1815_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1815_a_HPC2_and_n9), 
        .ZN(cell_1815_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1815_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1815_a_HPC2_and_n9), 
        .ZN(cell_1815_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1815_a_HPC2_and_U8 ( .A(Fresh[101]), .ZN(cell_1815_a_HPC2_and_n9) );
  AND2_X1 cell_1815_a_HPC2_and_U7 ( .A1(cell_1815_and_in[1]), .A2(n418), .ZN(
        cell_1815_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1815_a_HPC2_and_U6 ( .A1(cell_1815_and_in[0]), .A2(n401), .ZN(
        cell_1815_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1815_a_HPC2_and_U5 ( .A(cell_1815_a_HPC2_and_n8), .B(
        cell_1815_a_HPC2_and_z_1__1_), .ZN(cell_1815_and_out[1]) );
  XNOR2_X1 cell_1815_a_HPC2_and_U4 ( .A(
        cell_1815_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1815_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1815_a_HPC2_and_n8) );
  XNOR2_X1 cell_1815_a_HPC2_and_U3 ( .A(cell_1815_a_HPC2_and_n7), .B(
        cell_1815_a_HPC2_and_z_0__0_), .ZN(cell_1815_and_out[0]) );
  XNOR2_X1 cell_1815_a_HPC2_and_U2 ( .A(
        cell_1815_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1815_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1815_a_HPC2_and_n7) );
  DFF_X1 cell_1815_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1815_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1815_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1815_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1815_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1815_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1815_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1815_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1815_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1815_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1816_U4 ( .A(n378), .B(cell_1816_and_out[1]), .Z(signal_3522)
         );
  XOR2_X1 cell_1816_U3 ( .A(n376), .B(cell_1816_and_out[0]), .Z(signal_2084)
         );
  XOR2_X1 cell_1816_U2 ( .A(n378), .B(n361), .Z(cell_1816_and_in[1]) );
  XOR2_X1 cell_1816_U1 ( .A(n376), .B(n359), .Z(cell_1816_and_in[0]) );
  XOR2_X1 cell_1816_a_HPC2_and_U14 ( .A(Fresh[102]), .B(cell_1816_and_in[0]), 
        .Z(cell_1816_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1816_a_HPC2_and_U13 ( .A(Fresh[102]), .B(cell_1816_and_in[1]), 
        .Z(cell_1816_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1816_a_HPC2_and_U12 ( .A1(cell_1816_a_HPC2_and_a_reg[1]), .A2(
        cell_1816_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1816_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1816_a_HPC2_and_U11 ( .A1(cell_1816_a_HPC2_and_a_reg[0]), .A2(
        cell_1816_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1816_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1816_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1816_a_HPC2_and_n9), 
        .ZN(cell_1816_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1816_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1816_a_HPC2_and_n9), 
        .ZN(cell_1816_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1816_a_HPC2_and_U8 ( .A(Fresh[102]), .ZN(cell_1816_a_HPC2_and_n9) );
  AND2_X1 cell_1816_a_HPC2_and_U7 ( .A1(cell_1816_and_in[1]), .A2(n418), .ZN(
        cell_1816_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1816_a_HPC2_and_U6 ( .A1(cell_1816_and_in[0]), .A2(n401), .ZN(
        cell_1816_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1816_a_HPC2_and_U5 ( .A(cell_1816_a_HPC2_and_n8), .B(
        cell_1816_a_HPC2_and_z_1__1_), .ZN(cell_1816_and_out[1]) );
  XNOR2_X1 cell_1816_a_HPC2_and_U4 ( .A(
        cell_1816_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1816_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1816_a_HPC2_and_n8) );
  XNOR2_X1 cell_1816_a_HPC2_and_U3 ( .A(cell_1816_a_HPC2_and_n7), .B(
        cell_1816_a_HPC2_and_z_0__0_), .ZN(cell_1816_and_out[0]) );
  XNOR2_X1 cell_1816_a_HPC2_and_U2 ( .A(
        cell_1816_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1816_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1816_a_HPC2_and_n7) );
  DFF_X1 cell_1816_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1816_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1816_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1816_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1816_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1816_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1816_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1816_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1816_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1816_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1817_U4 ( .A(n370), .B(cell_1817_and_out[1]), .Z(signal_3523)
         );
  XOR2_X1 cell_1817_U3 ( .A(n368), .B(cell_1817_and_out[0]), .Z(signal_2085)
         );
  XOR2_X1 cell_1817_U2 ( .A(n370), .B(n355), .Z(cell_1817_and_in[1]) );
  XOR2_X1 cell_1817_U1 ( .A(n368), .B(n353), .Z(cell_1817_and_in[0]) );
  XOR2_X1 cell_1817_a_HPC2_and_U14 ( .A(Fresh[103]), .B(cell_1817_and_in[0]), 
        .Z(cell_1817_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1817_a_HPC2_and_U13 ( .A(Fresh[103]), .B(cell_1817_and_in[1]), 
        .Z(cell_1817_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1817_a_HPC2_and_U12 ( .A1(cell_1817_a_HPC2_and_a_reg[1]), .A2(
        cell_1817_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1817_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1817_a_HPC2_and_U11 ( .A1(cell_1817_a_HPC2_and_a_reg[0]), .A2(
        cell_1817_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1817_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1817_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1817_a_HPC2_and_n9), 
        .ZN(cell_1817_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1817_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1817_a_HPC2_and_n9), 
        .ZN(cell_1817_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1817_a_HPC2_and_U8 ( .A(Fresh[103]), .ZN(cell_1817_a_HPC2_and_n9) );
  AND2_X1 cell_1817_a_HPC2_and_U7 ( .A1(cell_1817_and_in[1]), .A2(n418), .ZN(
        cell_1817_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1817_a_HPC2_and_U6 ( .A1(cell_1817_and_in[0]), .A2(n401), .ZN(
        cell_1817_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1817_a_HPC2_and_U5 ( .A(cell_1817_a_HPC2_and_n8), .B(
        cell_1817_a_HPC2_and_z_1__1_), .ZN(cell_1817_and_out[1]) );
  XNOR2_X1 cell_1817_a_HPC2_and_U4 ( .A(
        cell_1817_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1817_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1817_a_HPC2_and_n8) );
  XNOR2_X1 cell_1817_a_HPC2_and_U3 ( .A(cell_1817_a_HPC2_and_n7), .B(
        cell_1817_a_HPC2_and_z_0__0_), .ZN(cell_1817_and_out[0]) );
  XNOR2_X1 cell_1817_a_HPC2_and_U2 ( .A(
        cell_1817_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1817_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1817_a_HPC2_and_n7) );
  DFF_X1 cell_1817_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1817_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1817_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1817_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1817_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1817_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1817_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1817_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1817_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1817_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1818_U4 ( .A(n374), .B(cell_1818_and_out[1]), .Z(signal_3524)
         );
  XOR2_X1 cell_1818_U3 ( .A(n372), .B(cell_1818_and_out[0]), .Z(signal_2086)
         );
  XOR2_X1 cell_1818_U2 ( .A(n374), .B(signal_3261), .Z(cell_1818_and_in[1]) );
  XOR2_X1 cell_1818_U1 ( .A(n372), .B(signal_1987), .Z(cell_1818_and_in[0]) );
  XOR2_X1 cell_1818_a_HPC2_and_U14 ( .A(Fresh[104]), .B(cell_1818_and_in[0]), 
        .Z(cell_1818_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1818_a_HPC2_and_U13 ( .A(Fresh[104]), .B(cell_1818_and_in[1]), 
        .Z(cell_1818_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1818_a_HPC2_and_U12 ( .A1(cell_1818_a_HPC2_and_a_reg[1]), .A2(
        cell_1818_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1818_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1818_a_HPC2_and_U11 ( .A1(cell_1818_a_HPC2_and_a_reg[0]), .A2(
        cell_1818_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1818_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1818_a_HPC2_and_U10 ( .A1(n418), .A2(cell_1818_a_HPC2_and_n9), 
        .ZN(cell_1818_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1818_a_HPC2_and_U9 ( .A1(n401), .A2(cell_1818_a_HPC2_and_n9), 
        .ZN(cell_1818_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1818_a_HPC2_and_U8 ( .A(Fresh[104]), .ZN(cell_1818_a_HPC2_and_n9) );
  AND2_X1 cell_1818_a_HPC2_and_U7 ( .A1(cell_1818_and_in[1]), .A2(n418), .ZN(
        cell_1818_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1818_a_HPC2_and_U6 ( .A1(cell_1818_and_in[0]), .A2(n401), .ZN(
        cell_1818_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1818_a_HPC2_and_U5 ( .A(cell_1818_a_HPC2_and_n8), .B(
        cell_1818_a_HPC2_and_z_1__1_), .ZN(cell_1818_and_out[1]) );
  XNOR2_X1 cell_1818_a_HPC2_and_U4 ( .A(
        cell_1818_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1818_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1818_a_HPC2_and_n8) );
  XNOR2_X1 cell_1818_a_HPC2_and_U3 ( .A(cell_1818_a_HPC2_and_n7), .B(
        cell_1818_a_HPC2_and_z_0__0_), .ZN(cell_1818_and_out[0]) );
  XNOR2_X1 cell_1818_a_HPC2_and_U2 ( .A(
        cell_1818_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1818_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1818_a_HPC2_and_n7) );
  DFF_X1 cell_1818_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1818_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1818_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n401), .CK(clk), 
        .Q(cell_1818_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1818_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1818_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n418), .CK(clk), 
        .Q(cell_1818_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1818_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1818_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1818_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1819_U4 ( .A(n367), .B(cell_1819_and_out[1]), .Z(signal_3525)
         );
  XOR2_X1 cell_1819_U3 ( .A(n366), .B(cell_1819_and_out[0]), .Z(signal_2087)
         );
  XOR2_X1 cell_1819_U2 ( .A(n367), .B(n355), .Z(cell_1819_and_in[1]) );
  XOR2_X1 cell_1819_U1 ( .A(n366), .B(n353), .Z(cell_1819_and_in[0]) );
  XOR2_X1 cell_1819_a_HPC2_and_U14 ( .A(Fresh[105]), .B(cell_1819_and_in[0]), 
        .Z(cell_1819_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1819_a_HPC2_and_U13 ( .A(Fresh[105]), .B(cell_1819_and_in[1]), 
        .Z(cell_1819_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1819_a_HPC2_and_U12 ( .A1(cell_1819_a_HPC2_and_a_reg[1]), .A2(
        cell_1819_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1819_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1819_a_HPC2_and_U11 ( .A1(cell_1819_a_HPC2_and_a_reg[0]), .A2(
        cell_1819_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1819_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1819_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1819_a_HPC2_and_n9), 
        .ZN(cell_1819_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1819_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1819_a_HPC2_and_n9), 
        .ZN(cell_1819_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1819_a_HPC2_and_U8 ( .A(Fresh[105]), .ZN(cell_1819_a_HPC2_and_n9) );
  AND2_X1 cell_1819_a_HPC2_and_U7 ( .A1(cell_1819_and_in[1]), .A2(n419), .ZN(
        cell_1819_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1819_a_HPC2_and_U6 ( .A1(cell_1819_and_in[0]), .A2(n402), .ZN(
        cell_1819_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1819_a_HPC2_and_U5 ( .A(cell_1819_a_HPC2_and_n8), .B(
        cell_1819_a_HPC2_and_z_1__1_), .ZN(cell_1819_and_out[1]) );
  XNOR2_X1 cell_1819_a_HPC2_and_U4 ( .A(
        cell_1819_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1819_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1819_a_HPC2_and_n8) );
  XNOR2_X1 cell_1819_a_HPC2_and_U3 ( .A(cell_1819_a_HPC2_and_n7), .B(
        cell_1819_a_HPC2_and_z_0__0_), .ZN(cell_1819_and_out[0]) );
  XNOR2_X1 cell_1819_a_HPC2_and_U2 ( .A(
        cell_1819_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1819_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1819_a_HPC2_and_n7) );
  DFF_X1 cell_1819_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1819_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1819_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1819_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1819_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1819_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1819_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1819_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1819_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1819_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1820_U4 ( .A(n371), .B(cell_1820_and_out[1]), .Z(signal_3526)
         );
  XOR2_X1 cell_1820_U3 ( .A(n369), .B(cell_1820_and_out[0]), .Z(signal_2088)
         );
  XOR2_X1 cell_1820_U2 ( .A(n371), .B(n389), .Z(cell_1820_and_in[1]) );
  XOR2_X1 cell_1820_U1 ( .A(n369), .B(n388), .Z(cell_1820_and_in[0]) );
  XOR2_X1 cell_1820_a_HPC2_and_U14 ( .A(Fresh[106]), .B(cell_1820_and_in[0]), 
        .Z(cell_1820_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1820_a_HPC2_and_U13 ( .A(Fresh[106]), .B(cell_1820_and_in[1]), 
        .Z(cell_1820_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1820_a_HPC2_and_U12 ( .A1(cell_1820_a_HPC2_and_a_reg[1]), .A2(
        cell_1820_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1820_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1820_a_HPC2_and_U11 ( .A1(cell_1820_a_HPC2_and_a_reg[0]), .A2(
        cell_1820_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1820_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1820_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1820_a_HPC2_and_n9), 
        .ZN(cell_1820_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1820_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1820_a_HPC2_and_n9), 
        .ZN(cell_1820_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1820_a_HPC2_and_U8 ( .A(Fresh[106]), .ZN(cell_1820_a_HPC2_and_n9) );
  AND2_X1 cell_1820_a_HPC2_and_U7 ( .A1(cell_1820_and_in[1]), .A2(n419), .ZN(
        cell_1820_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1820_a_HPC2_and_U6 ( .A1(cell_1820_and_in[0]), .A2(n402), .ZN(
        cell_1820_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1820_a_HPC2_and_U5 ( .A(cell_1820_a_HPC2_and_n8), .B(
        cell_1820_a_HPC2_and_z_1__1_), .ZN(cell_1820_and_out[1]) );
  XNOR2_X1 cell_1820_a_HPC2_and_U4 ( .A(
        cell_1820_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1820_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1820_a_HPC2_and_n8) );
  XNOR2_X1 cell_1820_a_HPC2_and_U3 ( .A(cell_1820_a_HPC2_and_n7), .B(
        cell_1820_a_HPC2_and_z_0__0_), .ZN(cell_1820_and_out[0]) );
  XNOR2_X1 cell_1820_a_HPC2_and_U2 ( .A(
        cell_1820_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1820_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1820_a_HPC2_and_n7) );
  DFF_X1 cell_1820_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1820_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1820_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1820_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1820_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1820_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1820_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1820_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1820_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1820_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1821_U4 ( .A(n354), .B(cell_1821_and_out[1]), .Z(signal_3527)
         );
  XOR2_X1 cell_1821_U3 ( .A(n352), .B(cell_1821_and_out[0]), .Z(signal_2089)
         );
  XOR2_X1 cell_1821_U2 ( .A(n354), .B(n365), .Z(cell_1821_and_in[1]) );
  XOR2_X1 cell_1821_U1 ( .A(n352), .B(n363), .Z(cell_1821_and_in[0]) );
  XOR2_X1 cell_1821_a_HPC2_and_U14 ( .A(Fresh[107]), .B(cell_1821_and_in[0]), 
        .Z(cell_1821_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1821_a_HPC2_and_U13 ( .A(Fresh[107]), .B(cell_1821_and_in[1]), 
        .Z(cell_1821_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1821_a_HPC2_and_U12 ( .A1(cell_1821_a_HPC2_and_a_reg[1]), .A2(
        cell_1821_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1821_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1821_a_HPC2_and_U11 ( .A1(cell_1821_a_HPC2_and_a_reg[0]), .A2(
        cell_1821_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1821_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1821_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1821_a_HPC2_and_n9), 
        .ZN(cell_1821_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1821_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1821_a_HPC2_and_n9), 
        .ZN(cell_1821_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1821_a_HPC2_and_U8 ( .A(Fresh[107]), .ZN(cell_1821_a_HPC2_and_n9) );
  AND2_X1 cell_1821_a_HPC2_and_U7 ( .A1(cell_1821_and_in[1]), .A2(n419), .ZN(
        cell_1821_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1821_a_HPC2_and_U6 ( .A1(cell_1821_and_in[0]), .A2(n402), .ZN(
        cell_1821_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1821_a_HPC2_and_U5 ( .A(cell_1821_a_HPC2_and_n8), .B(
        cell_1821_a_HPC2_and_z_1__1_), .ZN(cell_1821_and_out[1]) );
  XNOR2_X1 cell_1821_a_HPC2_and_U4 ( .A(
        cell_1821_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1821_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1821_a_HPC2_and_n8) );
  XNOR2_X1 cell_1821_a_HPC2_and_U3 ( .A(cell_1821_a_HPC2_and_n7), .B(
        cell_1821_a_HPC2_and_z_0__0_), .ZN(cell_1821_and_out[0]) );
  XNOR2_X1 cell_1821_a_HPC2_and_U2 ( .A(
        cell_1821_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1821_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1821_a_HPC2_and_n7) );
  DFF_X1 cell_1821_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1821_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1821_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1821_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1821_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1821_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1821_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1821_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1821_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1821_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1822_U4 ( .A(n354), .B(cell_1822_and_out[1]), .Z(signal_3528)
         );
  XOR2_X1 cell_1822_U3 ( .A(n352), .B(cell_1822_and_out[0]), .Z(signal_2090)
         );
  XOR2_X1 cell_1822_U2 ( .A(n354), .B(signal_3413), .Z(cell_1822_and_in[1]) );
  XOR2_X1 cell_1822_U1 ( .A(n352), .B(signal_1999), .Z(cell_1822_and_in[0]) );
  XOR2_X1 cell_1822_a_HPC2_and_U14 ( .A(Fresh[108]), .B(cell_1822_and_in[0]), 
        .Z(cell_1822_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1822_a_HPC2_and_U13 ( .A(Fresh[108]), .B(cell_1822_and_in[1]), 
        .Z(cell_1822_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1822_a_HPC2_and_U12 ( .A1(cell_1822_a_HPC2_and_a_reg[1]), .A2(
        cell_1822_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1822_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1822_a_HPC2_and_U11 ( .A1(cell_1822_a_HPC2_and_a_reg[0]), .A2(
        cell_1822_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1822_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1822_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1822_a_HPC2_and_n9), 
        .ZN(cell_1822_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1822_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1822_a_HPC2_and_n9), 
        .ZN(cell_1822_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1822_a_HPC2_and_U8 ( .A(Fresh[108]), .ZN(cell_1822_a_HPC2_and_n9) );
  AND2_X1 cell_1822_a_HPC2_and_U7 ( .A1(cell_1822_and_in[1]), .A2(n419), .ZN(
        cell_1822_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1822_a_HPC2_and_U6 ( .A1(cell_1822_and_in[0]), .A2(n402), .ZN(
        cell_1822_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1822_a_HPC2_and_U5 ( .A(cell_1822_a_HPC2_and_n8), .B(
        cell_1822_a_HPC2_and_z_1__1_), .ZN(cell_1822_and_out[1]) );
  XNOR2_X1 cell_1822_a_HPC2_and_U4 ( .A(
        cell_1822_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1822_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1822_a_HPC2_and_n8) );
  XNOR2_X1 cell_1822_a_HPC2_and_U3 ( .A(cell_1822_a_HPC2_and_n7), .B(
        cell_1822_a_HPC2_and_z_0__0_), .ZN(cell_1822_and_out[0]) );
  XNOR2_X1 cell_1822_a_HPC2_and_U2 ( .A(
        cell_1822_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1822_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1822_a_HPC2_and_n7) );
  DFF_X1 cell_1822_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1822_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1822_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1822_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1822_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1822_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1822_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1822_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1822_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1822_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1823_U4 ( .A(n386), .B(cell_1823_and_out[1]), .Z(signal_3529)
         );
  XOR2_X1 cell_1823_U3 ( .A(n384), .B(cell_1823_and_out[0]), .Z(signal_2091)
         );
  XOR2_X1 cell_1823_U2 ( .A(n386), .B(signal_3406), .Z(cell_1823_and_in[1]) );
  XOR2_X1 cell_1823_U1 ( .A(n384), .B(signal_1992), .Z(cell_1823_and_in[0]) );
  XOR2_X1 cell_1823_a_HPC2_and_U14 ( .A(Fresh[109]), .B(cell_1823_and_in[0]), 
        .Z(cell_1823_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1823_a_HPC2_and_U13 ( .A(Fresh[109]), .B(cell_1823_and_in[1]), 
        .Z(cell_1823_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1823_a_HPC2_and_U12 ( .A1(cell_1823_a_HPC2_and_a_reg[1]), .A2(
        cell_1823_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1823_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1823_a_HPC2_and_U11 ( .A1(cell_1823_a_HPC2_and_a_reg[0]), .A2(
        cell_1823_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1823_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1823_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1823_a_HPC2_and_n9), 
        .ZN(cell_1823_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1823_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1823_a_HPC2_and_n9), 
        .ZN(cell_1823_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1823_a_HPC2_and_U8 ( .A(Fresh[109]), .ZN(cell_1823_a_HPC2_and_n9) );
  AND2_X1 cell_1823_a_HPC2_and_U7 ( .A1(cell_1823_and_in[1]), .A2(n419), .ZN(
        cell_1823_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1823_a_HPC2_and_U6 ( .A1(cell_1823_and_in[0]), .A2(n402), .ZN(
        cell_1823_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1823_a_HPC2_and_U5 ( .A(cell_1823_a_HPC2_and_n8), .B(
        cell_1823_a_HPC2_and_z_1__1_), .ZN(cell_1823_and_out[1]) );
  XNOR2_X1 cell_1823_a_HPC2_and_U4 ( .A(
        cell_1823_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1823_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1823_a_HPC2_and_n8) );
  XNOR2_X1 cell_1823_a_HPC2_and_U3 ( .A(cell_1823_a_HPC2_and_n7), .B(
        cell_1823_a_HPC2_and_z_0__0_), .ZN(cell_1823_and_out[0]) );
  XNOR2_X1 cell_1823_a_HPC2_and_U2 ( .A(
        cell_1823_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1823_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1823_a_HPC2_and_n7) );
  DFF_X1 cell_1823_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1823_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1823_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1823_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1823_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1823_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1823_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1823_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1823_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1823_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1824_U6 ( .A(cell_1824_n4), .B(cell_1824_and_out[1]), .Z(
        signal_3530) );
  XOR2_X1 cell_1824_U5 ( .A(cell_1824_n3), .B(cell_1824_and_out[0]), .Z(
        signal_2092) );
  XOR2_X1 cell_1824_U4 ( .A(cell_1824_n4), .B(1'b0), .Z(cell_1824_and_in[1])
         );
  XOR2_X1 cell_1824_U3 ( .A(cell_1824_n3), .B(1'b0), .Z(cell_1824_and_in[0])
         );
  BUF_X1 cell_1824_U2 ( .A(signal_3426), .Z(cell_1824_n4) );
  BUF_X1 cell_1824_U1 ( .A(signal_2012), .Z(cell_1824_n3) );
  XOR2_X1 cell_1824_a_HPC2_and_U14 ( .A(Fresh[110]), .B(cell_1824_and_in[0]), 
        .Z(cell_1824_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1824_a_HPC2_and_U13 ( .A(Fresh[110]), .B(cell_1824_and_in[1]), 
        .Z(cell_1824_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1824_a_HPC2_and_U12 ( .A1(cell_1824_a_HPC2_and_a_reg[1]), .A2(
        cell_1824_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1824_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1824_a_HPC2_and_U11 ( .A1(cell_1824_a_HPC2_and_a_reg[0]), .A2(
        cell_1824_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1824_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1824_a_HPC2_and_U10 ( .A1(n413), .A2(cell_1824_a_HPC2_and_n9), 
        .ZN(cell_1824_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1824_a_HPC2_and_U9 ( .A1(n396), .A2(cell_1824_a_HPC2_and_n9), 
        .ZN(cell_1824_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1824_a_HPC2_and_U8 ( .A(Fresh[110]), .ZN(cell_1824_a_HPC2_and_n9) );
  AND2_X1 cell_1824_a_HPC2_and_U7 ( .A1(cell_1824_and_in[1]), .A2(n413), .ZN(
        cell_1824_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1824_a_HPC2_and_U6 ( .A1(cell_1824_and_in[0]), .A2(n396), .ZN(
        cell_1824_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1824_a_HPC2_and_U5 ( .A(cell_1824_a_HPC2_and_n8), .B(
        cell_1824_a_HPC2_and_z_1__1_), .ZN(cell_1824_and_out[1]) );
  XNOR2_X1 cell_1824_a_HPC2_and_U4 ( .A(
        cell_1824_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1824_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1824_a_HPC2_and_n8) );
  XNOR2_X1 cell_1824_a_HPC2_and_U3 ( .A(cell_1824_a_HPC2_and_n7), .B(
        cell_1824_a_HPC2_and_z_0__0_), .ZN(cell_1824_and_out[0]) );
  XNOR2_X1 cell_1824_a_HPC2_and_U2 ( .A(
        cell_1824_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1824_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1824_a_HPC2_and_n7) );
  DFF_X1 cell_1824_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1824_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1824_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n396), .CK(clk), 
        .Q(cell_1824_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1824_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1824_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n413), .CK(clk), 
        .Q(cell_1824_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1824_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1824_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1824_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1825_U4 ( .A(1'b0), .B(cell_1825_and_out[1]), .Z(signal_3531)
         );
  XOR2_X1 cell_1825_U3 ( .A(1'b1), .B(cell_1825_and_out[0]), .Z(signal_2093)
         );
  XOR2_X1 cell_1825_U2 ( .A(1'b0), .B(n365), .Z(cell_1825_and_in[1]) );
  XOR2_X1 cell_1825_U1 ( .A(1'b1), .B(n363), .Z(cell_1825_and_in[0]) );
  XOR2_X1 cell_1825_a_HPC2_and_U14 ( .A(Fresh[111]), .B(cell_1825_and_in[0]), 
        .Z(cell_1825_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1825_a_HPC2_and_U13 ( .A(Fresh[111]), .B(cell_1825_and_in[1]), 
        .Z(cell_1825_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1825_a_HPC2_and_U12 ( .A1(cell_1825_a_HPC2_and_a_reg[1]), .A2(
        cell_1825_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1825_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1825_a_HPC2_and_U11 ( .A1(cell_1825_a_HPC2_and_a_reg[0]), .A2(
        cell_1825_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1825_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1825_a_HPC2_and_U10 ( .A1(signal_3237), .A2(
        cell_1825_a_HPC2_and_n9), .ZN(cell_1825_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1825_a_HPC2_and_U9 ( .A1(signal_1512), .A2(
        cell_1825_a_HPC2_and_n9), .ZN(cell_1825_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1825_a_HPC2_and_U8 ( .A(Fresh[111]), .ZN(cell_1825_a_HPC2_and_n9) );
  AND2_X1 cell_1825_a_HPC2_and_U7 ( .A1(cell_1825_and_in[1]), .A2(signal_3237), 
        .ZN(cell_1825_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1825_a_HPC2_and_U6 ( .A1(cell_1825_and_in[0]), .A2(signal_1512), 
        .ZN(cell_1825_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1825_a_HPC2_and_U5 ( .A(cell_1825_a_HPC2_and_n8), .B(
        cell_1825_a_HPC2_and_z_1__1_), .ZN(cell_1825_and_out[1]) );
  XNOR2_X1 cell_1825_a_HPC2_and_U4 ( .A(
        cell_1825_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1825_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1825_a_HPC2_and_n8) );
  XNOR2_X1 cell_1825_a_HPC2_and_U3 ( .A(cell_1825_a_HPC2_and_n7), .B(
        cell_1825_a_HPC2_and_z_0__0_), .ZN(cell_1825_and_out[0]) );
  XNOR2_X1 cell_1825_a_HPC2_and_U2 ( .A(
        cell_1825_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1825_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1825_a_HPC2_and_n7) );
  DFF_X1 cell_1825_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1825_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1825_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1512), 
        .CK(clk), .Q(cell_1825_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1825_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1825_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3237), 
        .CK(clk), .Q(cell_1825_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1825_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1825_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1825_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1826_U4 ( .A(n381), .B(cell_1826_and_out[1]), .Z(signal_3532)
         );
  XOR2_X1 cell_1826_U3 ( .A(n380), .B(cell_1826_and_out[0]), .Z(signal_2094)
         );
  XOR2_X1 cell_1826_U2 ( .A(n381), .B(n371), .Z(cell_1826_and_in[1]) );
  XOR2_X1 cell_1826_U1 ( .A(n380), .B(n369), .Z(cell_1826_and_in[0]) );
  XOR2_X1 cell_1826_a_HPC2_and_U14 ( .A(Fresh[112]), .B(cell_1826_and_in[0]), 
        .Z(cell_1826_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1826_a_HPC2_and_U13 ( .A(Fresh[112]), .B(cell_1826_and_in[1]), 
        .Z(cell_1826_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1826_a_HPC2_and_U12 ( .A1(cell_1826_a_HPC2_and_a_reg[1]), .A2(
        cell_1826_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1826_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1826_a_HPC2_and_U11 ( .A1(cell_1826_a_HPC2_and_a_reg[0]), .A2(
        cell_1826_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1826_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1826_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1826_a_HPC2_and_n9), 
        .ZN(cell_1826_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1826_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1826_a_HPC2_and_n9), 
        .ZN(cell_1826_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1826_a_HPC2_and_U8 ( .A(Fresh[112]), .ZN(cell_1826_a_HPC2_and_n9) );
  AND2_X1 cell_1826_a_HPC2_and_U7 ( .A1(cell_1826_and_in[1]), .A2(n419), .ZN(
        cell_1826_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1826_a_HPC2_and_U6 ( .A1(cell_1826_and_in[0]), .A2(n402), .ZN(
        cell_1826_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1826_a_HPC2_and_U5 ( .A(cell_1826_a_HPC2_and_n8), .B(
        cell_1826_a_HPC2_and_z_1__1_), .ZN(cell_1826_and_out[1]) );
  XNOR2_X1 cell_1826_a_HPC2_and_U4 ( .A(
        cell_1826_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1826_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1826_a_HPC2_and_n8) );
  XNOR2_X1 cell_1826_a_HPC2_and_U3 ( .A(cell_1826_a_HPC2_and_n7), .B(
        cell_1826_a_HPC2_and_z_0__0_), .ZN(cell_1826_and_out[0]) );
  XNOR2_X1 cell_1826_a_HPC2_and_U2 ( .A(
        cell_1826_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1826_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1826_a_HPC2_and_n7) );
  DFF_X1 cell_1826_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1826_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1826_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1826_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1826_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1826_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1826_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1826_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1826_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1826_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1827_U4 ( .A(n389), .B(cell_1827_and_out[1]), .Z(signal_3533)
         );
  XOR2_X1 cell_1827_U3 ( .A(n388), .B(cell_1827_and_out[0]), .Z(signal_2095)
         );
  XOR2_X1 cell_1827_U2 ( .A(n389), .B(n355), .Z(cell_1827_and_in[1]) );
  XOR2_X1 cell_1827_U1 ( .A(n388), .B(n353), .Z(cell_1827_and_in[0]) );
  XOR2_X1 cell_1827_a_HPC2_and_U14 ( .A(Fresh[113]), .B(cell_1827_and_in[0]), 
        .Z(cell_1827_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1827_a_HPC2_and_U13 ( .A(Fresh[113]), .B(cell_1827_and_in[1]), 
        .Z(cell_1827_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1827_a_HPC2_and_U12 ( .A1(cell_1827_a_HPC2_and_a_reg[1]), .A2(
        cell_1827_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1827_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1827_a_HPC2_and_U11 ( .A1(cell_1827_a_HPC2_and_a_reg[0]), .A2(
        cell_1827_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1827_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1827_a_HPC2_and_U10 ( .A1(n419), .A2(cell_1827_a_HPC2_and_n9), 
        .ZN(cell_1827_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1827_a_HPC2_and_U9 ( .A1(n402), .A2(cell_1827_a_HPC2_and_n9), 
        .ZN(cell_1827_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1827_a_HPC2_and_U8 ( .A(Fresh[113]), .ZN(cell_1827_a_HPC2_and_n9) );
  AND2_X1 cell_1827_a_HPC2_and_U7 ( .A1(cell_1827_and_in[1]), .A2(n419), .ZN(
        cell_1827_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1827_a_HPC2_and_U6 ( .A1(cell_1827_and_in[0]), .A2(n402), .ZN(
        cell_1827_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1827_a_HPC2_and_U5 ( .A(cell_1827_a_HPC2_and_n8), .B(
        cell_1827_a_HPC2_and_z_1__1_), .ZN(cell_1827_and_out[1]) );
  XNOR2_X1 cell_1827_a_HPC2_and_U4 ( .A(
        cell_1827_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1827_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1827_a_HPC2_and_n8) );
  XNOR2_X1 cell_1827_a_HPC2_and_U3 ( .A(cell_1827_a_HPC2_and_n7), .B(
        cell_1827_a_HPC2_and_z_0__0_), .ZN(cell_1827_and_out[0]) );
  XNOR2_X1 cell_1827_a_HPC2_and_U2 ( .A(
        cell_1827_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1827_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1827_a_HPC2_and_n7) );
  DFF_X1 cell_1827_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1827_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1827_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n402), .CK(clk), 
        .Q(cell_1827_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1827_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1827_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n419), .CK(clk), 
        .Q(cell_1827_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1827_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1827_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1827_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1828_U4 ( .A(n357), .B(cell_1828_and_out[1]), .Z(signal_3534)
         );
  XOR2_X1 cell_1828_U3 ( .A(n356), .B(cell_1828_and_out[0]), .Z(signal_2096)
         );
  XOR2_X1 cell_1828_U2 ( .A(n357), .B(n355), .Z(cell_1828_and_in[1]) );
  XOR2_X1 cell_1828_U1 ( .A(n356), .B(n353), .Z(cell_1828_and_in[0]) );
  XOR2_X1 cell_1828_a_HPC2_and_U14 ( .A(Fresh[114]), .B(cell_1828_and_in[0]), 
        .Z(cell_1828_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1828_a_HPC2_and_U13 ( .A(Fresh[114]), .B(cell_1828_and_in[1]), 
        .Z(cell_1828_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1828_a_HPC2_and_U12 ( .A1(cell_1828_a_HPC2_and_a_reg[1]), .A2(
        cell_1828_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1828_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1828_a_HPC2_and_U11 ( .A1(cell_1828_a_HPC2_and_a_reg[0]), .A2(
        cell_1828_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1828_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1828_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1828_a_HPC2_and_n9), 
        .ZN(cell_1828_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1828_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1828_a_HPC2_and_n9), 
        .ZN(cell_1828_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1828_a_HPC2_and_U8 ( .A(Fresh[114]), .ZN(cell_1828_a_HPC2_and_n9) );
  AND2_X1 cell_1828_a_HPC2_and_U7 ( .A1(cell_1828_and_in[1]), .A2(n420), .ZN(
        cell_1828_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1828_a_HPC2_and_U6 ( .A1(cell_1828_and_in[0]), .A2(n403), .ZN(
        cell_1828_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1828_a_HPC2_and_U5 ( .A(cell_1828_a_HPC2_and_n8), .B(
        cell_1828_a_HPC2_and_z_1__1_), .ZN(cell_1828_and_out[1]) );
  XNOR2_X1 cell_1828_a_HPC2_and_U4 ( .A(
        cell_1828_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1828_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1828_a_HPC2_and_n8) );
  XNOR2_X1 cell_1828_a_HPC2_and_U3 ( .A(cell_1828_a_HPC2_and_n7), .B(
        cell_1828_a_HPC2_and_z_0__0_), .ZN(cell_1828_and_out[0]) );
  XNOR2_X1 cell_1828_a_HPC2_and_U2 ( .A(
        cell_1828_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1828_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1828_a_HPC2_and_n7) );
  DFF_X1 cell_1828_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1828_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1828_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1828_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1828_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1828_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1828_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1828_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1828_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1828_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1829_U4 ( .A(signal_3418), .B(cell_1829_and_out[1]), .Z(
        signal_3535) );
  XOR2_X1 cell_1829_U3 ( .A(signal_2004), .B(cell_1829_and_out[0]), .Z(
        signal_2097) );
  XOR2_X1 cell_1829_U2 ( .A(signal_3418), .B(signal_3258), .Z(
        cell_1829_and_in[1]) );
  XOR2_X1 cell_1829_U1 ( .A(signal_2004), .B(signal_1984), .Z(
        cell_1829_and_in[0]) );
  XOR2_X1 cell_1829_a_HPC2_and_U14 ( .A(Fresh[115]), .B(cell_1829_and_in[0]), 
        .Z(cell_1829_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1829_a_HPC2_and_U13 ( .A(Fresh[115]), .B(cell_1829_and_in[1]), 
        .Z(cell_1829_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1829_a_HPC2_and_U12 ( .A1(cell_1829_a_HPC2_and_a_reg[1]), .A2(
        cell_1829_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1829_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1829_a_HPC2_and_U11 ( .A1(cell_1829_a_HPC2_and_a_reg[0]), .A2(
        cell_1829_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1829_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1829_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1829_a_HPC2_and_n9), 
        .ZN(cell_1829_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1829_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1829_a_HPC2_and_n9), 
        .ZN(cell_1829_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1829_a_HPC2_and_U8 ( .A(Fresh[115]), .ZN(cell_1829_a_HPC2_and_n9) );
  AND2_X1 cell_1829_a_HPC2_and_U7 ( .A1(cell_1829_and_in[1]), .A2(n442), .ZN(
        cell_1829_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1829_a_HPC2_and_U6 ( .A1(cell_1829_and_in[0]), .A2(n428), .ZN(
        cell_1829_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1829_a_HPC2_and_U5 ( .A(cell_1829_a_HPC2_and_n8), .B(
        cell_1829_a_HPC2_and_z_1__1_), .ZN(cell_1829_and_out[1]) );
  XNOR2_X1 cell_1829_a_HPC2_and_U4 ( .A(
        cell_1829_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1829_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1829_a_HPC2_and_n8) );
  XNOR2_X1 cell_1829_a_HPC2_and_U3 ( .A(cell_1829_a_HPC2_and_n7), .B(
        cell_1829_a_HPC2_and_z_0__0_), .ZN(cell_1829_and_out[0]) );
  XNOR2_X1 cell_1829_a_HPC2_and_U2 ( .A(
        cell_1829_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1829_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1829_a_HPC2_and_n7) );
  DFF_X1 cell_1829_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1829_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1829_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1829_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1829_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1829_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1829_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1829_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1829_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1829_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1830_U4 ( .A(signal_3406), .B(cell_1830_and_out[1]), .Z(
        signal_3536) );
  XOR2_X1 cell_1830_U3 ( .A(signal_1992), .B(cell_1830_and_out[0]), .Z(
        signal_2098) );
  XOR2_X1 cell_1830_U2 ( .A(signal_3406), .B(1'b0), .Z(cell_1830_and_in[1]) );
  XOR2_X1 cell_1830_U1 ( .A(signal_1992), .B(1'b0), .Z(cell_1830_and_in[0]) );
  XOR2_X1 cell_1830_a_HPC2_and_U14 ( .A(Fresh[116]), .B(cell_1830_and_in[0]), 
        .Z(cell_1830_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1830_a_HPC2_and_U13 ( .A(Fresh[116]), .B(cell_1830_and_in[1]), 
        .Z(cell_1830_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1830_a_HPC2_and_U12 ( .A1(cell_1830_a_HPC2_and_a_reg[1]), .A2(
        cell_1830_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1830_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1830_a_HPC2_and_U11 ( .A1(cell_1830_a_HPC2_and_a_reg[0]), .A2(
        cell_1830_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1830_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1830_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1830_a_HPC2_and_n9), 
        .ZN(cell_1830_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1830_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1830_a_HPC2_and_n9), 
        .ZN(cell_1830_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1830_a_HPC2_and_U8 ( .A(Fresh[116]), .ZN(cell_1830_a_HPC2_and_n9) );
  AND2_X1 cell_1830_a_HPC2_and_U7 ( .A1(cell_1830_and_in[1]), .A2(n412), .ZN(
        cell_1830_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1830_a_HPC2_and_U6 ( .A1(cell_1830_and_in[0]), .A2(n395), .ZN(
        cell_1830_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1830_a_HPC2_and_U5 ( .A(cell_1830_a_HPC2_and_n8), .B(
        cell_1830_a_HPC2_and_z_1__1_), .ZN(cell_1830_and_out[1]) );
  XNOR2_X1 cell_1830_a_HPC2_and_U4 ( .A(
        cell_1830_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1830_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1830_a_HPC2_and_n8) );
  XNOR2_X1 cell_1830_a_HPC2_and_U3 ( .A(cell_1830_a_HPC2_and_n7), .B(
        cell_1830_a_HPC2_and_z_0__0_), .ZN(cell_1830_and_out[0]) );
  XNOR2_X1 cell_1830_a_HPC2_and_U2 ( .A(
        cell_1830_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1830_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1830_a_HPC2_and_n7) );
  DFF_X1 cell_1830_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1830_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1830_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1830_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1830_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1830_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1830_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1830_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1830_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1830_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1831_U4 ( .A(n383), .B(cell_1831_and_out[1]), .Z(signal_3537)
         );
  XOR2_X1 cell_1831_U3 ( .A(n382), .B(cell_1831_and_out[0]), .Z(signal_2099)
         );
  XOR2_X1 cell_1831_U2 ( .A(n383), .B(signal_3426), .Z(cell_1831_and_in[1]) );
  XOR2_X1 cell_1831_U1 ( .A(n382), .B(signal_2012), .Z(cell_1831_and_in[0]) );
  XOR2_X1 cell_1831_a_HPC2_and_U14 ( .A(Fresh[117]), .B(cell_1831_and_in[0]), 
        .Z(cell_1831_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1831_a_HPC2_and_U13 ( .A(Fresh[117]), .B(cell_1831_and_in[1]), 
        .Z(cell_1831_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1831_a_HPC2_and_U12 ( .A1(cell_1831_a_HPC2_and_a_reg[1]), .A2(
        cell_1831_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1831_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1831_a_HPC2_and_U11 ( .A1(cell_1831_a_HPC2_and_a_reg[0]), .A2(
        cell_1831_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1831_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1831_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1831_a_HPC2_and_n9), 
        .ZN(cell_1831_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1831_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1831_a_HPC2_and_n9), 
        .ZN(cell_1831_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1831_a_HPC2_and_U8 ( .A(Fresh[117]), .ZN(cell_1831_a_HPC2_and_n9) );
  AND2_X1 cell_1831_a_HPC2_and_U7 ( .A1(cell_1831_and_in[1]), .A2(n420), .ZN(
        cell_1831_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1831_a_HPC2_and_U6 ( .A1(cell_1831_and_in[0]), .A2(n403), .ZN(
        cell_1831_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1831_a_HPC2_and_U5 ( .A(cell_1831_a_HPC2_and_n8), .B(
        cell_1831_a_HPC2_and_z_1__1_), .ZN(cell_1831_and_out[1]) );
  XNOR2_X1 cell_1831_a_HPC2_and_U4 ( .A(
        cell_1831_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1831_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1831_a_HPC2_and_n8) );
  XNOR2_X1 cell_1831_a_HPC2_and_U3 ( .A(cell_1831_a_HPC2_and_n7), .B(
        cell_1831_a_HPC2_and_z_0__0_), .ZN(cell_1831_and_out[0]) );
  XNOR2_X1 cell_1831_a_HPC2_and_U2 ( .A(
        cell_1831_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1831_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1831_a_HPC2_and_n7) );
  DFF_X1 cell_1831_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1831_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1831_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1831_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1831_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1831_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1831_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1831_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1831_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1831_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1832_U4 ( .A(n386), .B(cell_1832_and_out[1]), .Z(signal_3538)
         );
  XOR2_X1 cell_1832_U3 ( .A(n384), .B(cell_1832_and_out[0]), .Z(signal_2100)
         );
  XOR2_X1 cell_1832_U2 ( .A(n386), .B(n361), .Z(cell_1832_and_in[1]) );
  XOR2_X1 cell_1832_U1 ( .A(n384), .B(n359), .Z(cell_1832_and_in[0]) );
  XOR2_X1 cell_1832_a_HPC2_and_U14 ( .A(Fresh[118]), .B(cell_1832_and_in[0]), 
        .Z(cell_1832_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1832_a_HPC2_and_U13 ( .A(Fresh[118]), .B(cell_1832_and_in[1]), 
        .Z(cell_1832_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1832_a_HPC2_and_U12 ( .A1(cell_1832_a_HPC2_and_a_reg[1]), .A2(
        cell_1832_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1832_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1832_a_HPC2_and_U11 ( .A1(cell_1832_a_HPC2_and_a_reg[0]), .A2(
        cell_1832_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1832_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1832_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1832_a_HPC2_and_n9), 
        .ZN(cell_1832_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1832_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1832_a_HPC2_and_n9), 
        .ZN(cell_1832_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1832_a_HPC2_and_U8 ( .A(Fresh[118]), .ZN(cell_1832_a_HPC2_and_n9) );
  AND2_X1 cell_1832_a_HPC2_and_U7 ( .A1(cell_1832_and_in[1]), .A2(n420), .ZN(
        cell_1832_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1832_a_HPC2_and_U6 ( .A1(cell_1832_and_in[0]), .A2(n403), .ZN(
        cell_1832_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1832_a_HPC2_and_U5 ( .A(cell_1832_a_HPC2_and_n8), .B(
        cell_1832_a_HPC2_and_z_1__1_), .ZN(cell_1832_and_out[1]) );
  XNOR2_X1 cell_1832_a_HPC2_and_U4 ( .A(
        cell_1832_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1832_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1832_a_HPC2_and_n8) );
  XNOR2_X1 cell_1832_a_HPC2_and_U3 ( .A(cell_1832_a_HPC2_and_n7), .B(
        cell_1832_a_HPC2_and_z_0__0_), .ZN(cell_1832_and_out[0]) );
  XNOR2_X1 cell_1832_a_HPC2_and_U2 ( .A(
        cell_1832_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1832_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1832_a_HPC2_and_n7) );
  DFF_X1 cell_1832_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1832_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1832_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1832_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1832_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1832_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1832_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1832_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1832_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1832_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1833_U4 ( .A(n381), .B(cell_1833_and_out[1]), .Z(signal_3539)
         );
  XOR2_X1 cell_1833_U3 ( .A(n380), .B(cell_1833_and_out[0]), .Z(signal_2101)
         );
  XOR2_X1 cell_1833_U2 ( .A(n381), .B(n365), .Z(cell_1833_and_in[1]) );
  XOR2_X1 cell_1833_U1 ( .A(n380), .B(n363), .Z(cell_1833_and_in[0]) );
  XOR2_X1 cell_1833_a_HPC2_and_U14 ( .A(Fresh[119]), .B(cell_1833_and_in[0]), 
        .Z(cell_1833_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1833_a_HPC2_and_U13 ( .A(Fresh[119]), .B(cell_1833_and_in[1]), 
        .Z(cell_1833_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1833_a_HPC2_and_U12 ( .A1(cell_1833_a_HPC2_and_a_reg[1]), .A2(
        cell_1833_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1833_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1833_a_HPC2_and_U11 ( .A1(cell_1833_a_HPC2_and_a_reg[0]), .A2(
        cell_1833_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1833_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1833_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1833_a_HPC2_and_n9), 
        .ZN(cell_1833_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1833_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1833_a_HPC2_and_n9), 
        .ZN(cell_1833_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1833_a_HPC2_and_U8 ( .A(Fresh[119]), .ZN(cell_1833_a_HPC2_and_n9) );
  AND2_X1 cell_1833_a_HPC2_and_U7 ( .A1(cell_1833_and_in[1]), .A2(n420), .ZN(
        cell_1833_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1833_a_HPC2_and_U6 ( .A1(cell_1833_and_in[0]), .A2(n403), .ZN(
        cell_1833_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1833_a_HPC2_and_U5 ( .A(cell_1833_a_HPC2_and_n8), .B(
        cell_1833_a_HPC2_and_z_1__1_), .ZN(cell_1833_and_out[1]) );
  XNOR2_X1 cell_1833_a_HPC2_and_U4 ( .A(
        cell_1833_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1833_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1833_a_HPC2_and_n8) );
  XNOR2_X1 cell_1833_a_HPC2_and_U3 ( .A(cell_1833_a_HPC2_and_n7), .B(
        cell_1833_a_HPC2_and_z_0__0_), .ZN(cell_1833_and_out[0]) );
  XNOR2_X1 cell_1833_a_HPC2_and_U2 ( .A(
        cell_1833_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1833_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1833_a_HPC2_and_n7) );
  DFF_X1 cell_1833_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1833_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1833_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1833_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1833_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1833_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1833_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1833_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1833_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1833_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1834_U4 ( .A(n375), .B(cell_1834_and_out[1]), .Z(signal_3540)
         );
  XOR2_X1 cell_1834_U3 ( .A(n373), .B(cell_1834_and_out[0]), .Z(signal_2102)
         );
  XOR2_X1 cell_1834_U2 ( .A(n375), .B(n371), .Z(cell_1834_and_in[1]) );
  XOR2_X1 cell_1834_U1 ( .A(n373), .B(n369), .Z(cell_1834_and_in[0]) );
  XOR2_X1 cell_1834_a_HPC2_and_U14 ( .A(Fresh[120]), .B(cell_1834_and_in[0]), 
        .Z(cell_1834_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1834_a_HPC2_and_U13 ( .A(Fresh[120]), .B(cell_1834_and_in[1]), 
        .Z(cell_1834_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1834_a_HPC2_and_U12 ( .A1(cell_1834_a_HPC2_and_a_reg[1]), .A2(
        cell_1834_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1834_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1834_a_HPC2_and_U11 ( .A1(cell_1834_a_HPC2_and_a_reg[0]), .A2(
        cell_1834_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1834_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1834_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1834_a_HPC2_and_n9), 
        .ZN(cell_1834_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1834_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1834_a_HPC2_and_n9), 
        .ZN(cell_1834_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1834_a_HPC2_and_U8 ( .A(Fresh[120]), .ZN(cell_1834_a_HPC2_and_n9) );
  AND2_X1 cell_1834_a_HPC2_and_U7 ( .A1(cell_1834_and_in[1]), .A2(n420), .ZN(
        cell_1834_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1834_a_HPC2_and_U6 ( .A1(cell_1834_and_in[0]), .A2(n403), .ZN(
        cell_1834_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1834_a_HPC2_and_U5 ( .A(cell_1834_a_HPC2_and_n8), .B(
        cell_1834_a_HPC2_and_z_1__1_), .ZN(cell_1834_and_out[1]) );
  XNOR2_X1 cell_1834_a_HPC2_and_U4 ( .A(
        cell_1834_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1834_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1834_a_HPC2_and_n8) );
  XNOR2_X1 cell_1834_a_HPC2_and_U3 ( .A(cell_1834_a_HPC2_and_n7), .B(
        cell_1834_a_HPC2_and_z_0__0_), .ZN(cell_1834_and_out[0]) );
  XNOR2_X1 cell_1834_a_HPC2_and_U2 ( .A(
        cell_1834_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1834_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1834_a_HPC2_and_n7) );
  DFF_X1 cell_1834_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1834_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1834_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1834_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1834_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1834_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1834_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1834_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1834_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1834_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1835_U4 ( .A(n367), .B(cell_1835_and_out[1]), .Z(signal_3541)
         );
  XOR2_X1 cell_1835_U3 ( .A(n366), .B(cell_1835_and_out[0]), .Z(signal_2103)
         );
  XOR2_X1 cell_1835_U2 ( .A(n367), .B(1'b0), .Z(cell_1835_and_in[1]) );
  XOR2_X1 cell_1835_U1 ( .A(n366), .B(1'b0), .Z(cell_1835_and_in[0]) );
  XOR2_X1 cell_1835_a_HPC2_and_U14 ( .A(Fresh[121]), .B(cell_1835_and_in[0]), 
        .Z(cell_1835_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1835_a_HPC2_and_U13 ( .A(Fresh[121]), .B(cell_1835_and_in[1]), 
        .Z(cell_1835_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1835_a_HPC2_and_U12 ( .A1(cell_1835_a_HPC2_and_a_reg[1]), .A2(
        cell_1835_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1835_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1835_a_HPC2_and_U11 ( .A1(cell_1835_a_HPC2_and_a_reg[0]), .A2(
        cell_1835_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1835_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1835_a_HPC2_and_U10 ( .A1(n417), .A2(cell_1835_a_HPC2_and_n9), 
        .ZN(cell_1835_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1835_a_HPC2_and_U9 ( .A1(n400), .A2(cell_1835_a_HPC2_and_n9), 
        .ZN(cell_1835_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1835_a_HPC2_and_U8 ( .A(Fresh[121]), .ZN(cell_1835_a_HPC2_and_n9) );
  AND2_X1 cell_1835_a_HPC2_and_U7 ( .A1(cell_1835_and_in[1]), .A2(n417), .ZN(
        cell_1835_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1835_a_HPC2_and_U6 ( .A1(cell_1835_and_in[0]), .A2(n400), .ZN(
        cell_1835_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1835_a_HPC2_and_U5 ( .A(cell_1835_a_HPC2_and_n8), .B(
        cell_1835_a_HPC2_and_z_1__1_), .ZN(cell_1835_and_out[1]) );
  XNOR2_X1 cell_1835_a_HPC2_and_U4 ( .A(
        cell_1835_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1835_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1835_a_HPC2_and_n8) );
  XNOR2_X1 cell_1835_a_HPC2_and_U3 ( .A(cell_1835_a_HPC2_and_n7), .B(
        cell_1835_a_HPC2_and_z_0__0_), .ZN(cell_1835_and_out[0]) );
  XNOR2_X1 cell_1835_a_HPC2_and_U2 ( .A(
        cell_1835_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1835_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1835_a_HPC2_and_n7) );
  DFF_X1 cell_1835_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1835_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1835_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n400), .CK(clk), 
        .Q(cell_1835_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1835_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1835_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n417), .CK(clk), 
        .Q(cell_1835_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1835_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1835_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1835_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1836_U4 ( .A(n371), .B(cell_1836_and_out[1]), .Z(signal_3542)
         );
  XOR2_X1 cell_1836_U3 ( .A(n369), .B(cell_1836_and_out[0]), .Z(signal_2104)
         );
  XOR2_X1 cell_1836_U2 ( .A(n371), .B(signal_3258), .Z(cell_1836_and_in[1]) );
  XOR2_X1 cell_1836_U1 ( .A(n369), .B(signal_1984), .Z(cell_1836_and_in[0]) );
  XOR2_X1 cell_1836_a_HPC2_and_U14 ( .A(Fresh[122]), .B(cell_1836_and_in[0]), 
        .Z(cell_1836_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1836_a_HPC2_and_U13 ( .A(Fresh[122]), .B(cell_1836_and_in[1]), 
        .Z(cell_1836_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1836_a_HPC2_and_U12 ( .A1(cell_1836_a_HPC2_and_a_reg[1]), .A2(
        cell_1836_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1836_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1836_a_HPC2_and_U11 ( .A1(cell_1836_a_HPC2_and_a_reg[0]), .A2(
        cell_1836_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1836_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1836_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1836_a_HPC2_and_n9), 
        .ZN(cell_1836_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1836_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1836_a_HPC2_and_n9), 
        .ZN(cell_1836_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1836_a_HPC2_and_U8 ( .A(Fresh[122]), .ZN(cell_1836_a_HPC2_and_n9) );
  AND2_X1 cell_1836_a_HPC2_and_U7 ( .A1(cell_1836_and_in[1]), .A2(n420), .ZN(
        cell_1836_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1836_a_HPC2_and_U6 ( .A1(cell_1836_and_in[0]), .A2(n403), .ZN(
        cell_1836_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1836_a_HPC2_and_U5 ( .A(cell_1836_a_HPC2_and_n8), .B(
        cell_1836_a_HPC2_and_z_1__1_), .ZN(cell_1836_and_out[1]) );
  XNOR2_X1 cell_1836_a_HPC2_and_U4 ( .A(
        cell_1836_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1836_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1836_a_HPC2_and_n8) );
  XNOR2_X1 cell_1836_a_HPC2_and_U3 ( .A(cell_1836_a_HPC2_and_n7), .B(
        cell_1836_a_HPC2_and_z_0__0_), .ZN(cell_1836_and_out[0]) );
  XNOR2_X1 cell_1836_a_HPC2_and_U2 ( .A(
        cell_1836_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1836_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1836_a_HPC2_and_n7) );
  DFF_X1 cell_1836_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1836_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1836_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1836_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1836_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1836_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1836_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1836_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1836_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1836_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1837_U4 ( .A(n379), .B(cell_1837_and_out[1]), .Z(signal_3543)
         );
  XOR2_X1 cell_1837_U3 ( .A(n377), .B(cell_1837_and_out[0]), .Z(signal_2105)
         );
  XOR2_X1 cell_1837_U2 ( .A(n379), .B(n375), .Z(cell_1837_and_in[1]) );
  XOR2_X1 cell_1837_U1 ( .A(n377), .B(n373), .Z(cell_1837_and_in[0]) );
  XOR2_X1 cell_1837_a_HPC2_and_U14 ( .A(Fresh[123]), .B(cell_1837_and_in[0]), 
        .Z(cell_1837_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1837_a_HPC2_and_U13 ( .A(Fresh[123]), .B(cell_1837_and_in[1]), 
        .Z(cell_1837_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1837_a_HPC2_and_U12 ( .A1(cell_1837_a_HPC2_and_a_reg[1]), .A2(
        cell_1837_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1837_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1837_a_HPC2_and_U11 ( .A1(cell_1837_a_HPC2_and_a_reg[0]), .A2(
        cell_1837_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1837_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1837_a_HPC2_and_U10 ( .A1(n420), .A2(cell_1837_a_HPC2_and_n9), 
        .ZN(cell_1837_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1837_a_HPC2_and_U9 ( .A1(n403), .A2(cell_1837_a_HPC2_and_n9), 
        .ZN(cell_1837_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1837_a_HPC2_and_U8 ( .A(Fresh[123]), .ZN(cell_1837_a_HPC2_and_n9) );
  AND2_X1 cell_1837_a_HPC2_and_U7 ( .A1(cell_1837_and_in[1]), .A2(n420), .ZN(
        cell_1837_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1837_a_HPC2_and_U6 ( .A1(cell_1837_and_in[0]), .A2(n403), .ZN(
        cell_1837_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1837_a_HPC2_and_U5 ( .A(cell_1837_a_HPC2_and_n8), .B(
        cell_1837_a_HPC2_and_z_1__1_), .ZN(cell_1837_and_out[1]) );
  XNOR2_X1 cell_1837_a_HPC2_and_U4 ( .A(
        cell_1837_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1837_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1837_a_HPC2_and_n8) );
  XNOR2_X1 cell_1837_a_HPC2_and_U3 ( .A(cell_1837_a_HPC2_and_n7), .B(
        cell_1837_a_HPC2_and_z_0__0_), .ZN(cell_1837_and_out[0]) );
  XNOR2_X1 cell_1837_a_HPC2_and_U2 ( .A(
        cell_1837_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1837_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1837_a_HPC2_and_n7) );
  DFF_X1 cell_1837_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1837_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1837_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n403), .CK(clk), 
        .Q(cell_1837_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1837_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1837_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n420), .CK(clk), 
        .Q(cell_1837_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1837_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1837_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1837_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1838_U4 ( .A(n361), .B(cell_1838_and_out[1]), .Z(signal_3544)
         );
  XOR2_X1 cell_1838_U3 ( .A(n359), .B(cell_1838_and_out[0]), .Z(signal_2106)
         );
  XOR2_X1 cell_1838_U2 ( .A(n361), .B(signal_3426), .Z(cell_1838_and_in[1]) );
  XOR2_X1 cell_1838_U1 ( .A(n359), .B(signal_2012), .Z(cell_1838_and_in[0]) );
  XOR2_X1 cell_1838_a_HPC2_and_U14 ( .A(Fresh[124]), .B(cell_1838_and_in[0]), 
        .Z(cell_1838_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1838_a_HPC2_and_U13 ( .A(Fresh[124]), .B(cell_1838_and_in[1]), 
        .Z(cell_1838_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1838_a_HPC2_and_U12 ( .A1(cell_1838_a_HPC2_and_a_reg[1]), .A2(
        cell_1838_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1838_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1838_a_HPC2_and_U11 ( .A1(cell_1838_a_HPC2_and_a_reg[0]), .A2(
        cell_1838_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1838_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1838_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1838_a_HPC2_and_n9), 
        .ZN(cell_1838_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1838_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1838_a_HPC2_and_n9), 
        .ZN(cell_1838_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1838_a_HPC2_and_U8 ( .A(Fresh[124]), .ZN(cell_1838_a_HPC2_and_n9) );
  AND2_X1 cell_1838_a_HPC2_and_U7 ( .A1(cell_1838_and_in[1]), .A2(n421), .ZN(
        cell_1838_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1838_a_HPC2_and_U6 ( .A1(cell_1838_and_in[0]), .A2(n404), .ZN(
        cell_1838_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1838_a_HPC2_and_U5 ( .A(cell_1838_a_HPC2_and_n8), .B(
        cell_1838_a_HPC2_and_z_1__1_), .ZN(cell_1838_and_out[1]) );
  XNOR2_X1 cell_1838_a_HPC2_and_U4 ( .A(
        cell_1838_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1838_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1838_a_HPC2_and_n8) );
  XNOR2_X1 cell_1838_a_HPC2_and_U3 ( .A(cell_1838_a_HPC2_and_n7), .B(
        cell_1838_a_HPC2_and_z_0__0_), .ZN(cell_1838_and_out[0]) );
  XNOR2_X1 cell_1838_a_HPC2_and_U2 ( .A(
        cell_1838_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1838_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1838_a_HPC2_and_n7) );
  DFF_X1 cell_1838_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1838_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1838_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1838_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1838_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1838_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1838_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1838_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1838_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1838_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1839_U4 ( .A(n357), .B(cell_1839_and_out[1]), .Z(signal_3545)
         );
  XOR2_X1 cell_1839_U3 ( .A(n356), .B(cell_1839_and_out[0]), .Z(signal_2107)
         );
  XOR2_X1 cell_1839_U2 ( .A(n357), .B(n381), .Z(cell_1839_and_in[1]) );
  XOR2_X1 cell_1839_U1 ( .A(n356), .B(n380), .Z(cell_1839_and_in[0]) );
  XOR2_X1 cell_1839_a_HPC2_and_U14 ( .A(Fresh[125]), .B(cell_1839_and_in[0]), 
        .Z(cell_1839_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1839_a_HPC2_and_U13 ( .A(Fresh[125]), .B(cell_1839_and_in[1]), 
        .Z(cell_1839_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1839_a_HPC2_and_U12 ( .A1(cell_1839_a_HPC2_and_a_reg[1]), .A2(
        cell_1839_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1839_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1839_a_HPC2_and_U11 ( .A1(cell_1839_a_HPC2_and_a_reg[0]), .A2(
        cell_1839_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1839_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1839_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1839_a_HPC2_and_n9), 
        .ZN(cell_1839_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1839_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1839_a_HPC2_and_n9), 
        .ZN(cell_1839_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1839_a_HPC2_and_U8 ( .A(Fresh[125]), .ZN(cell_1839_a_HPC2_and_n9) );
  AND2_X1 cell_1839_a_HPC2_and_U7 ( .A1(cell_1839_and_in[1]), .A2(n421), .ZN(
        cell_1839_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1839_a_HPC2_and_U6 ( .A1(cell_1839_and_in[0]), .A2(n404), .ZN(
        cell_1839_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1839_a_HPC2_and_U5 ( .A(cell_1839_a_HPC2_and_n8), .B(
        cell_1839_a_HPC2_and_z_1__1_), .ZN(cell_1839_and_out[1]) );
  XNOR2_X1 cell_1839_a_HPC2_and_U4 ( .A(
        cell_1839_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1839_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1839_a_HPC2_and_n8) );
  XNOR2_X1 cell_1839_a_HPC2_and_U3 ( .A(cell_1839_a_HPC2_and_n7), .B(
        cell_1839_a_HPC2_and_z_0__0_), .ZN(cell_1839_and_out[0]) );
  XNOR2_X1 cell_1839_a_HPC2_and_U2 ( .A(
        cell_1839_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1839_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1839_a_HPC2_and_n7) );
  DFF_X1 cell_1839_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1839_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1839_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1839_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1839_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1839_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1839_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1839_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1839_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1839_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1840_U4 ( .A(n381), .B(cell_1840_and_out[1]), .Z(signal_3546)
         );
  XOR2_X1 cell_1840_U3 ( .A(n380), .B(cell_1840_and_out[0]), .Z(signal_2108)
         );
  XOR2_X1 cell_1840_U2 ( .A(n381), .B(n375), .Z(cell_1840_and_in[1]) );
  XOR2_X1 cell_1840_U1 ( .A(n380), .B(n373), .Z(cell_1840_and_in[0]) );
  XOR2_X1 cell_1840_a_HPC2_and_U14 ( .A(Fresh[126]), .B(cell_1840_and_in[0]), 
        .Z(cell_1840_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1840_a_HPC2_and_U13 ( .A(Fresh[126]), .B(cell_1840_and_in[1]), 
        .Z(cell_1840_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1840_a_HPC2_and_U12 ( .A1(cell_1840_a_HPC2_and_a_reg[1]), .A2(
        cell_1840_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1840_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1840_a_HPC2_and_U11 ( .A1(cell_1840_a_HPC2_and_a_reg[0]), .A2(
        cell_1840_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1840_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1840_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1840_a_HPC2_and_n9), 
        .ZN(cell_1840_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1840_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1840_a_HPC2_and_n9), 
        .ZN(cell_1840_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1840_a_HPC2_and_U8 ( .A(Fresh[126]), .ZN(cell_1840_a_HPC2_and_n9) );
  AND2_X1 cell_1840_a_HPC2_and_U7 ( .A1(cell_1840_and_in[1]), .A2(n421), .ZN(
        cell_1840_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1840_a_HPC2_and_U6 ( .A1(cell_1840_and_in[0]), .A2(n404), .ZN(
        cell_1840_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1840_a_HPC2_and_U5 ( .A(cell_1840_a_HPC2_and_n8), .B(
        cell_1840_a_HPC2_and_z_1__1_), .ZN(cell_1840_and_out[1]) );
  XNOR2_X1 cell_1840_a_HPC2_and_U4 ( .A(
        cell_1840_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1840_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1840_a_HPC2_and_n8) );
  XNOR2_X1 cell_1840_a_HPC2_and_U3 ( .A(cell_1840_a_HPC2_and_n7), .B(
        cell_1840_a_HPC2_and_z_0__0_), .ZN(cell_1840_and_out[0]) );
  XNOR2_X1 cell_1840_a_HPC2_and_U2 ( .A(
        cell_1840_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1840_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1840_a_HPC2_and_n7) );
  DFF_X1 cell_1840_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1840_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1840_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1840_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1840_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1840_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1840_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1840_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1840_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1840_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1841_U4 ( .A(n386), .B(cell_1841_and_out[1]), .Z(signal_3547)
         );
  XOR2_X1 cell_1841_U3 ( .A(n384), .B(cell_1841_and_out[0]), .Z(signal_2109)
         );
  XOR2_X1 cell_1841_U2 ( .A(n386), .B(n357), .Z(cell_1841_and_in[1]) );
  XOR2_X1 cell_1841_U1 ( .A(n384), .B(n356), .Z(cell_1841_and_in[0]) );
  XOR2_X1 cell_1841_a_HPC2_and_U14 ( .A(Fresh[127]), .B(cell_1841_and_in[0]), 
        .Z(cell_1841_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1841_a_HPC2_and_U13 ( .A(Fresh[127]), .B(cell_1841_and_in[1]), 
        .Z(cell_1841_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1841_a_HPC2_and_U12 ( .A1(cell_1841_a_HPC2_and_a_reg[1]), .A2(
        cell_1841_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1841_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1841_a_HPC2_and_U11 ( .A1(cell_1841_a_HPC2_and_a_reg[0]), .A2(
        cell_1841_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1841_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1841_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1841_a_HPC2_and_n9), 
        .ZN(cell_1841_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1841_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1841_a_HPC2_and_n9), 
        .ZN(cell_1841_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1841_a_HPC2_and_U8 ( .A(Fresh[127]), .ZN(cell_1841_a_HPC2_and_n9) );
  AND2_X1 cell_1841_a_HPC2_and_U7 ( .A1(cell_1841_and_in[1]), .A2(n421), .ZN(
        cell_1841_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1841_a_HPC2_and_U6 ( .A1(cell_1841_and_in[0]), .A2(n404), .ZN(
        cell_1841_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1841_a_HPC2_and_U5 ( .A(cell_1841_a_HPC2_and_n8), .B(
        cell_1841_a_HPC2_and_z_1__1_), .ZN(cell_1841_and_out[1]) );
  XNOR2_X1 cell_1841_a_HPC2_and_U4 ( .A(
        cell_1841_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1841_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1841_a_HPC2_and_n8) );
  XNOR2_X1 cell_1841_a_HPC2_and_U3 ( .A(cell_1841_a_HPC2_and_n7), .B(
        cell_1841_a_HPC2_and_z_0__0_), .ZN(cell_1841_and_out[0]) );
  XNOR2_X1 cell_1841_a_HPC2_and_U2 ( .A(
        cell_1841_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1841_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1841_a_HPC2_and_n7) );
  DFF_X1 cell_1841_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1841_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1841_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1841_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1841_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1841_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1841_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1841_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1841_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1841_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1842_U4 ( .A(n370), .B(cell_1842_and_out[1]), .Z(signal_3548)
         );
  XOR2_X1 cell_1842_U3 ( .A(n368), .B(cell_1842_and_out[0]), .Z(signal_2110)
         );
  XOR2_X1 cell_1842_U2 ( .A(n370), .B(signal_3426), .Z(cell_1842_and_in[1]) );
  XOR2_X1 cell_1842_U1 ( .A(n368), .B(signal_2012), .Z(cell_1842_and_in[0]) );
  XOR2_X1 cell_1842_a_HPC2_and_U14 ( .A(Fresh[128]), .B(cell_1842_and_in[0]), 
        .Z(cell_1842_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1842_a_HPC2_and_U13 ( .A(Fresh[128]), .B(cell_1842_and_in[1]), 
        .Z(cell_1842_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1842_a_HPC2_and_U12 ( .A1(cell_1842_a_HPC2_and_a_reg[1]), .A2(
        cell_1842_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1842_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1842_a_HPC2_and_U11 ( .A1(cell_1842_a_HPC2_and_a_reg[0]), .A2(
        cell_1842_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1842_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1842_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1842_a_HPC2_and_n9), 
        .ZN(cell_1842_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1842_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1842_a_HPC2_and_n9), 
        .ZN(cell_1842_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1842_a_HPC2_and_U8 ( .A(Fresh[128]), .ZN(cell_1842_a_HPC2_and_n9) );
  AND2_X1 cell_1842_a_HPC2_and_U7 ( .A1(cell_1842_and_in[1]), .A2(n421), .ZN(
        cell_1842_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1842_a_HPC2_and_U6 ( .A1(cell_1842_and_in[0]), .A2(n404), .ZN(
        cell_1842_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1842_a_HPC2_and_U5 ( .A(cell_1842_a_HPC2_and_n8), .B(
        cell_1842_a_HPC2_and_z_1__1_), .ZN(cell_1842_and_out[1]) );
  XNOR2_X1 cell_1842_a_HPC2_and_U4 ( .A(
        cell_1842_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1842_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1842_a_HPC2_and_n8) );
  XNOR2_X1 cell_1842_a_HPC2_and_U3 ( .A(cell_1842_a_HPC2_and_n7), .B(
        cell_1842_a_HPC2_and_z_0__0_), .ZN(cell_1842_and_out[0]) );
  XNOR2_X1 cell_1842_a_HPC2_and_U2 ( .A(
        cell_1842_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1842_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1842_a_HPC2_and_n7) );
  DFF_X1 cell_1842_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1842_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1842_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1842_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1842_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1842_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1842_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1842_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1842_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1842_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1843_U4 ( .A(n364), .B(cell_1843_and_out[1]), .Z(signal_3549)
         );
  XOR2_X1 cell_1843_U3 ( .A(n362), .B(cell_1843_and_out[0]), .Z(signal_2111)
         );
  XOR2_X1 cell_1843_U2 ( .A(n364), .B(n375), .Z(cell_1843_and_in[1]) );
  XOR2_X1 cell_1843_U1 ( .A(n362), .B(n373), .Z(cell_1843_and_in[0]) );
  XOR2_X1 cell_1843_a_HPC2_and_U14 ( .A(Fresh[129]), .B(cell_1843_and_in[0]), 
        .Z(cell_1843_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1843_a_HPC2_and_U13 ( .A(Fresh[129]), .B(cell_1843_and_in[1]), 
        .Z(cell_1843_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1843_a_HPC2_and_U12 ( .A1(cell_1843_a_HPC2_and_a_reg[1]), .A2(
        cell_1843_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1843_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1843_a_HPC2_and_U11 ( .A1(cell_1843_a_HPC2_and_a_reg[0]), .A2(
        cell_1843_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1843_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1843_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1843_a_HPC2_and_n9), 
        .ZN(cell_1843_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1843_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1843_a_HPC2_and_n9), 
        .ZN(cell_1843_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1843_a_HPC2_and_U8 ( .A(Fresh[129]), .ZN(cell_1843_a_HPC2_and_n9) );
  AND2_X1 cell_1843_a_HPC2_and_U7 ( .A1(cell_1843_and_in[1]), .A2(n421), .ZN(
        cell_1843_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1843_a_HPC2_and_U6 ( .A1(cell_1843_and_in[0]), .A2(n404), .ZN(
        cell_1843_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1843_a_HPC2_and_U5 ( .A(cell_1843_a_HPC2_and_n8), .B(
        cell_1843_a_HPC2_and_z_1__1_), .ZN(cell_1843_and_out[1]) );
  XNOR2_X1 cell_1843_a_HPC2_and_U4 ( .A(
        cell_1843_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1843_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1843_a_HPC2_and_n8) );
  XNOR2_X1 cell_1843_a_HPC2_and_U3 ( .A(cell_1843_a_HPC2_and_n7), .B(
        cell_1843_a_HPC2_and_z_0__0_), .ZN(cell_1843_and_out[0]) );
  XNOR2_X1 cell_1843_a_HPC2_and_U2 ( .A(
        cell_1843_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1843_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1843_a_HPC2_and_n7) );
  DFF_X1 cell_1843_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1843_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1843_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1843_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1843_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1843_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1843_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1843_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1843_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1843_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1844_U4 ( .A(signal_3426), .B(cell_1844_and_out[1]), .Z(
        signal_3550) );
  XOR2_X1 cell_1844_U3 ( .A(signal_2012), .B(cell_1844_and_out[0]), .Z(
        signal_2112) );
  XOR2_X1 cell_1844_U2 ( .A(signal_3426), .B(n379), .Z(cell_1844_and_in[1]) );
  XOR2_X1 cell_1844_U1 ( .A(signal_2012), .B(n377), .Z(cell_1844_and_in[0]) );
  XOR2_X1 cell_1844_a_HPC2_and_U14 ( .A(Fresh[130]), .B(cell_1844_and_in[0]), 
        .Z(cell_1844_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1844_a_HPC2_and_U13 ( .A(Fresh[130]), .B(cell_1844_and_in[1]), 
        .Z(cell_1844_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1844_a_HPC2_and_U12 ( .A1(cell_1844_a_HPC2_and_a_reg[1]), .A2(
        cell_1844_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1844_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1844_a_HPC2_and_U11 ( .A1(cell_1844_a_HPC2_and_a_reg[0]), .A2(
        cell_1844_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1844_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1844_a_HPC2_and_U10 ( .A1(n421), .A2(cell_1844_a_HPC2_and_n9), 
        .ZN(cell_1844_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1844_a_HPC2_and_U9 ( .A1(n404), .A2(cell_1844_a_HPC2_and_n9), 
        .ZN(cell_1844_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1844_a_HPC2_and_U8 ( .A(Fresh[130]), .ZN(cell_1844_a_HPC2_and_n9) );
  AND2_X1 cell_1844_a_HPC2_and_U7 ( .A1(cell_1844_and_in[1]), .A2(n421), .ZN(
        cell_1844_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1844_a_HPC2_and_U6 ( .A1(cell_1844_and_in[0]), .A2(n404), .ZN(
        cell_1844_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1844_a_HPC2_and_U5 ( .A(cell_1844_a_HPC2_and_n8), .B(
        cell_1844_a_HPC2_and_z_1__1_), .ZN(cell_1844_and_out[1]) );
  XNOR2_X1 cell_1844_a_HPC2_and_U4 ( .A(
        cell_1844_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1844_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1844_a_HPC2_and_n8) );
  XNOR2_X1 cell_1844_a_HPC2_and_U3 ( .A(cell_1844_a_HPC2_and_n7), .B(
        cell_1844_a_HPC2_and_z_0__0_), .ZN(cell_1844_and_out[0]) );
  XNOR2_X1 cell_1844_a_HPC2_and_U2 ( .A(
        cell_1844_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1844_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1844_a_HPC2_and_n7) );
  DFF_X1 cell_1844_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1844_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1844_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n404), .CK(clk), 
        .Q(cell_1844_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1844_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1844_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n421), .CK(clk), 
        .Q(cell_1844_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1844_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1844_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1844_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1845_U4 ( .A(n357), .B(cell_1845_and_out[1]), .Z(signal_3551)
         );
  XOR2_X1 cell_1845_U3 ( .A(n356), .B(cell_1845_and_out[0]), .Z(signal_2113)
         );
  XOR2_X1 cell_1845_U2 ( .A(n357), .B(1'b0), .Z(cell_1845_and_in[1]) );
  XOR2_X1 cell_1845_U1 ( .A(n356), .B(1'b0), .Z(cell_1845_and_in[0]) );
  XOR2_X1 cell_1845_a_HPC2_and_U14 ( .A(Fresh[131]), .B(cell_1845_and_in[0]), 
        .Z(cell_1845_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1845_a_HPC2_and_U13 ( .A(Fresh[131]), .B(cell_1845_and_in[1]), 
        .Z(cell_1845_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1845_a_HPC2_and_U12 ( .A1(cell_1845_a_HPC2_and_a_reg[1]), .A2(
        cell_1845_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1845_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1845_a_HPC2_and_U11 ( .A1(cell_1845_a_HPC2_and_a_reg[0]), .A2(
        cell_1845_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1845_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1845_a_HPC2_and_U10 ( .A1(n416), .A2(cell_1845_a_HPC2_and_n9), 
        .ZN(cell_1845_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1845_a_HPC2_and_U9 ( .A1(n399), .A2(cell_1845_a_HPC2_and_n9), 
        .ZN(cell_1845_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1845_a_HPC2_and_U8 ( .A(Fresh[131]), .ZN(cell_1845_a_HPC2_and_n9) );
  AND2_X1 cell_1845_a_HPC2_and_U7 ( .A1(cell_1845_and_in[1]), .A2(n416), .ZN(
        cell_1845_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1845_a_HPC2_and_U6 ( .A1(cell_1845_and_in[0]), .A2(n399), .ZN(
        cell_1845_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1845_a_HPC2_and_U5 ( .A(cell_1845_a_HPC2_and_n8), .B(
        cell_1845_a_HPC2_and_z_1__1_), .ZN(cell_1845_and_out[1]) );
  XNOR2_X1 cell_1845_a_HPC2_and_U4 ( .A(
        cell_1845_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1845_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1845_a_HPC2_and_n8) );
  XNOR2_X1 cell_1845_a_HPC2_and_U3 ( .A(cell_1845_a_HPC2_and_n7), .B(
        cell_1845_a_HPC2_and_z_0__0_), .ZN(cell_1845_and_out[0]) );
  XNOR2_X1 cell_1845_a_HPC2_and_U2 ( .A(
        cell_1845_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1845_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1845_a_HPC2_and_n7) );
  DFF_X1 cell_1845_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1845_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1845_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n399), .CK(clk), 
        .Q(cell_1845_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1845_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1845_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n416), .CK(clk), 
        .Q(cell_1845_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1845_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1845_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1845_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1846_U4 ( .A(signal_3406), .B(cell_1846_and_out[1]), .Z(
        signal_3552) );
  XOR2_X1 cell_1846_U3 ( .A(signal_1992), .B(cell_1846_and_out[0]), .Z(
        signal_2114) );
  XOR2_X1 cell_1846_U2 ( .A(signal_3406), .B(n367), .Z(cell_1846_and_in[1]) );
  XOR2_X1 cell_1846_U1 ( .A(signal_1992), .B(n366), .Z(cell_1846_and_in[0]) );
  XOR2_X1 cell_1846_a_HPC2_and_U14 ( .A(Fresh[132]), .B(cell_1846_and_in[0]), 
        .Z(cell_1846_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1846_a_HPC2_and_U13 ( .A(Fresh[132]), .B(cell_1846_and_in[1]), 
        .Z(cell_1846_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1846_a_HPC2_and_U12 ( .A1(cell_1846_a_HPC2_and_a_reg[1]), .A2(
        cell_1846_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1846_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1846_a_HPC2_and_U11 ( .A1(cell_1846_a_HPC2_and_a_reg[0]), .A2(
        cell_1846_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1846_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1846_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1846_a_HPC2_and_n9), 
        .ZN(cell_1846_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1846_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1846_a_HPC2_and_n9), 
        .ZN(cell_1846_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1846_a_HPC2_and_U8 ( .A(Fresh[132]), .ZN(cell_1846_a_HPC2_and_n9) );
  AND2_X1 cell_1846_a_HPC2_and_U7 ( .A1(cell_1846_and_in[1]), .A2(n411), .ZN(
        cell_1846_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1846_a_HPC2_and_U6 ( .A1(cell_1846_and_in[0]), .A2(n394), .ZN(
        cell_1846_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1846_a_HPC2_and_U5 ( .A(cell_1846_a_HPC2_and_n8), .B(
        cell_1846_a_HPC2_and_z_1__1_), .ZN(cell_1846_and_out[1]) );
  XNOR2_X1 cell_1846_a_HPC2_and_U4 ( .A(
        cell_1846_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1846_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1846_a_HPC2_and_n8) );
  XNOR2_X1 cell_1846_a_HPC2_and_U3 ( .A(cell_1846_a_HPC2_and_n7), .B(
        cell_1846_a_HPC2_and_z_0__0_), .ZN(cell_1846_and_out[0]) );
  XNOR2_X1 cell_1846_a_HPC2_and_U2 ( .A(
        cell_1846_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1846_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1846_a_HPC2_and_n7) );
  DFF_X1 cell_1846_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1846_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1846_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1846_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1846_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1846_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1846_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1846_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1846_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1846_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1847_U4 ( .A(n360), .B(cell_1847_and_out[1]), .Z(signal_3553)
         );
  XOR2_X1 cell_1847_U3 ( .A(n358), .B(cell_1847_and_out[0]), .Z(signal_2115)
         );
  XOR2_X1 cell_1847_U2 ( .A(n360), .B(n367), .Z(cell_1847_and_in[1]) );
  XOR2_X1 cell_1847_U1 ( .A(n358), .B(n366), .Z(cell_1847_and_in[0]) );
  XOR2_X1 cell_1847_a_HPC2_and_U14 ( .A(Fresh[133]), .B(cell_1847_and_in[0]), 
        .Z(cell_1847_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1847_a_HPC2_and_U13 ( .A(Fresh[133]), .B(cell_1847_and_in[1]), 
        .Z(cell_1847_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1847_a_HPC2_and_U12 ( .A1(cell_1847_a_HPC2_and_a_reg[1]), .A2(
        cell_1847_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1847_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1847_a_HPC2_and_U11 ( .A1(cell_1847_a_HPC2_and_a_reg[0]), .A2(
        cell_1847_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1847_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1847_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1847_a_HPC2_and_n9), 
        .ZN(cell_1847_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1847_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1847_a_HPC2_and_n9), 
        .ZN(cell_1847_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1847_a_HPC2_and_U8 ( .A(Fresh[133]), .ZN(cell_1847_a_HPC2_and_n9) );
  AND2_X1 cell_1847_a_HPC2_and_U7 ( .A1(cell_1847_and_in[1]), .A2(n422), .ZN(
        cell_1847_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1847_a_HPC2_and_U6 ( .A1(cell_1847_and_in[0]), .A2(n405), .ZN(
        cell_1847_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1847_a_HPC2_and_U5 ( .A(cell_1847_a_HPC2_and_n8), .B(
        cell_1847_a_HPC2_and_z_1__1_), .ZN(cell_1847_and_out[1]) );
  XNOR2_X1 cell_1847_a_HPC2_and_U4 ( .A(
        cell_1847_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1847_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1847_a_HPC2_and_n8) );
  XNOR2_X1 cell_1847_a_HPC2_and_U3 ( .A(cell_1847_a_HPC2_and_n7), .B(
        cell_1847_a_HPC2_and_z_0__0_), .ZN(cell_1847_and_out[0]) );
  XNOR2_X1 cell_1847_a_HPC2_and_U2 ( .A(
        cell_1847_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1847_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1847_a_HPC2_and_n7) );
  DFF_X1 cell_1847_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1847_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1847_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1847_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1847_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1847_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1847_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1847_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1847_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1847_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1848_U4 ( .A(signal_3406), .B(cell_1848_and_out[1]), .Z(
        signal_3554) );
  XOR2_X1 cell_1848_U3 ( .A(signal_1992), .B(cell_1848_and_out[0]), .Z(
        signal_2116) );
  XOR2_X1 cell_1848_U2 ( .A(signal_3406), .B(n387), .Z(cell_1848_and_in[1]) );
  XOR2_X1 cell_1848_U1 ( .A(signal_1992), .B(n385), .Z(cell_1848_and_in[0]) );
  XOR2_X1 cell_1848_a_HPC2_and_U14 ( .A(Fresh[134]), .B(cell_1848_and_in[0]), 
        .Z(cell_1848_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1848_a_HPC2_and_U13 ( .A(Fresh[134]), .B(cell_1848_and_in[1]), 
        .Z(cell_1848_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1848_a_HPC2_and_U12 ( .A1(cell_1848_a_HPC2_and_a_reg[1]), .A2(
        cell_1848_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1848_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1848_a_HPC2_and_U11 ( .A1(cell_1848_a_HPC2_and_a_reg[0]), .A2(
        cell_1848_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1848_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1848_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1848_a_HPC2_and_n9), 
        .ZN(cell_1848_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1848_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1848_a_HPC2_and_n9), 
        .ZN(cell_1848_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1848_a_HPC2_and_U8 ( .A(Fresh[134]), .ZN(cell_1848_a_HPC2_and_n9) );
  AND2_X1 cell_1848_a_HPC2_and_U7 ( .A1(cell_1848_and_in[1]), .A2(n411), .ZN(
        cell_1848_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1848_a_HPC2_and_U6 ( .A1(cell_1848_and_in[0]), .A2(n394), .ZN(
        cell_1848_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1848_a_HPC2_and_U5 ( .A(cell_1848_a_HPC2_and_n8), .B(
        cell_1848_a_HPC2_and_z_1__1_), .ZN(cell_1848_and_out[1]) );
  XNOR2_X1 cell_1848_a_HPC2_and_U4 ( .A(
        cell_1848_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1848_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1848_a_HPC2_and_n8) );
  XNOR2_X1 cell_1848_a_HPC2_and_U3 ( .A(cell_1848_a_HPC2_and_n7), .B(
        cell_1848_a_HPC2_and_z_0__0_), .ZN(cell_1848_and_out[0]) );
  XNOR2_X1 cell_1848_a_HPC2_and_U2 ( .A(
        cell_1848_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1848_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1848_a_HPC2_and_n7) );
  DFF_X1 cell_1848_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1848_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1848_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1848_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1848_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1848_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1848_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1848_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1848_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1848_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1849_U4 ( .A(signal_3426), .B(cell_1849_and_out[1]), .Z(
        signal_3555) );
  XOR2_X1 cell_1849_U3 ( .A(signal_2012), .B(cell_1849_and_out[0]), .Z(
        signal_2117) );
  XOR2_X1 cell_1849_U2 ( .A(signal_3426), .B(n371), .Z(cell_1849_and_in[1]) );
  XOR2_X1 cell_1849_U1 ( .A(signal_2012), .B(n369), .Z(cell_1849_and_in[0]) );
  XOR2_X1 cell_1849_a_HPC2_and_U14 ( .A(Fresh[135]), .B(cell_1849_and_in[0]), 
        .Z(cell_1849_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1849_a_HPC2_and_U13 ( .A(Fresh[135]), .B(cell_1849_and_in[1]), 
        .Z(cell_1849_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1849_a_HPC2_and_U12 ( .A1(cell_1849_a_HPC2_and_a_reg[1]), .A2(
        cell_1849_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1849_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1849_a_HPC2_and_U11 ( .A1(cell_1849_a_HPC2_and_a_reg[0]), .A2(
        cell_1849_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1849_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1849_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1849_a_HPC2_and_n9), 
        .ZN(cell_1849_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1849_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1849_a_HPC2_and_n9), 
        .ZN(cell_1849_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1849_a_HPC2_and_U8 ( .A(Fresh[135]), .ZN(cell_1849_a_HPC2_and_n9) );
  AND2_X1 cell_1849_a_HPC2_and_U7 ( .A1(cell_1849_and_in[1]), .A2(n422), .ZN(
        cell_1849_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1849_a_HPC2_and_U6 ( .A1(cell_1849_and_in[0]), .A2(n405), .ZN(
        cell_1849_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1849_a_HPC2_and_U5 ( .A(cell_1849_a_HPC2_and_n8), .B(
        cell_1849_a_HPC2_and_z_1__1_), .ZN(cell_1849_and_out[1]) );
  XNOR2_X1 cell_1849_a_HPC2_and_U4 ( .A(
        cell_1849_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1849_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1849_a_HPC2_and_n8) );
  XNOR2_X1 cell_1849_a_HPC2_and_U3 ( .A(cell_1849_a_HPC2_and_n7), .B(
        cell_1849_a_HPC2_and_z_0__0_), .ZN(cell_1849_and_out[0]) );
  XNOR2_X1 cell_1849_a_HPC2_and_U2 ( .A(
        cell_1849_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1849_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1849_a_HPC2_and_n7) );
  DFF_X1 cell_1849_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1849_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1849_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1849_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1849_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1849_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1849_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1849_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1849_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1849_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1850_U4 ( .A(n357), .B(cell_1850_and_out[1]), .Z(signal_3556)
         );
  XOR2_X1 cell_1850_U3 ( .A(n356), .B(cell_1850_and_out[0]), .Z(signal_2118)
         );
  XOR2_X1 cell_1850_U2 ( .A(n357), .B(n375), .Z(cell_1850_and_in[1]) );
  XOR2_X1 cell_1850_U1 ( .A(n356), .B(n373), .Z(cell_1850_and_in[0]) );
  XOR2_X1 cell_1850_a_HPC2_and_U14 ( .A(Fresh[136]), .B(cell_1850_and_in[0]), 
        .Z(cell_1850_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1850_a_HPC2_and_U13 ( .A(Fresh[136]), .B(cell_1850_and_in[1]), 
        .Z(cell_1850_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1850_a_HPC2_and_U12 ( .A1(cell_1850_a_HPC2_and_a_reg[1]), .A2(
        cell_1850_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1850_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1850_a_HPC2_and_U11 ( .A1(cell_1850_a_HPC2_and_a_reg[0]), .A2(
        cell_1850_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1850_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1850_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1850_a_HPC2_and_n9), 
        .ZN(cell_1850_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1850_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1850_a_HPC2_and_n9), 
        .ZN(cell_1850_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1850_a_HPC2_and_U8 ( .A(Fresh[136]), .ZN(cell_1850_a_HPC2_and_n9) );
  AND2_X1 cell_1850_a_HPC2_and_U7 ( .A1(cell_1850_and_in[1]), .A2(n422), .ZN(
        cell_1850_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1850_a_HPC2_and_U6 ( .A1(cell_1850_and_in[0]), .A2(n405), .ZN(
        cell_1850_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1850_a_HPC2_and_U5 ( .A(cell_1850_a_HPC2_and_n8), .B(
        cell_1850_a_HPC2_and_z_1__1_), .ZN(cell_1850_and_out[1]) );
  XNOR2_X1 cell_1850_a_HPC2_and_U4 ( .A(
        cell_1850_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1850_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1850_a_HPC2_and_n8) );
  XNOR2_X1 cell_1850_a_HPC2_and_U3 ( .A(cell_1850_a_HPC2_and_n7), .B(
        cell_1850_a_HPC2_and_z_0__0_), .ZN(cell_1850_and_out[0]) );
  XNOR2_X1 cell_1850_a_HPC2_and_U2 ( .A(
        cell_1850_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1850_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1850_a_HPC2_and_n7) );
  DFF_X1 cell_1850_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1850_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1850_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1850_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1850_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1850_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1850_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1850_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1850_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1850_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1851_U4 ( .A(n367), .B(cell_1851_and_out[1]), .Z(signal_3557)
         );
  XOR2_X1 cell_1851_U3 ( .A(n366), .B(cell_1851_and_out[0]), .Z(signal_2119)
         );
  XOR2_X1 cell_1851_U2 ( .A(n367), .B(n365), .Z(cell_1851_and_in[1]) );
  XOR2_X1 cell_1851_U1 ( .A(n366), .B(n363), .Z(cell_1851_and_in[0]) );
  XOR2_X1 cell_1851_a_HPC2_and_U14 ( .A(Fresh[137]), .B(cell_1851_and_in[0]), 
        .Z(cell_1851_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1851_a_HPC2_and_U13 ( .A(Fresh[137]), .B(cell_1851_and_in[1]), 
        .Z(cell_1851_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1851_a_HPC2_and_U12 ( .A1(cell_1851_a_HPC2_and_a_reg[1]), .A2(
        cell_1851_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1851_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1851_a_HPC2_and_U11 ( .A1(cell_1851_a_HPC2_and_a_reg[0]), .A2(
        cell_1851_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1851_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1851_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1851_a_HPC2_and_n9), 
        .ZN(cell_1851_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1851_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1851_a_HPC2_and_n9), 
        .ZN(cell_1851_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1851_a_HPC2_and_U8 ( .A(Fresh[137]), .ZN(cell_1851_a_HPC2_and_n9) );
  AND2_X1 cell_1851_a_HPC2_and_U7 ( .A1(cell_1851_and_in[1]), .A2(n422), .ZN(
        cell_1851_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1851_a_HPC2_and_U6 ( .A1(cell_1851_and_in[0]), .A2(n405), .ZN(
        cell_1851_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1851_a_HPC2_and_U5 ( .A(cell_1851_a_HPC2_and_n8), .B(
        cell_1851_a_HPC2_and_z_1__1_), .ZN(cell_1851_and_out[1]) );
  XNOR2_X1 cell_1851_a_HPC2_and_U4 ( .A(
        cell_1851_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1851_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1851_a_HPC2_and_n8) );
  XNOR2_X1 cell_1851_a_HPC2_and_U3 ( .A(cell_1851_a_HPC2_and_n7), .B(
        cell_1851_a_HPC2_and_z_0__0_), .ZN(cell_1851_and_out[0]) );
  XNOR2_X1 cell_1851_a_HPC2_and_U2 ( .A(
        cell_1851_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1851_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1851_a_HPC2_and_n7) );
  DFF_X1 cell_1851_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1851_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1851_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1851_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1851_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1851_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1851_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1851_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1851_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1851_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1852_U4 ( .A(n364), .B(cell_1852_and_out[1]), .Z(signal_3558)
         );
  XOR2_X1 cell_1852_U3 ( .A(n362), .B(cell_1852_and_out[0]), .Z(signal_2120)
         );
  XOR2_X1 cell_1852_U2 ( .A(n364), .B(n371), .Z(cell_1852_and_in[1]) );
  XOR2_X1 cell_1852_U1 ( .A(n362), .B(n369), .Z(cell_1852_and_in[0]) );
  XOR2_X1 cell_1852_a_HPC2_and_U14 ( .A(Fresh[138]), .B(cell_1852_and_in[0]), 
        .Z(cell_1852_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1852_a_HPC2_and_U13 ( .A(Fresh[138]), .B(cell_1852_and_in[1]), 
        .Z(cell_1852_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1852_a_HPC2_and_U12 ( .A1(cell_1852_a_HPC2_and_a_reg[1]), .A2(
        cell_1852_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1852_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1852_a_HPC2_and_U11 ( .A1(cell_1852_a_HPC2_and_a_reg[0]), .A2(
        cell_1852_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1852_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1852_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1852_a_HPC2_and_n9), 
        .ZN(cell_1852_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1852_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1852_a_HPC2_and_n9), 
        .ZN(cell_1852_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1852_a_HPC2_and_U8 ( .A(Fresh[138]), .ZN(cell_1852_a_HPC2_and_n9) );
  AND2_X1 cell_1852_a_HPC2_and_U7 ( .A1(cell_1852_and_in[1]), .A2(n422), .ZN(
        cell_1852_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1852_a_HPC2_and_U6 ( .A1(cell_1852_and_in[0]), .A2(n405), .ZN(
        cell_1852_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1852_a_HPC2_and_U5 ( .A(cell_1852_a_HPC2_and_n8), .B(
        cell_1852_a_HPC2_and_z_1__1_), .ZN(cell_1852_and_out[1]) );
  XNOR2_X1 cell_1852_a_HPC2_and_U4 ( .A(
        cell_1852_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1852_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1852_a_HPC2_and_n8) );
  XNOR2_X1 cell_1852_a_HPC2_and_U3 ( .A(cell_1852_a_HPC2_and_n7), .B(
        cell_1852_a_HPC2_and_z_0__0_), .ZN(cell_1852_and_out[0]) );
  XNOR2_X1 cell_1852_a_HPC2_and_U2 ( .A(
        cell_1852_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1852_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1852_a_HPC2_and_n7) );
  DFF_X1 cell_1852_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1852_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1852_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1852_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1852_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1852_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1852_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1852_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1852_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1852_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1853_U4 ( .A(signal_3404), .B(cell_1853_and_out[1]), .Z(
        signal_3559) );
  XOR2_X1 cell_1853_U3 ( .A(signal_1990), .B(cell_1853_and_out[0]), .Z(
        signal_2121) );
  XOR2_X1 cell_1853_U2 ( .A(signal_3404), .B(n379), .Z(cell_1853_and_in[1]) );
  XOR2_X1 cell_1853_U1 ( .A(signal_1990), .B(n377), .Z(cell_1853_and_in[0]) );
  XOR2_X1 cell_1853_a_HPC2_and_U14 ( .A(Fresh[139]), .B(cell_1853_and_in[0]), 
        .Z(cell_1853_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1853_a_HPC2_and_U13 ( .A(Fresh[139]), .B(cell_1853_and_in[1]), 
        .Z(cell_1853_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1853_a_HPC2_and_U12 ( .A1(cell_1853_a_HPC2_and_a_reg[1]), .A2(
        cell_1853_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1853_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1853_a_HPC2_and_U11 ( .A1(cell_1853_a_HPC2_and_a_reg[0]), .A2(
        cell_1853_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1853_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1853_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1853_a_HPC2_and_n9), 
        .ZN(cell_1853_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1853_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1853_a_HPC2_and_n9), 
        .ZN(cell_1853_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1853_a_HPC2_and_U8 ( .A(Fresh[139]), .ZN(cell_1853_a_HPC2_and_n9) );
  AND2_X1 cell_1853_a_HPC2_and_U7 ( .A1(cell_1853_and_in[1]), .A2(n442), .ZN(
        cell_1853_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1853_a_HPC2_and_U6 ( .A1(cell_1853_and_in[0]), .A2(n428), .ZN(
        cell_1853_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1853_a_HPC2_and_U5 ( .A(cell_1853_a_HPC2_and_n8), .B(
        cell_1853_a_HPC2_and_z_1__1_), .ZN(cell_1853_and_out[1]) );
  XNOR2_X1 cell_1853_a_HPC2_and_U4 ( .A(
        cell_1853_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1853_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1853_a_HPC2_and_n8) );
  XNOR2_X1 cell_1853_a_HPC2_and_U3 ( .A(cell_1853_a_HPC2_and_n7), .B(
        cell_1853_a_HPC2_and_z_0__0_), .ZN(cell_1853_and_out[0]) );
  XNOR2_X1 cell_1853_a_HPC2_and_U2 ( .A(
        cell_1853_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1853_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1853_a_HPC2_and_n7) );
  DFF_X1 cell_1853_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1853_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1853_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1853_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1853_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1853_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1853_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1853_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1853_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1853_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1854_U4 ( .A(n379), .B(cell_1854_and_out[1]), .Z(signal_3560)
         );
  XOR2_X1 cell_1854_U3 ( .A(n377), .B(cell_1854_and_out[0]), .Z(signal_2122)
         );
  XOR2_X1 cell_1854_U2 ( .A(n379), .B(n357), .Z(cell_1854_and_in[1]) );
  XOR2_X1 cell_1854_U1 ( .A(n377), .B(n356), .Z(cell_1854_and_in[0]) );
  XOR2_X1 cell_1854_a_HPC2_and_U14 ( .A(Fresh[140]), .B(cell_1854_and_in[0]), 
        .Z(cell_1854_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1854_a_HPC2_and_U13 ( .A(Fresh[140]), .B(cell_1854_and_in[1]), 
        .Z(cell_1854_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1854_a_HPC2_and_U12 ( .A1(cell_1854_a_HPC2_and_a_reg[1]), .A2(
        cell_1854_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1854_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1854_a_HPC2_and_U11 ( .A1(cell_1854_a_HPC2_and_a_reg[0]), .A2(
        cell_1854_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1854_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1854_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1854_a_HPC2_and_n9), 
        .ZN(cell_1854_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1854_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1854_a_HPC2_and_n9), 
        .ZN(cell_1854_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1854_a_HPC2_and_U8 ( .A(Fresh[140]), .ZN(cell_1854_a_HPC2_and_n9) );
  AND2_X1 cell_1854_a_HPC2_and_U7 ( .A1(cell_1854_and_in[1]), .A2(n422), .ZN(
        cell_1854_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1854_a_HPC2_and_U6 ( .A1(cell_1854_and_in[0]), .A2(n405), .ZN(
        cell_1854_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1854_a_HPC2_and_U5 ( .A(cell_1854_a_HPC2_and_n8), .B(
        cell_1854_a_HPC2_and_z_1__1_), .ZN(cell_1854_and_out[1]) );
  XNOR2_X1 cell_1854_a_HPC2_and_U4 ( .A(
        cell_1854_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1854_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1854_a_HPC2_and_n8) );
  XNOR2_X1 cell_1854_a_HPC2_and_U3 ( .A(cell_1854_a_HPC2_and_n7), .B(
        cell_1854_a_HPC2_and_z_0__0_), .ZN(cell_1854_and_out[0]) );
  XNOR2_X1 cell_1854_a_HPC2_and_U2 ( .A(
        cell_1854_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1854_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1854_a_HPC2_and_n7) );
  DFF_X1 cell_1854_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1854_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1854_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1854_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1854_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1854_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1854_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1854_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1854_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1854_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1855_U4 ( .A(n360), .B(cell_1855_and_out[1]), .Z(signal_3561)
         );
  XOR2_X1 cell_1855_U3 ( .A(n358), .B(cell_1855_and_out[0]), .Z(signal_2123)
         );
  XOR2_X1 cell_1855_U2 ( .A(n360), .B(n375), .Z(cell_1855_and_in[1]) );
  XOR2_X1 cell_1855_U1 ( .A(n358), .B(n373), .Z(cell_1855_and_in[0]) );
  XOR2_X1 cell_1855_a_HPC2_and_U14 ( .A(Fresh[141]), .B(cell_1855_and_in[0]), 
        .Z(cell_1855_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1855_a_HPC2_and_U13 ( .A(Fresh[141]), .B(cell_1855_and_in[1]), 
        .Z(cell_1855_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1855_a_HPC2_and_U12 ( .A1(cell_1855_a_HPC2_and_a_reg[1]), .A2(
        cell_1855_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1855_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1855_a_HPC2_and_U11 ( .A1(cell_1855_a_HPC2_and_a_reg[0]), .A2(
        cell_1855_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1855_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1855_a_HPC2_and_U10 ( .A1(n422), .A2(cell_1855_a_HPC2_and_n9), 
        .ZN(cell_1855_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1855_a_HPC2_and_U9 ( .A1(n405), .A2(cell_1855_a_HPC2_and_n9), 
        .ZN(cell_1855_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1855_a_HPC2_and_U8 ( .A(Fresh[141]), .ZN(cell_1855_a_HPC2_and_n9) );
  AND2_X1 cell_1855_a_HPC2_and_U7 ( .A1(cell_1855_and_in[1]), .A2(n422), .ZN(
        cell_1855_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1855_a_HPC2_and_U6 ( .A1(cell_1855_and_in[0]), .A2(n405), .ZN(
        cell_1855_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1855_a_HPC2_and_U5 ( .A(cell_1855_a_HPC2_and_n8), .B(
        cell_1855_a_HPC2_and_z_1__1_), .ZN(cell_1855_and_out[1]) );
  XNOR2_X1 cell_1855_a_HPC2_and_U4 ( .A(
        cell_1855_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1855_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1855_a_HPC2_and_n8) );
  XNOR2_X1 cell_1855_a_HPC2_and_U3 ( .A(cell_1855_a_HPC2_and_n7), .B(
        cell_1855_a_HPC2_and_z_0__0_), .ZN(cell_1855_and_out[0]) );
  XNOR2_X1 cell_1855_a_HPC2_and_U2 ( .A(
        cell_1855_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1855_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1855_a_HPC2_and_n7) );
  DFF_X1 cell_1855_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1855_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1855_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n405), .CK(clk), 
        .Q(cell_1855_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1855_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1855_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n422), .CK(clk), 
        .Q(cell_1855_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1855_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1855_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1855_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1856_U4 ( .A(n381), .B(cell_1856_and_out[1]), .Z(signal_3562)
         );
  XOR2_X1 cell_1856_U3 ( .A(n380), .B(cell_1856_and_out[0]), .Z(signal_2124)
         );
  XOR2_X1 cell_1856_U2 ( .A(n381), .B(n361), .Z(cell_1856_and_in[1]) );
  XOR2_X1 cell_1856_U1 ( .A(n380), .B(n359), .Z(cell_1856_and_in[0]) );
  XOR2_X1 cell_1856_a_HPC2_and_U14 ( .A(Fresh[142]), .B(cell_1856_and_in[0]), 
        .Z(cell_1856_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1856_a_HPC2_and_U13 ( .A(Fresh[142]), .B(cell_1856_and_in[1]), 
        .Z(cell_1856_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1856_a_HPC2_and_U12 ( .A1(cell_1856_a_HPC2_and_a_reg[1]), .A2(
        cell_1856_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1856_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1856_a_HPC2_and_U11 ( .A1(cell_1856_a_HPC2_and_a_reg[0]), .A2(
        cell_1856_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1856_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1856_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1856_a_HPC2_and_n9), 
        .ZN(cell_1856_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1856_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1856_a_HPC2_and_n9), 
        .ZN(cell_1856_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1856_a_HPC2_and_U8 ( .A(Fresh[142]), .ZN(cell_1856_a_HPC2_and_n9) );
  AND2_X1 cell_1856_a_HPC2_and_U7 ( .A1(cell_1856_and_in[1]), .A2(n423), .ZN(
        cell_1856_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1856_a_HPC2_and_U6 ( .A1(cell_1856_and_in[0]), .A2(n406), .ZN(
        cell_1856_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1856_a_HPC2_and_U5 ( .A(cell_1856_a_HPC2_and_n8), .B(
        cell_1856_a_HPC2_and_z_1__1_), .ZN(cell_1856_and_out[1]) );
  XNOR2_X1 cell_1856_a_HPC2_and_U4 ( .A(
        cell_1856_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1856_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1856_a_HPC2_and_n8) );
  XNOR2_X1 cell_1856_a_HPC2_and_U3 ( .A(cell_1856_a_HPC2_and_n7), .B(
        cell_1856_a_HPC2_and_z_0__0_), .ZN(cell_1856_and_out[0]) );
  XNOR2_X1 cell_1856_a_HPC2_and_U2 ( .A(
        cell_1856_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1856_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1856_a_HPC2_and_n7) );
  DFF_X1 cell_1856_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1856_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1856_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1856_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1856_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1856_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1856_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1856_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1856_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1856_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1857_U4 ( .A(n357), .B(cell_1857_and_out[1]), .Z(signal_3563)
         );
  XOR2_X1 cell_1857_U3 ( .A(n356), .B(cell_1857_and_out[0]), .Z(signal_2125)
         );
  XOR2_X1 cell_1857_U2 ( .A(n357), .B(n361), .Z(cell_1857_and_in[1]) );
  XOR2_X1 cell_1857_U1 ( .A(n356), .B(n359), .Z(cell_1857_and_in[0]) );
  XOR2_X1 cell_1857_a_HPC2_and_U14 ( .A(Fresh[143]), .B(cell_1857_and_in[0]), 
        .Z(cell_1857_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1857_a_HPC2_and_U13 ( .A(Fresh[143]), .B(cell_1857_and_in[1]), 
        .Z(cell_1857_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1857_a_HPC2_and_U12 ( .A1(cell_1857_a_HPC2_and_a_reg[1]), .A2(
        cell_1857_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1857_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1857_a_HPC2_and_U11 ( .A1(cell_1857_a_HPC2_and_a_reg[0]), .A2(
        cell_1857_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1857_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1857_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1857_a_HPC2_and_n9), 
        .ZN(cell_1857_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1857_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1857_a_HPC2_and_n9), 
        .ZN(cell_1857_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1857_a_HPC2_and_U8 ( .A(Fresh[143]), .ZN(cell_1857_a_HPC2_and_n9) );
  AND2_X1 cell_1857_a_HPC2_and_U7 ( .A1(cell_1857_and_in[1]), .A2(n423), .ZN(
        cell_1857_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1857_a_HPC2_and_U6 ( .A1(cell_1857_and_in[0]), .A2(n406), .ZN(
        cell_1857_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1857_a_HPC2_and_U5 ( .A(cell_1857_a_HPC2_and_n8), .B(
        cell_1857_a_HPC2_and_z_1__1_), .ZN(cell_1857_and_out[1]) );
  XNOR2_X1 cell_1857_a_HPC2_and_U4 ( .A(
        cell_1857_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1857_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1857_a_HPC2_and_n8) );
  XNOR2_X1 cell_1857_a_HPC2_and_U3 ( .A(cell_1857_a_HPC2_and_n7), .B(
        cell_1857_a_HPC2_and_z_0__0_), .ZN(cell_1857_and_out[0]) );
  XNOR2_X1 cell_1857_a_HPC2_and_U2 ( .A(
        cell_1857_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1857_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1857_a_HPC2_and_n7) );
  DFF_X1 cell_1857_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1857_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1857_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1857_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1857_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1857_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1857_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1857_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1857_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1857_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1858_U4 ( .A(n367), .B(cell_1858_and_out[1]), .Z(signal_3564)
         );
  XOR2_X1 cell_1858_U3 ( .A(n366), .B(cell_1858_and_out[0]), .Z(signal_2126)
         );
  XOR2_X1 cell_1858_U2 ( .A(n367), .B(1'b0), .Z(cell_1858_and_in[1]) );
  XOR2_X1 cell_1858_U1 ( .A(n366), .B(1'b1), .Z(cell_1858_and_in[0]) );
  XOR2_X1 cell_1858_a_HPC2_and_U14 ( .A(Fresh[144]), .B(cell_1858_and_in[0]), 
        .Z(cell_1858_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1858_a_HPC2_and_U13 ( .A(Fresh[144]), .B(cell_1858_and_in[1]), 
        .Z(cell_1858_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1858_a_HPC2_and_U12 ( .A1(cell_1858_a_HPC2_and_a_reg[1]), .A2(
        cell_1858_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1858_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1858_a_HPC2_and_U11 ( .A1(cell_1858_a_HPC2_and_a_reg[0]), .A2(
        cell_1858_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1858_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1858_a_HPC2_and_U10 ( .A1(n411), .A2(cell_1858_a_HPC2_and_n9), 
        .ZN(cell_1858_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1858_a_HPC2_and_U9 ( .A1(n394), .A2(cell_1858_a_HPC2_and_n9), 
        .ZN(cell_1858_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1858_a_HPC2_and_U8 ( .A(Fresh[144]), .ZN(cell_1858_a_HPC2_and_n9) );
  AND2_X1 cell_1858_a_HPC2_and_U7 ( .A1(cell_1858_and_in[1]), .A2(n411), .ZN(
        cell_1858_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1858_a_HPC2_and_U6 ( .A1(cell_1858_and_in[0]), .A2(n394), .ZN(
        cell_1858_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1858_a_HPC2_and_U5 ( .A(cell_1858_a_HPC2_and_n8), .B(
        cell_1858_a_HPC2_and_z_1__1_), .ZN(cell_1858_and_out[1]) );
  XNOR2_X1 cell_1858_a_HPC2_and_U4 ( .A(
        cell_1858_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1858_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1858_a_HPC2_and_n8) );
  XNOR2_X1 cell_1858_a_HPC2_and_U3 ( .A(cell_1858_a_HPC2_and_n7), .B(
        cell_1858_a_HPC2_and_z_0__0_), .ZN(cell_1858_and_out[0]) );
  XNOR2_X1 cell_1858_a_HPC2_and_U2 ( .A(
        cell_1858_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1858_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1858_a_HPC2_and_n7) );
  DFF_X1 cell_1858_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1858_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1858_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n394), .CK(clk), 
        .Q(cell_1858_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1858_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1858_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n411), .CK(clk), 
        .Q(cell_1858_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1858_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1858_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1858_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1859_U4 ( .A(n360), .B(cell_1859_and_out[1]), .Z(signal_3565)
         );
  XOR2_X1 cell_1859_U3 ( .A(n358), .B(cell_1859_and_out[0]), .Z(signal_2127)
         );
  XOR2_X1 cell_1859_U2 ( .A(n360), .B(1'b0), .Z(cell_1859_and_in[1]) );
  XOR2_X1 cell_1859_U1 ( .A(n358), .B(1'b0), .Z(cell_1859_and_in[0]) );
  XOR2_X1 cell_1859_a_HPC2_and_U14 ( .A(Fresh[145]), .B(cell_1859_and_in[0]), 
        .Z(cell_1859_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1859_a_HPC2_and_U13 ( .A(Fresh[145]), .B(cell_1859_and_in[1]), 
        .Z(cell_1859_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1859_a_HPC2_and_U12 ( .A1(cell_1859_a_HPC2_and_a_reg[1]), .A2(
        cell_1859_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1859_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1859_a_HPC2_and_U11 ( .A1(cell_1859_a_HPC2_and_a_reg[0]), .A2(
        cell_1859_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1859_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1859_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1859_a_HPC2_and_n9), 
        .ZN(cell_1859_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1859_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1859_a_HPC2_and_n9), 
        .ZN(cell_1859_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1859_a_HPC2_and_U8 ( .A(Fresh[145]), .ZN(cell_1859_a_HPC2_and_n9) );
  AND2_X1 cell_1859_a_HPC2_and_U7 ( .A1(cell_1859_and_in[1]), .A2(n426), .ZN(
        cell_1859_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1859_a_HPC2_and_U6 ( .A1(cell_1859_and_in[0]), .A2(n409), .ZN(
        cell_1859_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1859_a_HPC2_and_U5 ( .A(cell_1859_a_HPC2_and_n8), .B(
        cell_1859_a_HPC2_and_z_1__1_), .ZN(cell_1859_and_out[1]) );
  XNOR2_X1 cell_1859_a_HPC2_and_U4 ( .A(
        cell_1859_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1859_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1859_a_HPC2_and_n8) );
  XNOR2_X1 cell_1859_a_HPC2_and_U3 ( .A(cell_1859_a_HPC2_and_n7), .B(
        cell_1859_a_HPC2_and_z_0__0_), .ZN(cell_1859_and_out[0]) );
  XNOR2_X1 cell_1859_a_HPC2_and_U2 ( .A(
        cell_1859_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1859_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1859_a_HPC2_and_n7) );
  DFF_X1 cell_1859_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1859_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1859_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1859_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1859_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1859_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1859_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1859_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1859_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1859_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1860_U4 ( .A(n354), .B(cell_1860_and_out[1]), .Z(signal_3566)
         );
  XOR2_X1 cell_1860_U3 ( .A(n352), .B(cell_1860_and_out[0]), .Z(signal_2128)
         );
  XOR2_X1 cell_1860_U2 ( .A(n354), .B(n379), .Z(cell_1860_and_in[1]) );
  XOR2_X1 cell_1860_U1 ( .A(n352), .B(n377), .Z(cell_1860_and_in[0]) );
  XOR2_X1 cell_1860_a_HPC2_and_U14 ( .A(Fresh[146]), .B(cell_1860_and_in[0]), 
        .Z(cell_1860_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1860_a_HPC2_and_U13 ( .A(Fresh[146]), .B(cell_1860_and_in[1]), 
        .Z(cell_1860_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1860_a_HPC2_and_U12 ( .A1(cell_1860_a_HPC2_and_a_reg[1]), .A2(
        cell_1860_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1860_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1860_a_HPC2_and_U11 ( .A1(cell_1860_a_HPC2_and_a_reg[0]), .A2(
        cell_1860_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1860_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1860_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1860_a_HPC2_and_n9), 
        .ZN(cell_1860_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1860_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1860_a_HPC2_and_n9), 
        .ZN(cell_1860_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1860_a_HPC2_and_U8 ( .A(Fresh[146]), .ZN(cell_1860_a_HPC2_and_n9) );
  AND2_X1 cell_1860_a_HPC2_and_U7 ( .A1(cell_1860_and_in[1]), .A2(n423), .ZN(
        cell_1860_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1860_a_HPC2_and_U6 ( .A1(cell_1860_and_in[0]), .A2(n406), .ZN(
        cell_1860_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1860_a_HPC2_and_U5 ( .A(cell_1860_a_HPC2_and_n8), .B(
        cell_1860_a_HPC2_and_z_1__1_), .ZN(cell_1860_and_out[1]) );
  XNOR2_X1 cell_1860_a_HPC2_and_U4 ( .A(
        cell_1860_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1860_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1860_a_HPC2_and_n8) );
  XNOR2_X1 cell_1860_a_HPC2_and_U3 ( .A(cell_1860_a_HPC2_and_n7), .B(
        cell_1860_a_HPC2_and_z_0__0_), .ZN(cell_1860_and_out[0]) );
  XNOR2_X1 cell_1860_a_HPC2_and_U2 ( .A(
        cell_1860_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1860_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1860_a_HPC2_and_n7) );
  DFF_X1 cell_1860_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1860_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1860_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1860_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1860_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1860_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1860_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1860_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1860_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1860_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1861_U4 ( .A(n357), .B(cell_1861_and_out[1]), .Z(signal_3567)
         );
  XOR2_X1 cell_1861_U3 ( .A(n356), .B(cell_1861_and_out[0]), .Z(signal_2129)
         );
  XOR2_X1 cell_1861_U2 ( .A(n357), .B(signal_3426), .Z(cell_1861_and_in[1]) );
  XOR2_X1 cell_1861_U1 ( .A(n356), .B(signal_2012), .Z(cell_1861_and_in[0]) );
  XOR2_X1 cell_1861_a_HPC2_and_U14 ( .A(Fresh[147]), .B(cell_1861_and_in[0]), 
        .Z(cell_1861_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1861_a_HPC2_and_U13 ( .A(Fresh[147]), .B(cell_1861_and_in[1]), 
        .Z(cell_1861_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1861_a_HPC2_and_U12 ( .A1(cell_1861_a_HPC2_and_a_reg[1]), .A2(
        cell_1861_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1861_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1861_a_HPC2_and_U11 ( .A1(cell_1861_a_HPC2_and_a_reg[0]), .A2(
        cell_1861_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1861_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1861_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1861_a_HPC2_and_n9), 
        .ZN(cell_1861_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1861_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1861_a_HPC2_and_n9), 
        .ZN(cell_1861_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1861_a_HPC2_and_U8 ( .A(Fresh[147]), .ZN(cell_1861_a_HPC2_and_n9) );
  AND2_X1 cell_1861_a_HPC2_and_U7 ( .A1(cell_1861_and_in[1]), .A2(n423), .ZN(
        cell_1861_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1861_a_HPC2_and_U6 ( .A1(cell_1861_and_in[0]), .A2(n406), .ZN(
        cell_1861_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1861_a_HPC2_and_U5 ( .A(cell_1861_a_HPC2_and_n8), .B(
        cell_1861_a_HPC2_and_z_1__1_), .ZN(cell_1861_and_out[1]) );
  XNOR2_X1 cell_1861_a_HPC2_and_U4 ( .A(
        cell_1861_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1861_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1861_a_HPC2_and_n8) );
  XNOR2_X1 cell_1861_a_HPC2_and_U3 ( .A(cell_1861_a_HPC2_and_n7), .B(
        cell_1861_a_HPC2_and_z_0__0_), .ZN(cell_1861_and_out[0]) );
  XNOR2_X1 cell_1861_a_HPC2_and_U2 ( .A(
        cell_1861_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1861_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1861_a_HPC2_and_n7) );
  DFF_X1 cell_1861_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1861_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1861_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1861_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1861_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1861_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1861_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1861_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1861_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1861_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1862_U4 ( .A(n364), .B(cell_1862_and_out[1]), .Z(signal_3568)
         );
  XOR2_X1 cell_1862_U3 ( .A(n362), .B(cell_1862_and_out[0]), .Z(signal_2130)
         );
  XOR2_X1 cell_1862_U2 ( .A(n364), .B(n355), .Z(cell_1862_and_in[1]) );
  XOR2_X1 cell_1862_U1 ( .A(n362), .B(n353), .Z(cell_1862_and_in[0]) );
  XOR2_X1 cell_1862_a_HPC2_and_U14 ( .A(Fresh[148]), .B(cell_1862_and_in[0]), 
        .Z(cell_1862_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1862_a_HPC2_and_U13 ( .A(Fresh[148]), .B(cell_1862_and_in[1]), 
        .Z(cell_1862_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1862_a_HPC2_and_U12 ( .A1(cell_1862_a_HPC2_and_a_reg[1]), .A2(
        cell_1862_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1862_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1862_a_HPC2_and_U11 ( .A1(cell_1862_a_HPC2_and_a_reg[0]), .A2(
        cell_1862_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1862_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1862_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1862_a_HPC2_and_n9), 
        .ZN(cell_1862_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1862_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1862_a_HPC2_and_n9), 
        .ZN(cell_1862_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1862_a_HPC2_and_U8 ( .A(Fresh[148]), .ZN(cell_1862_a_HPC2_and_n9) );
  AND2_X1 cell_1862_a_HPC2_and_U7 ( .A1(cell_1862_and_in[1]), .A2(n423), .ZN(
        cell_1862_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1862_a_HPC2_and_U6 ( .A1(cell_1862_and_in[0]), .A2(n406), .ZN(
        cell_1862_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1862_a_HPC2_and_U5 ( .A(cell_1862_a_HPC2_and_n8), .B(
        cell_1862_a_HPC2_and_z_1__1_), .ZN(cell_1862_and_out[1]) );
  XNOR2_X1 cell_1862_a_HPC2_and_U4 ( .A(
        cell_1862_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1862_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1862_a_HPC2_and_n8) );
  XNOR2_X1 cell_1862_a_HPC2_and_U3 ( .A(cell_1862_a_HPC2_and_n7), .B(
        cell_1862_a_HPC2_and_z_0__0_), .ZN(cell_1862_and_out[0]) );
  XNOR2_X1 cell_1862_a_HPC2_and_U2 ( .A(
        cell_1862_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1862_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1862_a_HPC2_and_n7) );
  DFF_X1 cell_1862_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1862_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1862_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1862_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1862_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1862_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1862_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1862_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1862_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1862_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1863_U4 ( .A(n361), .B(cell_1863_and_out[1]), .Z(signal_3569)
         );
  XOR2_X1 cell_1863_U3 ( .A(n359), .B(cell_1863_and_out[0]), .Z(signal_2131)
         );
  XOR2_X1 cell_1863_U2 ( .A(n361), .B(signal_3261), .Z(cell_1863_and_in[1]) );
  XOR2_X1 cell_1863_U1 ( .A(n359), .B(signal_1987), .Z(cell_1863_and_in[0]) );
  XOR2_X1 cell_1863_a_HPC2_and_U14 ( .A(Fresh[149]), .B(cell_1863_and_in[0]), 
        .Z(cell_1863_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1863_a_HPC2_and_U13 ( .A(Fresh[149]), .B(cell_1863_and_in[1]), 
        .Z(cell_1863_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1863_a_HPC2_and_U12 ( .A1(cell_1863_a_HPC2_and_a_reg[1]), .A2(
        cell_1863_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1863_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1863_a_HPC2_and_U11 ( .A1(cell_1863_a_HPC2_and_a_reg[0]), .A2(
        cell_1863_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1863_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1863_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1863_a_HPC2_and_n9), 
        .ZN(cell_1863_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1863_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1863_a_HPC2_and_n9), 
        .ZN(cell_1863_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1863_a_HPC2_and_U8 ( .A(Fresh[149]), .ZN(cell_1863_a_HPC2_and_n9) );
  AND2_X1 cell_1863_a_HPC2_and_U7 ( .A1(cell_1863_and_in[1]), .A2(n423), .ZN(
        cell_1863_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1863_a_HPC2_and_U6 ( .A1(cell_1863_and_in[0]), .A2(n406), .ZN(
        cell_1863_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1863_a_HPC2_and_U5 ( .A(cell_1863_a_HPC2_and_n8), .B(
        cell_1863_a_HPC2_and_z_1__1_), .ZN(cell_1863_and_out[1]) );
  XNOR2_X1 cell_1863_a_HPC2_and_U4 ( .A(
        cell_1863_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1863_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1863_a_HPC2_and_n8) );
  XNOR2_X1 cell_1863_a_HPC2_and_U3 ( .A(cell_1863_a_HPC2_and_n7), .B(
        cell_1863_a_HPC2_and_z_0__0_), .ZN(cell_1863_and_out[0]) );
  XNOR2_X1 cell_1863_a_HPC2_and_U2 ( .A(
        cell_1863_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1863_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1863_a_HPC2_and_n7) );
  DFF_X1 cell_1863_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1863_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1863_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1863_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1863_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1863_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1863_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1863_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1863_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1863_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1864_U4 ( .A(n367), .B(cell_1864_and_out[1]), .Z(signal_3570)
         );
  XOR2_X1 cell_1864_U3 ( .A(n366), .B(cell_1864_and_out[0]), .Z(signal_2132)
         );
  XOR2_X1 cell_1864_U2 ( .A(n367), .B(n379), .Z(cell_1864_and_in[1]) );
  XOR2_X1 cell_1864_U1 ( .A(n366), .B(n377), .Z(cell_1864_and_in[0]) );
  XOR2_X1 cell_1864_a_HPC2_and_U14 ( .A(Fresh[150]), .B(cell_1864_and_in[0]), 
        .Z(cell_1864_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1864_a_HPC2_and_U13 ( .A(Fresh[150]), .B(cell_1864_and_in[1]), 
        .Z(cell_1864_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1864_a_HPC2_and_U12 ( .A1(cell_1864_a_HPC2_and_a_reg[1]), .A2(
        cell_1864_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1864_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1864_a_HPC2_and_U11 ( .A1(cell_1864_a_HPC2_and_a_reg[0]), .A2(
        cell_1864_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1864_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1864_a_HPC2_and_U10 ( .A1(n423), .A2(cell_1864_a_HPC2_and_n9), 
        .ZN(cell_1864_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1864_a_HPC2_and_U9 ( .A1(n406), .A2(cell_1864_a_HPC2_and_n9), 
        .ZN(cell_1864_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1864_a_HPC2_and_U8 ( .A(Fresh[150]), .ZN(cell_1864_a_HPC2_and_n9) );
  AND2_X1 cell_1864_a_HPC2_and_U7 ( .A1(cell_1864_and_in[1]), .A2(n423), .ZN(
        cell_1864_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1864_a_HPC2_and_U6 ( .A1(cell_1864_and_in[0]), .A2(n406), .ZN(
        cell_1864_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1864_a_HPC2_and_U5 ( .A(cell_1864_a_HPC2_and_n8), .B(
        cell_1864_a_HPC2_and_z_1__1_), .ZN(cell_1864_and_out[1]) );
  XNOR2_X1 cell_1864_a_HPC2_and_U4 ( .A(
        cell_1864_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1864_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1864_a_HPC2_and_n8) );
  XNOR2_X1 cell_1864_a_HPC2_and_U3 ( .A(cell_1864_a_HPC2_and_n7), .B(
        cell_1864_a_HPC2_and_z_0__0_), .ZN(cell_1864_and_out[0]) );
  XNOR2_X1 cell_1864_a_HPC2_and_U2 ( .A(
        cell_1864_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1864_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1864_a_HPC2_and_n7) );
  DFF_X1 cell_1864_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1864_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1864_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n406), .CK(clk), 
        .Q(cell_1864_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1864_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1864_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n423), .CK(clk), 
        .Q(cell_1864_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1864_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1864_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1864_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1865_U4 ( .A(1'b0), .B(cell_1865_and_out[1]), .Z(signal_3571)
         );
  XOR2_X1 cell_1865_U3 ( .A(1'b0), .B(cell_1865_and_out[0]), .Z(signal_2133)
         );
  XOR2_X1 cell_1865_U2 ( .A(1'b0), .B(n357), .Z(cell_1865_and_in[1]) );
  XOR2_X1 cell_1865_U1 ( .A(1'b0), .B(n356), .Z(cell_1865_and_in[0]) );
  XOR2_X1 cell_1865_a_HPC2_and_U14 ( .A(Fresh[151]), .B(cell_1865_and_in[0]), 
        .Z(cell_1865_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1865_a_HPC2_and_U13 ( .A(Fresh[151]), .B(cell_1865_and_in[1]), 
        .Z(cell_1865_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1865_a_HPC2_and_U12 ( .A1(cell_1865_a_HPC2_and_a_reg[1]), .A2(
        cell_1865_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1865_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1865_a_HPC2_and_U11 ( .A1(cell_1865_a_HPC2_and_a_reg[0]), .A2(
        cell_1865_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1865_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1865_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1865_a_HPC2_and_n9), 
        .ZN(cell_1865_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1865_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1865_a_HPC2_and_n9), 
        .ZN(cell_1865_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1865_a_HPC2_and_U8 ( .A(Fresh[151]), .ZN(cell_1865_a_HPC2_and_n9) );
  AND2_X1 cell_1865_a_HPC2_and_U7 ( .A1(cell_1865_and_in[1]), .A2(n425), .ZN(
        cell_1865_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1865_a_HPC2_and_U6 ( .A1(cell_1865_and_in[0]), .A2(n408), .ZN(
        cell_1865_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1865_a_HPC2_and_U5 ( .A(cell_1865_a_HPC2_and_n8), .B(
        cell_1865_a_HPC2_and_z_1__1_), .ZN(cell_1865_and_out[1]) );
  XNOR2_X1 cell_1865_a_HPC2_and_U4 ( .A(
        cell_1865_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1865_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1865_a_HPC2_and_n8) );
  XNOR2_X1 cell_1865_a_HPC2_and_U3 ( .A(cell_1865_a_HPC2_and_n7), .B(
        cell_1865_a_HPC2_and_z_0__0_), .ZN(cell_1865_and_out[0]) );
  XNOR2_X1 cell_1865_a_HPC2_and_U2 ( .A(
        cell_1865_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1865_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1865_a_HPC2_and_n7) );
  DFF_X1 cell_1865_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1865_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1865_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1865_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1865_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1865_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1865_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1865_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1865_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1865_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1866_U4 ( .A(n360), .B(cell_1866_and_out[1]), .Z(signal_3572)
         );
  XOR2_X1 cell_1866_U3 ( .A(n358), .B(cell_1866_and_out[0]), .Z(signal_2134)
         );
  XOR2_X1 cell_1866_U2 ( .A(n360), .B(n365), .Z(cell_1866_and_in[1]) );
  XOR2_X1 cell_1866_U1 ( .A(n358), .B(n363), .Z(cell_1866_and_in[0]) );
  XOR2_X1 cell_1866_a_HPC2_and_U14 ( .A(Fresh[152]), .B(cell_1866_and_in[0]), 
        .Z(cell_1866_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1866_a_HPC2_and_U13 ( .A(Fresh[152]), .B(cell_1866_and_in[1]), 
        .Z(cell_1866_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1866_a_HPC2_and_U12 ( .A1(cell_1866_a_HPC2_and_a_reg[1]), .A2(
        cell_1866_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1866_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1866_a_HPC2_and_U11 ( .A1(cell_1866_a_HPC2_and_a_reg[0]), .A2(
        cell_1866_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1866_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1866_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1866_a_HPC2_and_n9), 
        .ZN(cell_1866_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1866_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1866_a_HPC2_and_n9), 
        .ZN(cell_1866_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1866_a_HPC2_and_U8 ( .A(Fresh[152]), .ZN(cell_1866_a_HPC2_and_n9) );
  AND2_X1 cell_1866_a_HPC2_and_U7 ( .A1(cell_1866_and_in[1]), .A2(n424), .ZN(
        cell_1866_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1866_a_HPC2_and_U6 ( .A1(cell_1866_and_in[0]), .A2(n407), .ZN(
        cell_1866_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1866_a_HPC2_and_U5 ( .A(cell_1866_a_HPC2_and_n8), .B(
        cell_1866_a_HPC2_and_z_1__1_), .ZN(cell_1866_and_out[1]) );
  XNOR2_X1 cell_1866_a_HPC2_and_U4 ( .A(
        cell_1866_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1866_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1866_a_HPC2_and_n8) );
  XNOR2_X1 cell_1866_a_HPC2_and_U3 ( .A(cell_1866_a_HPC2_and_n7), .B(
        cell_1866_a_HPC2_and_z_0__0_), .ZN(cell_1866_and_out[0]) );
  XNOR2_X1 cell_1866_a_HPC2_and_U2 ( .A(
        cell_1866_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1866_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1866_a_HPC2_and_n7) );
  DFF_X1 cell_1866_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1866_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1866_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1866_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1866_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1866_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1866_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1866_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1866_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1866_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1867_U4 ( .A(n383), .B(cell_1867_and_out[1]), .Z(signal_3573)
         );
  XOR2_X1 cell_1867_U3 ( .A(n382), .B(cell_1867_and_out[0]), .Z(signal_2135)
         );
  XOR2_X1 cell_1867_U2 ( .A(n383), .B(n360), .Z(cell_1867_and_in[1]) );
  XOR2_X1 cell_1867_U1 ( .A(n382), .B(n358), .Z(cell_1867_and_in[0]) );
  XOR2_X1 cell_1867_a_HPC2_and_U14 ( .A(Fresh[153]), .B(cell_1867_and_in[0]), 
        .Z(cell_1867_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1867_a_HPC2_and_U13 ( .A(Fresh[153]), .B(cell_1867_and_in[1]), 
        .Z(cell_1867_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1867_a_HPC2_and_U12 ( .A1(cell_1867_a_HPC2_and_a_reg[1]), .A2(
        cell_1867_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1867_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1867_a_HPC2_and_U11 ( .A1(cell_1867_a_HPC2_and_a_reg[0]), .A2(
        cell_1867_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1867_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1867_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1867_a_HPC2_and_n9), 
        .ZN(cell_1867_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1867_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1867_a_HPC2_and_n9), 
        .ZN(cell_1867_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1867_a_HPC2_and_U8 ( .A(Fresh[153]), .ZN(cell_1867_a_HPC2_and_n9) );
  AND2_X1 cell_1867_a_HPC2_and_U7 ( .A1(cell_1867_and_in[1]), .A2(n424), .ZN(
        cell_1867_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1867_a_HPC2_and_U6 ( .A1(cell_1867_and_in[0]), .A2(n407), .ZN(
        cell_1867_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1867_a_HPC2_and_U5 ( .A(cell_1867_a_HPC2_and_n8), .B(
        cell_1867_a_HPC2_and_z_1__1_), .ZN(cell_1867_and_out[1]) );
  XNOR2_X1 cell_1867_a_HPC2_and_U4 ( .A(
        cell_1867_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1867_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1867_a_HPC2_and_n8) );
  XNOR2_X1 cell_1867_a_HPC2_and_U3 ( .A(cell_1867_a_HPC2_and_n7), .B(
        cell_1867_a_HPC2_and_z_0__0_), .ZN(cell_1867_and_out[0]) );
  XNOR2_X1 cell_1867_a_HPC2_and_U2 ( .A(
        cell_1867_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1867_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1867_a_HPC2_and_n7) );
  DFF_X1 cell_1867_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1867_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1867_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1867_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1867_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1867_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1867_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1867_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1867_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1867_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1868_U4 ( .A(n379), .B(cell_1868_and_out[1]), .Z(signal_3574)
         );
  XOR2_X1 cell_1868_U3 ( .A(n377), .B(cell_1868_and_out[0]), .Z(signal_2136)
         );
  XOR2_X1 cell_1868_U2 ( .A(n379), .B(n367), .Z(cell_1868_and_in[1]) );
  XOR2_X1 cell_1868_U1 ( .A(n377), .B(n366), .Z(cell_1868_and_in[0]) );
  XOR2_X1 cell_1868_a_HPC2_and_U14 ( .A(Fresh[154]), .B(cell_1868_and_in[0]), 
        .Z(cell_1868_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1868_a_HPC2_and_U13 ( .A(Fresh[154]), .B(cell_1868_and_in[1]), 
        .Z(cell_1868_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1868_a_HPC2_and_U12 ( .A1(cell_1868_a_HPC2_and_a_reg[1]), .A2(
        cell_1868_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1868_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1868_a_HPC2_and_U11 ( .A1(cell_1868_a_HPC2_and_a_reg[0]), .A2(
        cell_1868_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1868_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1868_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1868_a_HPC2_and_n9), 
        .ZN(cell_1868_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1868_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1868_a_HPC2_and_n9), 
        .ZN(cell_1868_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1868_a_HPC2_and_U8 ( .A(Fresh[154]), .ZN(cell_1868_a_HPC2_and_n9) );
  AND2_X1 cell_1868_a_HPC2_and_U7 ( .A1(cell_1868_and_in[1]), .A2(n424), .ZN(
        cell_1868_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1868_a_HPC2_and_U6 ( .A1(cell_1868_and_in[0]), .A2(n407), .ZN(
        cell_1868_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1868_a_HPC2_and_U5 ( .A(cell_1868_a_HPC2_and_n8), .B(
        cell_1868_a_HPC2_and_z_1__1_), .ZN(cell_1868_and_out[1]) );
  XNOR2_X1 cell_1868_a_HPC2_and_U4 ( .A(
        cell_1868_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1868_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1868_a_HPC2_and_n8) );
  XNOR2_X1 cell_1868_a_HPC2_and_U3 ( .A(cell_1868_a_HPC2_and_n7), .B(
        cell_1868_a_HPC2_and_z_0__0_), .ZN(cell_1868_and_out[0]) );
  XNOR2_X1 cell_1868_a_HPC2_and_U2 ( .A(
        cell_1868_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1868_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1868_a_HPC2_and_n7) );
  DFF_X1 cell_1868_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1868_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1868_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1868_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1868_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1868_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1868_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1868_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1868_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1868_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1869_U4 ( .A(n364), .B(cell_1869_and_out[1]), .Z(signal_3575)
         );
  XOR2_X1 cell_1869_U3 ( .A(n362), .B(cell_1869_and_out[0]), .Z(signal_2137)
         );
  XOR2_X1 cell_1869_U2 ( .A(n364), .B(signal_3413), .Z(cell_1869_and_in[1]) );
  XOR2_X1 cell_1869_U1 ( .A(n362), .B(signal_1999), .Z(cell_1869_and_in[0]) );
  XOR2_X1 cell_1869_a_HPC2_and_U14 ( .A(Fresh[155]), .B(cell_1869_and_in[0]), 
        .Z(cell_1869_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1869_a_HPC2_and_U13 ( .A(Fresh[155]), .B(cell_1869_and_in[1]), 
        .Z(cell_1869_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1869_a_HPC2_and_U12 ( .A1(cell_1869_a_HPC2_and_a_reg[1]), .A2(
        cell_1869_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1869_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1869_a_HPC2_and_U11 ( .A1(cell_1869_a_HPC2_and_a_reg[0]), .A2(
        cell_1869_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1869_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1869_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1869_a_HPC2_and_n9), 
        .ZN(cell_1869_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1869_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1869_a_HPC2_and_n9), 
        .ZN(cell_1869_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1869_a_HPC2_and_U8 ( .A(Fresh[155]), .ZN(cell_1869_a_HPC2_and_n9) );
  AND2_X1 cell_1869_a_HPC2_and_U7 ( .A1(cell_1869_and_in[1]), .A2(n424), .ZN(
        cell_1869_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1869_a_HPC2_and_U6 ( .A1(cell_1869_and_in[0]), .A2(n407), .ZN(
        cell_1869_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1869_a_HPC2_and_U5 ( .A(cell_1869_a_HPC2_and_n8), .B(
        cell_1869_a_HPC2_and_z_1__1_), .ZN(cell_1869_and_out[1]) );
  XNOR2_X1 cell_1869_a_HPC2_and_U4 ( .A(
        cell_1869_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1869_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1869_a_HPC2_and_n8) );
  XNOR2_X1 cell_1869_a_HPC2_and_U3 ( .A(cell_1869_a_HPC2_and_n7), .B(
        cell_1869_a_HPC2_and_z_0__0_), .ZN(cell_1869_and_out[0]) );
  XNOR2_X1 cell_1869_a_HPC2_and_U2 ( .A(
        cell_1869_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1869_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1869_a_HPC2_and_n7) );
  DFF_X1 cell_1869_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1869_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1869_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1869_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1869_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1869_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1869_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1869_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1869_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1869_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1870_U4 ( .A(n370), .B(cell_1870_and_out[1]), .Z(signal_3576)
         );
  XOR2_X1 cell_1870_U3 ( .A(n368), .B(cell_1870_and_out[0]), .Z(signal_2138)
         );
  XOR2_X1 cell_1870_U2 ( .A(n370), .B(signal_3406), .Z(cell_1870_and_in[1]) );
  XOR2_X1 cell_1870_U1 ( .A(n368), .B(signal_1992), .Z(cell_1870_and_in[0]) );
  XOR2_X1 cell_1870_a_HPC2_and_U14 ( .A(Fresh[156]), .B(cell_1870_and_in[0]), 
        .Z(cell_1870_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1870_a_HPC2_and_U13 ( .A(Fresh[156]), .B(cell_1870_and_in[1]), 
        .Z(cell_1870_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1870_a_HPC2_and_U12 ( .A1(cell_1870_a_HPC2_and_a_reg[1]), .A2(
        cell_1870_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1870_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1870_a_HPC2_and_U11 ( .A1(cell_1870_a_HPC2_and_a_reg[0]), .A2(
        cell_1870_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1870_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1870_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1870_a_HPC2_and_n9), 
        .ZN(cell_1870_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1870_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1870_a_HPC2_and_n9), 
        .ZN(cell_1870_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1870_a_HPC2_and_U8 ( .A(Fresh[156]), .ZN(cell_1870_a_HPC2_and_n9) );
  AND2_X1 cell_1870_a_HPC2_and_U7 ( .A1(cell_1870_and_in[1]), .A2(n424), .ZN(
        cell_1870_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1870_a_HPC2_and_U6 ( .A1(cell_1870_and_in[0]), .A2(n407), .ZN(
        cell_1870_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1870_a_HPC2_and_U5 ( .A(cell_1870_a_HPC2_and_n8), .B(
        cell_1870_a_HPC2_and_z_1__1_), .ZN(cell_1870_and_out[1]) );
  XNOR2_X1 cell_1870_a_HPC2_and_U4 ( .A(
        cell_1870_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1870_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1870_a_HPC2_and_n8) );
  XNOR2_X1 cell_1870_a_HPC2_and_U3 ( .A(cell_1870_a_HPC2_and_n7), .B(
        cell_1870_a_HPC2_and_z_0__0_), .ZN(cell_1870_and_out[0]) );
  XNOR2_X1 cell_1870_a_HPC2_and_U2 ( .A(
        cell_1870_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1870_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1870_a_HPC2_and_n7) );
  DFF_X1 cell_1870_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1870_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1870_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1870_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1870_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1870_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1870_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1870_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1870_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1870_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1871_U4 ( .A(n370), .B(cell_1871_and_out[1]), .Z(signal_3577)
         );
  XOR2_X1 cell_1871_U3 ( .A(n368), .B(cell_1871_and_out[0]), .Z(signal_2139)
         );
  XOR2_X1 cell_1871_U2 ( .A(n370), .B(signal_3413), .Z(cell_1871_and_in[1]) );
  XOR2_X1 cell_1871_U1 ( .A(n368), .B(signal_1999), .Z(cell_1871_and_in[0]) );
  XOR2_X1 cell_1871_a_HPC2_and_U14 ( .A(Fresh[157]), .B(cell_1871_and_in[0]), 
        .Z(cell_1871_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1871_a_HPC2_and_U13 ( .A(Fresh[157]), .B(cell_1871_and_in[1]), 
        .Z(cell_1871_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1871_a_HPC2_and_U12 ( .A1(cell_1871_a_HPC2_and_a_reg[1]), .A2(
        cell_1871_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1871_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1871_a_HPC2_and_U11 ( .A1(cell_1871_a_HPC2_and_a_reg[0]), .A2(
        cell_1871_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1871_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1871_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1871_a_HPC2_and_n9), 
        .ZN(cell_1871_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1871_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1871_a_HPC2_and_n9), 
        .ZN(cell_1871_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1871_a_HPC2_and_U8 ( .A(Fresh[157]), .ZN(cell_1871_a_HPC2_and_n9) );
  AND2_X1 cell_1871_a_HPC2_and_U7 ( .A1(cell_1871_and_in[1]), .A2(n424), .ZN(
        cell_1871_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1871_a_HPC2_and_U6 ( .A1(cell_1871_and_in[0]), .A2(n407), .ZN(
        cell_1871_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1871_a_HPC2_and_U5 ( .A(cell_1871_a_HPC2_and_n8), .B(
        cell_1871_a_HPC2_and_z_1__1_), .ZN(cell_1871_and_out[1]) );
  XNOR2_X1 cell_1871_a_HPC2_and_U4 ( .A(
        cell_1871_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1871_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1871_a_HPC2_and_n8) );
  XNOR2_X1 cell_1871_a_HPC2_and_U3 ( .A(cell_1871_a_HPC2_and_n7), .B(
        cell_1871_a_HPC2_and_z_0__0_), .ZN(cell_1871_and_out[0]) );
  XNOR2_X1 cell_1871_a_HPC2_and_U2 ( .A(
        cell_1871_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1871_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1871_a_HPC2_and_n7) );
  DFF_X1 cell_1871_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1871_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1871_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1871_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1871_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1871_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1871_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1871_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1871_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1871_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1872_U4 ( .A(n360), .B(cell_1872_and_out[1]), .Z(signal_3578)
         );
  XOR2_X1 cell_1872_U3 ( .A(n358), .B(cell_1872_and_out[0]), .Z(signal_2140)
         );
  XOR2_X1 cell_1872_U2 ( .A(n360), .B(n383), .Z(cell_1872_and_in[1]) );
  XOR2_X1 cell_1872_U1 ( .A(n358), .B(n382), .Z(cell_1872_and_in[0]) );
  XOR2_X1 cell_1872_a_HPC2_and_U14 ( .A(Fresh[158]), .B(cell_1872_and_in[0]), 
        .Z(cell_1872_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1872_a_HPC2_and_U13 ( .A(Fresh[158]), .B(cell_1872_and_in[1]), 
        .Z(cell_1872_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1872_a_HPC2_and_U12 ( .A1(cell_1872_a_HPC2_and_a_reg[1]), .A2(
        cell_1872_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1872_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1872_a_HPC2_and_U11 ( .A1(cell_1872_a_HPC2_and_a_reg[0]), .A2(
        cell_1872_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1872_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1872_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1872_a_HPC2_and_n9), 
        .ZN(cell_1872_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1872_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1872_a_HPC2_and_n9), 
        .ZN(cell_1872_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1872_a_HPC2_and_U8 ( .A(Fresh[158]), .ZN(cell_1872_a_HPC2_and_n9) );
  AND2_X1 cell_1872_a_HPC2_and_U7 ( .A1(cell_1872_and_in[1]), .A2(n424), .ZN(
        cell_1872_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1872_a_HPC2_and_U6 ( .A1(cell_1872_and_in[0]), .A2(n407), .ZN(
        cell_1872_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1872_a_HPC2_and_U5 ( .A(cell_1872_a_HPC2_and_n8), .B(
        cell_1872_a_HPC2_and_z_1__1_), .ZN(cell_1872_and_out[1]) );
  XNOR2_X1 cell_1872_a_HPC2_and_U4 ( .A(
        cell_1872_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1872_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1872_a_HPC2_and_n8) );
  XNOR2_X1 cell_1872_a_HPC2_and_U3 ( .A(cell_1872_a_HPC2_and_n7), .B(
        cell_1872_a_HPC2_and_z_0__0_), .ZN(cell_1872_and_out[0]) );
  XNOR2_X1 cell_1872_a_HPC2_and_U2 ( .A(
        cell_1872_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1872_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1872_a_HPC2_and_n7) );
  DFF_X1 cell_1872_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1872_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1872_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1872_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1872_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1872_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1872_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1872_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1872_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1872_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1873_U4 ( .A(n357), .B(cell_1873_and_out[1]), .Z(signal_3579)
         );
  XOR2_X1 cell_1873_U3 ( .A(n356), .B(cell_1873_and_out[0]), .Z(signal_2141)
         );
  XOR2_X1 cell_1873_U2 ( .A(n357), .B(n379), .Z(cell_1873_and_in[1]) );
  XOR2_X1 cell_1873_U1 ( .A(n356), .B(n377), .Z(cell_1873_and_in[0]) );
  XOR2_X1 cell_1873_a_HPC2_and_U14 ( .A(Fresh[159]), .B(cell_1873_and_in[0]), 
        .Z(cell_1873_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1873_a_HPC2_and_U13 ( .A(Fresh[159]), .B(cell_1873_and_in[1]), 
        .Z(cell_1873_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1873_a_HPC2_and_U12 ( .A1(cell_1873_a_HPC2_and_a_reg[1]), .A2(
        cell_1873_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1873_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1873_a_HPC2_and_U11 ( .A1(cell_1873_a_HPC2_and_a_reg[0]), .A2(
        cell_1873_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1873_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1873_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1873_a_HPC2_and_n9), 
        .ZN(cell_1873_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1873_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1873_a_HPC2_and_n9), 
        .ZN(cell_1873_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1873_a_HPC2_and_U8 ( .A(Fresh[159]), .ZN(cell_1873_a_HPC2_and_n9) );
  AND2_X1 cell_1873_a_HPC2_and_U7 ( .A1(cell_1873_and_in[1]), .A2(n425), .ZN(
        cell_1873_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1873_a_HPC2_and_U6 ( .A1(cell_1873_and_in[0]), .A2(n408), .ZN(
        cell_1873_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1873_a_HPC2_and_U5 ( .A(cell_1873_a_HPC2_and_n8), .B(
        cell_1873_a_HPC2_and_z_1__1_), .ZN(cell_1873_and_out[1]) );
  XNOR2_X1 cell_1873_a_HPC2_and_U4 ( .A(
        cell_1873_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1873_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1873_a_HPC2_and_n8) );
  XNOR2_X1 cell_1873_a_HPC2_and_U3 ( .A(cell_1873_a_HPC2_and_n7), .B(
        cell_1873_a_HPC2_and_z_0__0_), .ZN(cell_1873_and_out[0]) );
  XNOR2_X1 cell_1873_a_HPC2_and_U2 ( .A(
        cell_1873_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1873_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1873_a_HPC2_and_n7) );
  DFF_X1 cell_1873_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1873_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1873_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1873_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1873_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1873_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1873_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1873_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1873_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1873_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1874_U4 ( .A(n367), .B(cell_1874_and_out[1]), .Z(signal_3580)
         );
  XOR2_X1 cell_1874_U3 ( .A(n366), .B(cell_1874_and_out[0]), .Z(signal_2142)
         );
  XOR2_X1 cell_1874_U2 ( .A(n367), .B(signal_3261), .Z(cell_1874_and_in[1]) );
  XOR2_X1 cell_1874_U1 ( .A(n366), .B(signal_1987), .Z(cell_1874_and_in[0]) );
  XOR2_X1 cell_1874_a_HPC2_and_U14 ( .A(Fresh[160]), .B(cell_1874_and_in[0]), 
        .Z(cell_1874_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1874_a_HPC2_and_U13 ( .A(Fresh[160]), .B(cell_1874_and_in[1]), 
        .Z(cell_1874_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1874_a_HPC2_and_U12 ( .A1(cell_1874_a_HPC2_and_a_reg[1]), .A2(
        cell_1874_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1874_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1874_a_HPC2_and_U11 ( .A1(cell_1874_a_HPC2_and_a_reg[0]), .A2(
        cell_1874_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1874_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1874_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1874_a_HPC2_and_n9), 
        .ZN(cell_1874_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1874_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1874_a_HPC2_and_n9), 
        .ZN(cell_1874_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1874_a_HPC2_and_U8 ( .A(Fresh[160]), .ZN(cell_1874_a_HPC2_and_n9) );
  AND2_X1 cell_1874_a_HPC2_and_U7 ( .A1(cell_1874_and_in[1]), .A2(n425), .ZN(
        cell_1874_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1874_a_HPC2_and_U6 ( .A1(cell_1874_and_in[0]), .A2(n408), .ZN(
        cell_1874_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1874_a_HPC2_and_U5 ( .A(cell_1874_a_HPC2_and_n8), .B(
        cell_1874_a_HPC2_and_z_1__1_), .ZN(cell_1874_and_out[1]) );
  XNOR2_X1 cell_1874_a_HPC2_and_U4 ( .A(
        cell_1874_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1874_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1874_a_HPC2_and_n8) );
  XNOR2_X1 cell_1874_a_HPC2_and_U3 ( .A(cell_1874_a_HPC2_and_n7), .B(
        cell_1874_a_HPC2_and_z_0__0_), .ZN(cell_1874_and_out[0]) );
  XNOR2_X1 cell_1874_a_HPC2_and_U2 ( .A(
        cell_1874_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1874_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1874_a_HPC2_and_n7) );
  DFF_X1 cell_1874_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1874_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1874_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1874_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1874_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1874_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1874_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1874_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1874_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1874_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1875_U4 ( .A(n364), .B(cell_1875_and_out[1]), .Z(signal_3581)
         );
  XOR2_X1 cell_1875_U3 ( .A(n362), .B(cell_1875_and_out[0]), .Z(signal_2143)
         );
  XOR2_X1 cell_1875_U2 ( .A(n364), .B(n360), .Z(cell_1875_and_in[1]) );
  XOR2_X1 cell_1875_U1 ( .A(n362), .B(n358), .Z(cell_1875_and_in[0]) );
  XOR2_X1 cell_1875_a_HPC2_and_U14 ( .A(Fresh[161]), .B(cell_1875_and_in[0]), 
        .Z(cell_1875_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1875_a_HPC2_and_U13 ( .A(Fresh[161]), .B(cell_1875_and_in[1]), 
        .Z(cell_1875_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1875_a_HPC2_and_U12 ( .A1(cell_1875_a_HPC2_and_a_reg[1]), .A2(
        cell_1875_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1875_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1875_a_HPC2_and_U11 ( .A1(cell_1875_a_HPC2_and_a_reg[0]), .A2(
        cell_1875_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1875_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1875_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1875_a_HPC2_and_n9), 
        .ZN(cell_1875_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1875_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1875_a_HPC2_and_n9), 
        .ZN(cell_1875_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1875_a_HPC2_and_U8 ( .A(Fresh[161]), .ZN(cell_1875_a_HPC2_and_n9) );
  AND2_X1 cell_1875_a_HPC2_and_U7 ( .A1(cell_1875_and_in[1]), .A2(n425), .ZN(
        cell_1875_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1875_a_HPC2_and_U6 ( .A1(cell_1875_and_in[0]), .A2(n408), .ZN(
        cell_1875_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1875_a_HPC2_and_U5 ( .A(cell_1875_a_HPC2_and_n8), .B(
        cell_1875_a_HPC2_and_z_1__1_), .ZN(cell_1875_and_out[1]) );
  XNOR2_X1 cell_1875_a_HPC2_and_U4 ( .A(
        cell_1875_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1875_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1875_a_HPC2_and_n8) );
  XNOR2_X1 cell_1875_a_HPC2_and_U3 ( .A(cell_1875_a_HPC2_and_n7), .B(
        cell_1875_a_HPC2_and_z_0__0_), .ZN(cell_1875_and_out[0]) );
  XNOR2_X1 cell_1875_a_HPC2_and_U2 ( .A(
        cell_1875_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1875_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1875_a_HPC2_and_n7) );
  DFF_X1 cell_1875_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1875_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1875_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1875_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1875_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1875_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1875_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1875_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1875_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1875_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1876_U4 ( .A(n367), .B(cell_1876_and_out[1]), .Z(signal_3582)
         );
  XOR2_X1 cell_1876_U3 ( .A(n366), .B(cell_1876_and_out[0]), .Z(signal_2144)
         );
  XOR2_X1 cell_1876_U2 ( .A(n367), .B(signal_3406), .Z(cell_1876_and_in[1]) );
  XOR2_X1 cell_1876_U1 ( .A(n366), .B(signal_1992), .Z(cell_1876_and_in[0]) );
  XOR2_X1 cell_1876_a_HPC2_and_U14 ( .A(Fresh[162]), .B(cell_1876_and_in[0]), 
        .Z(cell_1876_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1876_a_HPC2_and_U13 ( .A(Fresh[162]), .B(cell_1876_and_in[1]), 
        .Z(cell_1876_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1876_a_HPC2_and_U12 ( .A1(cell_1876_a_HPC2_and_a_reg[1]), .A2(
        cell_1876_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1876_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1876_a_HPC2_and_U11 ( .A1(cell_1876_a_HPC2_and_a_reg[0]), .A2(
        cell_1876_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1876_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1876_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1876_a_HPC2_and_n9), 
        .ZN(cell_1876_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1876_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1876_a_HPC2_and_n9), 
        .ZN(cell_1876_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1876_a_HPC2_and_U8 ( .A(Fresh[162]), .ZN(cell_1876_a_HPC2_and_n9) );
  AND2_X1 cell_1876_a_HPC2_and_U7 ( .A1(cell_1876_and_in[1]), .A2(n425), .ZN(
        cell_1876_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1876_a_HPC2_and_U6 ( .A1(cell_1876_and_in[0]), .A2(n408), .ZN(
        cell_1876_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1876_a_HPC2_and_U5 ( .A(cell_1876_a_HPC2_and_n8), .B(
        cell_1876_a_HPC2_and_z_1__1_), .ZN(cell_1876_and_out[1]) );
  XNOR2_X1 cell_1876_a_HPC2_and_U4 ( .A(
        cell_1876_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1876_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1876_a_HPC2_and_n8) );
  XNOR2_X1 cell_1876_a_HPC2_and_U3 ( .A(cell_1876_a_HPC2_and_n7), .B(
        cell_1876_a_HPC2_and_z_0__0_), .ZN(cell_1876_and_out[0]) );
  XNOR2_X1 cell_1876_a_HPC2_and_U2 ( .A(
        cell_1876_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1876_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1876_a_HPC2_and_n7) );
  DFF_X1 cell_1876_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1876_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1876_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1876_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1876_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1876_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1876_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1876_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1876_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1876_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1877_U4 ( .A(signal_3406), .B(cell_1877_and_out[1]), .Z(
        signal_3583) );
  XOR2_X1 cell_1877_U3 ( .A(signal_1992), .B(cell_1877_and_out[0]), .Z(
        signal_2145) );
  XOR2_X1 cell_1877_U2 ( .A(signal_3406), .B(n360), .Z(cell_1877_and_in[1]) );
  XOR2_X1 cell_1877_U1 ( .A(signal_1992), .B(n358), .Z(cell_1877_and_in[0]) );
  XOR2_X1 cell_1877_a_HPC2_and_U14 ( .A(Fresh[163]), .B(cell_1877_and_in[0]), 
        .Z(cell_1877_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1877_a_HPC2_and_U13 ( .A(Fresh[163]), .B(cell_1877_and_in[1]), 
        .Z(cell_1877_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1877_a_HPC2_and_U12 ( .A1(cell_1877_a_HPC2_and_a_reg[1]), .A2(
        cell_1877_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1877_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1877_a_HPC2_and_U11 ( .A1(cell_1877_a_HPC2_and_a_reg[0]), .A2(
        cell_1877_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1877_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1877_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1877_a_HPC2_and_n9), 
        .ZN(cell_1877_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1877_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1877_a_HPC2_and_n9), 
        .ZN(cell_1877_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1877_a_HPC2_and_U8 ( .A(Fresh[163]), .ZN(cell_1877_a_HPC2_and_n9) );
  AND2_X1 cell_1877_a_HPC2_and_U7 ( .A1(cell_1877_and_in[1]), .A2(n425), .ZN(
        cell_1877_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1877_a_HPC2_and_U6 ( .A1(cell_1877_and_in[0]), .A2(n408), .ZN(
        cell_1877_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1877_a_HPC2_and_U5 ( .A(cell_1877_a_HPC2_and_n8), .B(
        cell_1877_a_HPC2_and_z_1__1_), .ZN(cell_1877_and_out[1]) );
  XNOR2_X1 cell_1877_a_HPC2_and_U4 ( .A(
        cell_1877_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1877_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1877_a_HPC2_and_n8) );
  XNOR2_X1 cell_1877_a_HPC2_and_U3 ( .A(cell_1877_a_HPC2_and_n7), .B(
        cell_1877_a_HPC2_and_z_0__0_), .ZN(cell_1877_and_out[0]) );
  XNOR2_X1 cell_1877_a_HPC2_and_U2 ( .A(
        cell_1877_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1877_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1877_a_HPC2_and_n7) );
  DFF_X1 cell_1877_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1877_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1877_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1877_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1877_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1877_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1877_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1877_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1877_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1877_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1878_U4 ( .A(n379), .B(cell_1878_and_out[1]), .Z(signal_3584)
         );
  XOR2_X1 cell_1878_U3 ( .A(n377), .B(cell_1878_and_out[0]), .Z(signal_2146)
         );
  XOR2_X1 cell_1878_U2 ( .A(n379), .B(n355), .Z(cell_1878_and_in[1]) );
  XOR2_X1 cell_1878_U1 ( .A(n377), .B(n353), .Z(cell_1878_and_in[0]) );
  XOR2_X1 cell_1878_a_HPC2_and_U14 ( .A(Fresh[164]), .B(cell_1878_and_in[0]), 
        .Z(cell_1878_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1878_a_HPC2_and_U13 ( .A(Fresh[164]), .B(cell_1878_and_in[1]), 
        .Z(cell_1878_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1878_a_HPC2_and_U12 ( .A1(cell_1878_a_HPC2_and_a_reg[1]), .A2(
        cell_1878_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1878_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1878_a_HPC2_and_U11 ( .A1(cell_1878_a_HPC2_and_a_reg[0]), .A2(
        cell_1878_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1878_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1878_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1878_a_HPC2_and_n9), 
        .ZN(cell_1878_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1878_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1878_a_HPC2_and_n9), 
        .ZN(cell_1878_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1878_a_HPC2_and_U8 ( .A(Fresh[164]), .ZN(cell_1878_a_HPC2_and_n9) );
  AND2_X1 cell_1878_a_HPC2_and_U7 ( .A1(cell_1878_and_in[1]), .A2(n425), .ZN(
        cell_1878_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1878_a_HPC2_and_U6 ( .A1(cell_1878_and_in[0]), .A2(n408), .ZN(
        cell_1878_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1878_a_HPC2_and_U5 ( .A(cell_1878_a_HPC2_and_n8), .B(
        cell_1878_a_HPC2_and_z_1__1_), .ZN(cell_1878_and_out[1]) );
  XNOR2_X1 cell_1878_a_HPC2_and_U4 ( .A(
        cell_1878_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1878_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1878_a_HPC2_and_n8) );
  XNOR2_X1 cell_1878_a_HPC2_and_U3 ( .A(cell_1878_a_HPC2_and_n7), .B(
        cell_1878_a_HPC2_and_z_0__0_), .ZN(cell_1878_and_out[0]) );
  XNOR2_X1 cell_1878_a_HPC2_and_U2 ( .A(
        cell_1878_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1878_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1878_a_HPC2_and_n7) );
  DFF_X1 cell_1878_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1878_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1878_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1878_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1878_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1878_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1878_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1878_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1878_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1878_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1879_U4 ( .A(n354), .B(cell_1879_and_out[1]), .Z(signal_3585)
         );
  XOR2_X1 cell_1879_U3 ( .A(n352), .B(cell_1879_and_out[0]), .Z(signal_2147)
         );
  XOR2_X1 cell_1879_U2 ( .A(n354), .B(1'b0), .Z(cell_1879_and_in[1]) );
  XOR2_X1 cell_1879_U1 ( .A(n352), .B(1'b1), .Z(cell_1879_and_in[0]) );
  XOR2_X1 cell_1879_a_HPC2_and_U14 ( .A(Fresh[165]), .B(cell_1879_and_in[0]), 
        .Z(cell_1879_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1879_a_HPC2_and_U13 ( .A(Fresh[165]), .B(cell_1879_and_in[1]), 
        .Z(cell_1879_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1879_a_HPC2_and_U12 ( .A1(cell_1879_a_HPC2_and_a_reg[1]), .A2(
        cell_1879_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1879_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1879_a_HPC2_and_U11 ( .A1(cell_1879_a_HPC2_and_a_reg[0]), .A2(
        cell_1879_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1879_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1879_a_HPC2_and_U10 ( .A1(n424), .A2(cell_1879_a_HPC2_and_n9), 
        .ZN(cell_1879_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1879_a_HPC2_and_U9 ( .A1(n407), .A2(cell_1879_a_HPC2_and_n9), 
        .ZN(cell_1879_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1879_a_HPC2_and_U8 ( .A(Fresh[165]), .ZN(cell_1879_a_HPC2_and_n9) );
  AND2_X1 cell_1879_a_HPC2_and_U7 ( .A1(cell_1879_and_in[1]), .A2(n424), .ZN(
        cell_1879_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1879_a_HPC2_and_U6 ( .A1(cell_1879_and_in[0]), .A2(n407), .ZN(
        cell_1879_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1879_a_HPC2_and_U5 ( .A(cell_1879_a_HPC2_and_n8), .B(
        cell_1879_a_HPC2_and_z_1__1_), .ZN(cell_1879_and_out[1]) );
  XNOR2_X1 cell_1879_a_HPC2_and_U4 ( .A(
        cell_1879_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1879_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1879_a_HPC2_and_n8) );
  XNOR2_X1 cell_1879_a_HPC2_and_U3 ( .A(cell_1879_a_HPC2_and_n7), .B(
        cell_1879_a_HPC2_and_z_0__0_), .ZN(cell_1879_and_out[0]) );
  XNOR2_X1 cell_1879_a_HPC2_and_U2 ( .A(
        cell_1879_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1879_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1879_a_HPC2_and_n7) );
  DFF_X1 cell_1879_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1879_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1879_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n407), .CK(clk), 
        .Q(cell_1879_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1879_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1879_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n424), .CK(clk), 
        .Q(cell_1879_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1879_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1879_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1879_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1880_U4 ( .A(n360), .B(cell_1880_and_out[1]), .Z(signal_3586)
         );
  XOR2_X1 cell_1880_U3 ( .A(n358), .B(cell_1880_and_out[0]), .Z(signal_2148)
         );
  XOR2_X1 cell_1880_U2 ( .A(n360), .B(n371), .Z(cell_1880_and_in[1]) );
  XOR2_X1 cell_1880_U1 ( .A(n358), .B(n369), .Z(cell_1880_and_in[0]) );
  XOR2_X1 cell_1880_a_HPC2_and_U14 ( .A(Fresh[166]), .B(cell_1880_and_in[0]), 
        .Z(cell_1880_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1880_a_HPC2_and_U13 ( .A(Fresh[166]), .B(cell_1880_and_in[1]), 
        .Z(cell_1880_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1880_a_HPC2_and_U12 ( .A1(cell_1880_a_HPC2_and_a_reg[1]), .A2(
        cell_1880_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1880_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1880_a_HPC2_and_U11 ( .A1(cell_1880_a_HPC2_and_a_reg[0]), .A2(
        cell_1880_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1880_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1880_a_HPC2_and_U10 ( .A1(n425), .A2(cell_1880_a_HPC2_and_n9), 
        .ZN(cell_1880_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1880_a_HPC2_and_U9 ( .A1(n408), .A2(cell_1880_a_HPC2_and_n9), 
        .ZN(cell_1880_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1880_a_HPC2_and_U8 ( .A(Fresh[166]), .ZN(cell_1880_a_HPC2_and_n9) );
  AND2_X1 cell_1880_a_HPC2_and_U7 ( .A1(cell_1880_and_in[1]), .A2(n425), .ZN(
        cell_1880_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1880_a_HPC2_and_U6 ( .A1(cell_1880_and_in[0]), .A2(n408), .ZN(
        cell_1880_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1880_a_HPC2_and_U5 ( .A(cell_1880_a_HPC2_and_n8), .B(
        cell_1880_a_HPC2_and_z_1__1_), .ZN(cell_1880_and_out[1]) );
  XNOR2_X1 cell_1880_a_HPC2_and_U4 ( .A(
        cell_1880_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1880_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1880_a_HPC2_and_n8) );
  XNOR2_X1 cell_1880_a_HPC2_and_U3 ( .A(cell_1880_a_HPC2_and_n7), .B(
        cell_1880_a_HPC2_and_z_0__0_), .ZN(cell_1880_and_out[0]) );
  XNOR2_X1 cell_1880_a_HPC2_and_U2 ( .A(
        cell_1880_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1880_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1880_a_HPC2_and_n7) );
  DFF_X1 cell_1880_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1880_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1880_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n408), .CK(clk), 
        .Q(cell_1880_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1880_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1880_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n425), .CK(clk), 
        .Q(cell_1880_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1880_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1880_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1880_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1881_U4 ( .A(1'b0), .B(cell_1881_and_out[1]), .Z(signal_3587)
         );
  XOR2_X1 cell_1881_U3 ( .A(1'b1), .B(cell_1881_and_out[0]), .Z(signal_2149)
         );
  XOR2_X1 cell_1881_U2 ( .A(1'b0), .B(n367), .Z(cell_1881_and_in[1]) );
  XOR2_X1 cell_1881_U1 ( .A(1'b1), .B(n366), .Z(cell_1881_and_in[0]) );
  XOR2_X1 cell_1881_a_HPC2_and_U14 ( .A(Fresh[167]), .B(cell_1881_and_in[0]), 
        .Z(cell_1881_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1881_a_HPC2_and_U13 ( .A(Fresh[167]), .B(cell_1881_and_in[1]), 
        .Z(cell_1881_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1881_a_HPC2_and_U12 ( .A1(cell_1881_a_HPC2_and_a_reg[1]), .A2(
        cell_1881_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1881_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1881_a_HPC2_and_U11 ( .A1(cell_1881_a_HPC2_and_a_reg[0]), .A2(
        cell_1881_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1881_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1881_a_HPC2_and_U10 ( .A1(n412), .A2(cell_1881_a_HPC2_and_n9), 
        .ZN(cell_1881_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1881_a_HPC2_and_U9 ( .A1(n395), .A2(cell_1881_a_HPC2_and_n9), 
        .ZN(cell_1881_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1881_a_HPC2_and_U8 ( .A(Fresh[167]), .ZN(cell_1881_a_HPC2_and_n9) );
  AND2_X1 cell_1881_a_HPC2_and_U7 ( .A1(cell_1881_and_in[1]), .A2(n412), .ZN(
        cell_1881_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1881_a_HPC2_and_U6 ( .A1(cell_1881_and_in[0]), .A2(n395), .ZN(
        cell_1881_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1881_a_HPC2_and_U5 ( .A(cell_1881_a_HPC2_and_n8), .B(
        cell_1881_a_HPC2_and_z_1__1_), .ZN(cell_1881_and_out[1]) );
  XNOR2_X1 cell_1881_a_HPC2_and_U4 ( .A(
        cell_1881_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1881_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1881_a_HPC2_and_n8) );
  XNOR2_X1 cell_1881_a_HPC2_and_U3 ( .A(cell_1881_a_HPC2_and_n7), .B(
        cell_1881_a_HPC2_and_z_0__0_), .ZN(cell_1881_and_out[0]) );
  XNOR2_X1 cell_1881_a_HPC2_and_U2 ( .A(
        cell_1881_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1881_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1881_a_HPC2_and_n7) );
  DFF_X1 cell_1881_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1881_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1881_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n395), .CK(clk), 
        .Q(cell_1881_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1881_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1881_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n412), .CK(clk), 
        .Q(cell_1881_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1881_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1881_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1881_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1882_U4 ( .A(n375), .B(cell_1882_and_out[1]), .Z(signal_3588)
         );
  XOR2_X1 cell_1882_U3 ( .A(n373), .B(cell_1882_and_out[0]), .Z(signal_2150)
         );
  XOR2_X1 cell_1882_U2 ( .A(n375), .B(1'b0), .Z(cell_1882_and_in[1]) );
  XOR2_X1 cell_1882_U1 ( .A(n373), .B(1'b0), .Z(cell_1882_and_in[0]) );
  XOR2_X1 cell_1882_a_HPC2_and_U14 ( .A(Fresh[168]), .B(cell_1882_and_in[0]), 
        .Z(cell_1882_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1882_a_HPC2_and_U13 ( .A(Fresh[168]), .B(cell_1882_and_in[1]), 
        .Z(cell_1882_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1882_a_HPC2_and_U12 ( .A1(cell_1882_a_HPC2_and_a_reg[1]), .A2(
        cell_1882_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1882_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1882_a_HPC2_and_U11 ( .A1(cell_1882_a_HPC2_and_a_reg[0]), .A2(
        cell_1882_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1882_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1882_a_HPC2_and_U10 ( .A1(n427), .A2(cell_1882_a_HPC2_and_n9), 
        .ZN(cell_1882_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1882_a_HPC2_and_U9 ( .A1(n410), .A2(cell_1882_a_HPC2_and_n9), 
        .ZN(cell_1882_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1882_a_HPC2_and_U8 ( .A(Fresh[168]), .ZN(cell_1882_a_HPC2_and_n9) );
  AND2_X1 cell_1882_a_HPC2_and_U7 ( .A1(cell_1882_and_in[1]), .A2(n427), .ZN(
        cell_1882_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1882_a_HPC2_and_U6 ( .A1(cell_1882_and_in[0]), .A2(n410), .ZN(
        cell_1882_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1882_a_HPC2_and_U5 ( .A(cell_1882_a_HPC2_and_n8), .B(
        cell_1882_a_HPC2_and_z_1__1_), .ZN(cell_1882_and_out[1]) );
  XNOR2_X1 cell_1882_a_HPC2_and_U4 ( .A(
        cell_1882_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1882_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1882_a_HPC2_and_n8) );
  XNOR2_X1 cell_1882_a_HPC2_and_U3 ( .A(cell_1882_a_HPC2_and_n7), .B(
        cell_1882_a_HPC2_and_z_0__0_), .ZN(cell_1882_and_out[0]) );
  XNOR2_X1 cell_1882_a_HPC2_and_U2 ( .A(
        cell_1882_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1882_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1882_a_HPC2_and_n7) );
  DFF_X1 cell_1882_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1882_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1882_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n410), .CK(clk), 
        .Q(cell_1882_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1882_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1882_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n427), .CK(clk), 
        .Q(cell_1882_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1882_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1882_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1882_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1883_U4 ( .A(n378), .B(cell_1883_and_out[1]), .Z(signal_3589)
         );
  XOR2_X1 cell_1883_U3 ( .A(n376), .B(cell_1883_and_out[0]), .Z(signal_2151)
         );
  XOR2_X1 cell_1883_U2 ( .A(n378), .B(n383), .Z(cell_1883_and_in[1]) );
  XOR2_X1 cell_1883_U1 ( .A(n376), .B(n382), .Z(cell_1883_and_in[0]) );
  XOR2_X1 cell_1883_a_HPC2_and_U14 ( .A(Fresh[169]), .B(cell_1883_and_in[0]), 
        .Z(cell_1883_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1883_a_HPC2_and_U13 ( .A(Fresh[169]), .B(cell_1883_and_in[1]), 
        .Z(cell_1883_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1883_a_HPC2_and_U12 ( .A1(cell_1883_a_HPC2_and_a_reg[1]), .A2(
        cell_1883_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1883_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1883_a_HPC2_and_U11 ( .A1(cell_1883_a_HPC2_and_a_reg[0]), .A2(
        cell_1883_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1883_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1883_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1883_a_HPC2_and_n9), 
        .ZN(cell_1883_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1883_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1883_a_HPC2_and_n9), 
        .ZN(cell_1883_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1883_a_HPC2_and_U8 ( .A(Fresh[169]), .ZN(cell_1883_a_HPC2_and_n9) );
  AND2_X1 cell_1883_a_HPC2_and_U7 ( .A1(cell_1883_and_in[1]), .A2(n426), .ZN(
        cell_1883_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1883_a_HPC2_and_U6 ( .A1(cell_1883_and_in[0]), .A2(n409), .ZN(
        cell_1883_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1883_a_HPC2_and_U5 ( .A(cell_1883_a_HPC2_and_n8), .B(
        cell_1883_a_HPC2_and_z_1__1_), .ZN(cell_1883_and_out[1]) );
  XNOR2_X1 cell_1883_a_HPC2_and_U4 ( .A(
        cell_1883_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1883_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1883_a_HPC2_and_n8) );
  XNOR2_X1 cell_1883_a_HPC2_and_U3 ( .A(cell_1883_a_HPC2_and_n7), .B(
        cell_1883_a_HPC2_and_z_0__0_), .ZN(cell_1883_and_out[0]) );
  XNOR2_X1 cell_1883_a_HPC2_and_U2 ( .A(
        cell_1883_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1883_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1883_a_HPC2_and_n7) );
  DFF_X1 cell_1883_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1883_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1883_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1883_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1883_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1883_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1883_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1883_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1883_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1883_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1884_U4 ( .A(n367), .B(cell_1884_and_out[1]), .Z(signal_3590)
         );
  XOR2_X1 cell_1884_U3 ( .A(n366), .B(cell_1884_and_out[0]), .Z(signal_2152)
         );
  XOR2_X1 cell_1884_U2 ( .A(n367), .B(n375), .Z(cell_1884_and_in[1]) );
  XOR2_X1 cell_1884_U1 ( .A(n366), .B(n373), .Z(cell_1884_and_in[0]) );
  XOR2_X1 cell_1884_a_HPC2_and_U14 ( .A(Fresh[170]), .B(cell_1884_and_in[0]), 
        .Z(cell_1884_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1884_a_HPC2_and_U13 ( .A(Fresh[170]), .B(cell_1884_and_in[1]), 
        .Z(cell_1884_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1884_a_HPC2_and_U12 ( .A1(cell_1884_a_HPC2_and_a_reg[1]), .A2(
        cell_1884_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1884_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1884_a_HPC2_and_U11 ( .A1(cell_1884_a_HPC2_and_a_reg[0]), .A2(
        cell_1884_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1884_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1884_a_HPC2_and_U10 ( .A1(n426), .A2(cell_1884_a_HPC2_and_n9), 
        .ZN(cell_1884_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1884_a_HPC2_and_U9 ( .A1(n409), .A2(cell_1884_a_HPC2_and_n9), 
        .ZN(cell_1884_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1884_a_HPC2_and_U8 ( .A(Fresh[170]), .ZN(cell_1884_a_HPC2_and_n9) );
  AND2_X1 cell_1884_a_HPC2_and_U7 ( .A1(cell_1884_and_in[1]), .A2(n426), .ZN(
        cell_1884_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1884_a_HPC2_and_U6 ( .A1(cell_1884_and_in[0]), .A2(n409), .ZN(
        cell_1884_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1884_a_HPC2_and_U5 ( .A(cell_1884_a_HPC2_and_n8), .B(
        cell_1884_a_HPC2_and_z_1__1_), .ZN(cell_1884_and_out[1]) );
  XNOR2_X1 cell_1884_a_HPC2_and_U4 ( .A(
        cell_1884_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1884_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1884_a_HPC2_and_n8) );
  XNOR2_X1 cell_1884_a_HPC2_and_U3 ( .A(cell_1884_a_HPC2_and_n7), .B(
        cell_1884_a_HPC2_and_z_0__0_), .ZN(cell_1884_and_out[0]) );
  XNOR2_X1 cell_1884_a_HPC2_and_U2 ( .A(
        cell_1884_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1884_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1884_a_HPC2_and_n7) );
  DFF_X1 cell_1884_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1884_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1884_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n409), .CK(clk), 
        .Q(cell_1884_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1884_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1884_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n426), .CK(clk), 
        .Q(cell_1884_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1884_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1884_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1884_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1885_U4 ( .A(signal_3462), .B(cell_1885_and_out[1]), .Z(
        signal_3663) );
  XOR2_X1 cell_1885_U3 ( .A(signal_2024), .B(cell_1885_and_out[0]), .Z(
        signal_2153) );
  XOR2_X1 cell_1885_U2 ( .A(signal_3462), .B(signal_3468), .Z(
        cell_1885_and_in[1]) );
  XOR2_X1 cell_1885_U1 ( .A(signal_2024), .B(signal_2030), .Z(
        cell_1885_and_in[0]) );
  XOR2_X1 cell_1885_a_HPC2_and_U14 ( .A(Fresh[171]), .B(cell_1885_and_in[0]), 
        .Z(cell_1885_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1885_a_HPC2_and_U13 ( .A(Fresh[171]), .B(cell_1885_and_in[1]), 
        .Z(cell_1885_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1885_a_HPC2_and_U12 ( .A1(cell_1885_a_HPC2_and_a_reg[1]), .A2(
        cell_1885_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1885_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1885_a_HPC2_and_U11 ( .A1(cell_1885_a_HPC2_and_a_reg[0]), .A2(
        cell_1885_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1885_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1885_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1885_a_HPC2_and_n9), 
        .ZN(cell_1885_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1885_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1885_a_HPC2_and_n9), 
        .ZN(cell_1885_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1885_a_HPC2_and_U8 ( .A(Fresh[171]), .ZN(cell_1885_a_HPC2_and_n9) );
  AND2_X1 cell_1885_a_HPC2_and_U7 ( .A1(cell_1885_and_in[1]), .A2(n451), .ZN(
        cell_1885_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1885_a_HPC2_and_U6 ( .A1(cell_1885_and_in[0]), .A2(n437), .ZN(
        cell_1885_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1885_a_HPC2_and_U5 ( .A(cell_1885_a_HPC2_and_n8), .B(
        cell_1885_a_HPC2_and_z_1__1_), .ZN(cell_1885_and_out[1]) );
  XNOR2_X1 cell_1885_a_HPC2_and_U4 ( .A(
        cell_1885_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1885_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1885_a_HPC2_and_n8) );
  XNOR2_X1 cell_1885_a_HPC2_and_U3 ( .A(cell_1885_a_HPC2_and_n7), .B(
        cell_1885_a_HPC2_and_z_0__0_), .ZN(cell_1885_and_out[0]) );
  XNOR2_X1 cell_1885_a_HPC2_and_U2 ( .A(
        cell_1885_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1885_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1885_a_HPC2_and_n7) );
  DFF_X1 cell_1885_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1885_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1885_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1885_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1885_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1885_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1885_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1885_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1885_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1885_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1886_U4 ( .A(signal_3569), .B(cell_1886_and_out[1]), .Z(
        signal_3664) );
  XOR2_X1 cell_1886_U3 ( .A(signal_2131), .B(cell_1886_and_out[0]), .Z(
        signal_2154) );
  XOR2_X1 cell_1886_U2 ( .A(signal_3569), .B(signal_3425), .Z(
        cell_1886_and_in[1]) );
  XOR2_X1 cell_1886_U1 ( .A(signal_2131), .B(signal_2011), .Z(
        cell_1886_and_in[0]) );
  XOR2_X1 cell_1886_a_HPC2_and_U14 ( .A(Fresh[172]), .B(cell_1886_and_in[0]), 
        .Z(cell_1886_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1886_a_HPC2_and_U13 ( .A(Fresh[172]), .B(cell_1886_and_in[1]), 
        .Z(cell_1886_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1886_a_HPC2_and_U12 ( .A1(cell_1886_a_HPC2_and_a_reg[1]), .A2(
        cell_1886_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1886_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1886_a_HPC2_and_U11 ( .A1(cell_1886_a_HPC2_and_a_reg[0]), .A2(
        cell_1886_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1886_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1886_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1886_a_HPC2_and_n9), 
        .ZN(cell_1886_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1886_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1886_a_HPC2_and_n9), 
        .ZN(cell_1886_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1886_a_HPC2_and_U8 ( .A(Fresh[172]), .ZN(cell_1886_a_HPC2_and_n9) );
  AND2_X1 cell_1886_a_HPC2_and_U7 ( .A1(cell_1886_and_in[1]), .A2(n442), .ZN(
        cell_1886_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1886_a_HPC2_and_U6 ( .A1(cell_1886_and_in[0]), .A2(n428), .ZN(
        cell_1886_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1886_a_HPC2_and_U5 ( .A(cell_1886_a_HPC2_and_n8), .B(
        cell_1886_a_HPC2_and_z_1__1_), .ZN(cell_1886_and_out[1]) );
  XNOR2_X1 cell_1886_a_HPC2_and_U4 ( .A(
        cell_1886_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1886_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1886_a_HPC2_and_n8) );
  XNOR2_X1 cell_1886_a_HPC2_and_U3 ( .A(cell_1886_a_HPC2_and_n7), .B(
        cell_1886_a_HPC2_and_z_0__0_), .ZN(cell_1886_and_out[0]) );
  XNOR2_X1 cell_1886_a_HPC2_and_U2 ( .A(
        cell_1886_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1886_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1886_a_HPC2_and_n7) );
  DFF_X1 cell_1886_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1886_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1886_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1886_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1886_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1886_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1886_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1886_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1886_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1886_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1887_U4 ( .A(signal_3549), .B(cell_1887_and_out[1]), .Z(
        signal_3665) );
  XOR2_X1 cell_1887_U3 ( .A(signal_2111), .B(cell_1887_and_out[0]), .Z(
        signal_2155) );
  XOR2_X1 cell_1887_U2 ( .A(signal_3549), .B(signal_3422), .Z(
        cell_1887_and_in[1]) );
  XOR2_X1 cell_1887_U1 ( .A(signal_2111), .B(signal_2008), .Z(
        cell_1887_and_in[0]) );
  XOR2_X1 cell_1887_a_HPC2_and_U14 ( .A(Fresh[173]), .B(cell_1887_and_in[0]), 
        .Z(cell_1887_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1887_a_HPC2_and_U13 ( .A(Fresh[173]), .B(cell_1887_and_in[1]), 
        .Z(cell_1887_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1887_a_HPC2_and_U12 ( .A1(cell_1887_a_HPC2_and_a_reg[1]), .A2(
        cell_1887_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1887_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1887_a_HPC2_and_U11 ( .A1(cell_1887_a_HPC2_and_a_reg[0]), .A2(
        cell_1887_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1887_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1887_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1887_a_HPC2_and_n9), 
        .ZN(cell_1887_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1887_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1887_a_HPC2_and_n9), 
        .ZN(cell_1887_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1887_a_HPC2_and_U8 ( .A(Fresh[173]), .ZN(cell_1887_a_HPC2_and_n9) );
  AND2_X1 cell_1887_a_HPC2_and_U7 ( .A1(cell_1887_and_in[1]), .A2(n442), .ZN(
        cell_1887_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1887_a_HPC2_and_U6 ( .A1(cell_1887_and_in[0]), .A2(n428), .ZN(
        cell_1887_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1887_a_HPC2_and_U5 ( .A(cell_1887_a_HPC2_and_n8), .B(
        cell_1887_a_HPC2_and_z_1__1_), .ZN(cell_1887_and_out[1]) );
  XNOR2_X1 cell_1887_a_HPC2_and_U4 ( .A(
        cell_1887_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1887_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1887_a_HPC2_and_n8) );
  XNOR2_X1 cell_1887_a_HPC2_and_U3 ( .A(cell_1887_a_HPC2_and_n7), .B(
        cell_1887_a_HPC2_and_z_0__0_), .ZN(cell_1887_and_out[0]) );
  XNOR2_X1 cell_1887_a_HPC2_and_U2 ( .A(
        cell_1887_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1887_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1887_a_HPC2_and_n7) );
  DFF_X1 cell_1887_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1887_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1887_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1887_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1887_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1887_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1887_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1887_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1887_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1887_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1888_U4 ( .A(signal_3517), .B(cell_1888_and_out[1]), .Z(
        signal_3666) );
  XOR2_X1 cell_1888_U3 ( .A(signal_2079), .B(cell_1888_and_out[0]), .Z(
        signal_2156) );
  XOR2_X1 cell_1888_U2 ( .A(signal_3517), .B(signal_3510), .Z(
        cell_1888_and_in[1]) );
  XOR2_X1 cell_1888_U1 ( .A(signal_2079), .B(signal_2072), .Z(
        cell_1888_and_in[0]) );
  XOR2_X1 cell_1888_a_HPC2_and_U14 ( .A(Fresh[174]), .B(cell_1888_and_in[0]), 
        .Z(cell_1888_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1888_a_HPC2_and_U13 ( .A(Fresh[174]), .B(cell_1888_and_in[1]), 
        .Z(cell_1888_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1888_a_HPC2_and_U12 ( .A1(cell_1888_a_HPC2_and_a_reg[1]), .A2(
        cell_1888_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1888_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1888_a_HPC2_and_U11 ( .A1(cell_1888_a_HPC2_and_a_reg[0]), .A2(
        cell_1888_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1888_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1888_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1888_a_HPC2_and_n9), 
        .ZN(cell_1888_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1888_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1888_a_HPC2_and_n9), 
        .ZN(cell_1888_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1888_a_HPC2_and_U8 ( .A(Fresh[174]), .ZN(cell_1888_a_HPC2_and_n9) );
  AND2_X1 cell_1888_a_HPC2_and_U7 ( .A1(cell_1888_and_in[1]), .A2(n442), .ZN(
        cell_1888_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1888_a_HPC2_and_U6 ( .A1(cell_1888_and_in[0]), .A2(n428), .ZN(
        cell_1888_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1888_a_HPC2_and_U5 ( .A(cell_1888_a_HPC2_and_n8), .B(
        cell_1888_a_HPC2_and_z_1__1_), .ZN(cell_1888_and_out[1]) );
  XNOR2_X1 cell_1888_a_HPC2_and_U4 ( .A(
        cell_1888_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1888_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1888_a_HPC2_and_n8) );
  XNOR2_X1 cell_1888_a_HPC2_and_U3 ( .A(cell_1888_a_HPC2_and_n7), .B(
        cell_1888_a_HPC2_and_z_0__0_), .ZN(cell_1888_and_out[0]) );
  XNOR2_X1 cell_1888_a_HPC2_and_U2 ( .A(
        cell_1888_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1888_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1888_a_HPC2_and_n7) );
  DFF_X1 cell_1888_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1888_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1888_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1888_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1888_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1888_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1888_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1888_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1888_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1888_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1889_U4 ( .A(signal_3491), .B(cell_1889_and_out[1]), .Z(
        signal_3667) );
  XOR2_X1 cell_1889_U3 ( .A(signal_2053), .B(cell_1889_and_out[0]), .Z(
        signal_2157) );
  XOR2_X1 cell_1889_U2 ( .A(signal_3491), .B(signal_3405), .Z(
        cell_1889_and_in[1]) );
  XOR2_X1 cell_1889_U1 ( .A(signal_2053), .B(signal_1991), .Z(
        cell_1889_and_in[0]) );
  XOR2_X1 cell_1889_a_HPC2_and_U14 ( .A(Fresh[175]), .B(cell_1889_and_in[0]), 
        .Z(cell_1889_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1889_a_HPC2_and_U13 ( .A(Fresh[175]), .B(cell_1889_and_in[1]), 
        .Z(cell_1889_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1889_a_HPC2_and_U12 ( .A1(cell_1889_a_HPC2_and_a_reg[1]), .A2(
        cell_1889_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1889_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1889_a_HPC2_and_U11 ( .A1(cell_1889_a_HPC2_and_a_reg[0]), .A2(
        cell_1889_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1889_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1889_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1889_a_HPC2_and_n9), 
        .ZN(cell_1889_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1889_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1889_a_HPC2_and_n9), 
        .ZN(cell_1889_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1889_a_HPC2_and_U8 ( .A(Fresh[175]), .ZN(cell_1889_a_HPC2_and_n9) );
  AND2_X1 cell_1889_a_HPC2_and_U7 ( .A1(cell_1889_and_in[1]), .A2(n443), .ZN(
        cell_1889_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1889_a_HPC2_and_U6 ( .A1(cell_1889_and_in[0]), .A2(n429), .ZN(
        cell_1889_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1889_a_HPC2_and_U5 ( .A(cell_1889_a_HPC2_and_n8), .B(
        cell_1889_a_HPC2_and_z_1__1_), .ZN(cell_1889_and_out[1]) );
  XNOR2_X1 cell_1889_a_HPC2_and_U4 ( .A(
        cell_1889_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1889_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1889_a_HPC2_and_n8) );
  XNOR2_X1 cell_1889_a_HPC2_and_U3 ( .A(cell_1889_a_HPC2_and_n7), .B(
        cell_1889_a_HPC2_and_z_0__0_), .ZN(cell_1889_and_out[0]) );
  XNOR2_X1 cell_1889_a_HPC2_and_U2 ( .A(
        cell_1889_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1889_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1889_a_HPC2_and_n7) );
  DFF_X1 cell_1889_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1889_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1889_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1889_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1889_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1889_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1889_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1889_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1889_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1889_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1890_U4 ( .A(signal_3538), .B(cell_1890_and_out[1]), .Z(
        signal_3668) );
  XOR2_X1 cell_1890_U3 ( .A(signal_2100), .B(cell_1890_and_out[0]), .Z(
        signal_2158) );
  XOR2_X1 cell_1890_U2 ( .A(signal_3538), .B(signal_3563), .Z(
        cell_1890_and_in[1]) );
  XOR2_X1 cell_1890_U1 ( .A(signal_2100), .B(signal_2125), .Z(
        cell_1890_and_in[0]) );
  XOR2_X1 cell_1890_a_HPC2_and_U14 ( .A(Fresh[176]), .B(cell_1890_and_in[0]), 
        .Z(cell_1890_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1890_a_HPC2_and_U13 ( .A(Fresh[176]), .B(cell_1890_and_in[1]), 
        .Z(cell_1890_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1890_a_HPC2_and_U12 ( .A1(cell_1890_a_HPC2_and_a_reg[1]), .A2(
        cell_1890_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1890_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1890_a_HPC2_and_U11 ( .A1(cell_1890_a_HPC2_and_a_reg[0]), .A2(
        cell_1890_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1890_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1890_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1890_a_HPC2_and_n9), 
        .ZN(cell_1890_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1890_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1890_a_HPC2_and_n9), 
        .ZN(cell_1890_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1890_a_HPC2_and_U8 ( .A(Fresh[176]), .ZN(cell_1890_a_HPC2_and_n9) );
  AND2_X1 cell_1890_a_HPC2_and_U7 ( .A1(cell_1890_and_in[1]), .A2(n443), .ZN(
        cell_1890_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1890_a_HPC2_and_U6 ( .A1(cell_1890_and_in[0]), .A2(n429), .ZN(
        cell_1890_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1890_a_HPC2_and_U5 ( .A(cell_1890_a_HPC2_and_n8), .B(
        cell_1890_a_HPC2_and_z_1__1_), .ZN(cell_1890_and_out[1]) );
  XNOR2_X1 cell_1890_a_HPC2_and_U4 ( .A(
        cell_1890_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1890_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1890_a_HPC2_and_n8) );
  XNOR2_X1 cell_1890_a_HPC2_and_U3 ( .A(cell_1890_a_HPC2_and_n7), .B(
        cell_1890_a_HPC2_and_z_0__0_), .ZN(cell_1890_and_out[0]) );
  XNOR2_X1 cell_1890_a_HPC2_and_U2 ( .A(
        cell_1890_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1890_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1890_a_HPC2_and_n7) );
  DFF_X1 cell_1890_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1890_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1890_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1890_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1890_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1890_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1890_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1890_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1890_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1890_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1891_U4 ( .A(signal_3521), .B(cell_1891_and_out[1]), .Z(
        signal_3669) );
  XOR2_X1 cell_1891_U3 ( .A(signal_2083), .B(cell_1891_and_out[0]), .Z(
        signal_2159) );
  XOR2_X1 cell_1891_U2 ( .A(signal_3521), .B(signal_3420), .Z(
        cell_1891_and_in[1]) );
  XOR2_X1 cell_1891_U1 ( .A(signal_2083), .B(signal_2006), .Z(
        cell_1891_and_in[0]) );
  XOR2_X1 cell_1891_a_HPC2_and_U14 ( .A(Fresh[177]), .B(cell_1891_and_in[0]), 
        .Z(cell_1891_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1891_a_HPC2_and_U13 ( .A(Fresh[177]), .B(cell_1891_and_in[1]), 
        .Z(cell_1891_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1891_a_HPC2_and_U12 ( .A1(cell_1891_a_HPC2_and_a_reg[1]), .A2(
        cell_1891_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1891_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1891_a_HPC2_and_U11 ( .A1(cell_1891_a_HPC2_and_a_reg[0]), .A2(
        cell_1891_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1891_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1891_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1891_a_HPC2_and_n9), 
        .ZN(cell_1891_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1891_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1891_a_HPC2_and_n9), 
        .ZN(cell_1891_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1891_a_HPC2_and_U8 ( .A(Fresh[177]), .ZN(cell_1891_a_HPC2_and_n9) );
  AND2_X1 cell_1891_a_HPC2_and_U7 ( .A1(cell_1891_and_in[1]), .A2(n451), .ZN(
        cell_1891_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1891_a_HPC2_and_U6 ( .A1(cell_1891_and_in[0]), .A2(n437), .ZN(
        cell_1891_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1891_a_HPC2_and_U5 ( .A(cell_1891_a_HPC2_and_n8), .B(
        cell_1891_a_HPC2_and_z_1__1_), .ZN(cell_1891_and_out[1]) );
  XNOR2_X1 cell_1891_a_HPC2_and_U4 ( .A(
        cell_1891_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1891_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1891_a_HPC2_and_n8) );
  XNOR2_X1 cell_1891_a_HPC2_and_U3 ( .A(cell_1891_a_HPC2_and_n7), .B(
        cell_1891_a_HPC2_and_z_0__0_), .ZN(cell_1891_and_out[0]) );
  XNOR2_X1 cell_1891_a_HPC2_and_U2 ( .A(
        cell_1891_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1891_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1891_a_HPC2_and_n7) );
  DFF_X1 cell_1891_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1891_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1891_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1891_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1891_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1891_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1891_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1891_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1891_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1891_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1892_U4 ( .A(signal_3474), .B(cell_1892_and_out[1]), .Z(
        signal_3670) );
  XOR2_X1 cell_1892_U3 ( .A(signal_2036), .B(cell_1892_and_out[0]), .Z(
        signal_2160) );
  XOR2_X1 cell_1892_U2 ( .A(signal_3474), .B(signal_3417), .Z(
        cell_1892_and_in[1]) );
  XOR2_X1 cell_1892_U1 ( .A(signal_2036), .B(signal_2003), .Z(
        cell_1892_and_in[0]) );
  XOR2_X1 cell_1892_a_HPC2_and_U14 ( .A(Fresh[178]), .B(cell_1892_and_in[0]), 
        .Z(cell_1892_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1892_a_HPC2_and_U13 ( .A(Fresh[178]), .B(cell_1892_and_in[1]), 
        .Z(cell_1892_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1892_a_HPC2_and_U12 ( .A1(cell_1892_a_HPC2_and_a_reg[1]), .A2(
        cell_1892_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1892_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1892_a_HPC2_and_U11 ( .A1(cell_1892_a_HPC2_and_a_reg[0]), .A2(
        cell_1892_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1892_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1892_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1892_a_HPC2_and_n9), 
        .ZN(cell_1892_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1892_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1892_a_HPC2_and_n9), 
        .ZN(cell_1892_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1892_a_HPC2_and_U8 ( .A(Fresh[178]), .ZN(cell_1892_a_HPC2_and_n9) );
  AND2_X1 cell_1892_a_HPC2_and_U7 ( .A1(cell_1892_and_in[1]), .A2(n451), .ZN(
        cell_1892_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1892_a_HPC2_and_U6 ( .A1(cell_1892_and_in[0]), .A2(n437), .ZN(
        cell_1892_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1892_a_HPC2_and_U5 ( .A(cell_1892_a_HPC2_and_n8), .B(
        cell_1892_a_HPC2_and_z_1__1_), .ZN(cell_1892_and_out[1]) );
  XNOR2_X1 cell_1892_a_HPC2_and_U4 ( .A(
        cell_1892_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1892_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1892_a_HPC2_and_n8) );
  XNOR2_X1 cell_1892_a_HPC2_and_U3 ( .A(cell_1892_a_HPC2_and_n7), .B(
        cell_1892_a_HPC2_and_z_0__0_), .ZN(cell_1892_and_out[0]) );
  XNOR2_X1 cell_1892_a_HPC2_and_U2 ( .A(
        cell_1892_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1892_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1892_a_HPC2_and_n7) );
  DFF_X1 cell_1892_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1892_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1892_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1892_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1892_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1892_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1892_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1892_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1892_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1892_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1893_U4 ( .A(signal_3555), .B(cell_1893_and_out[1]), .Z(
        signal_3671) );
  XOR2_X1 cell_1893_U3 ( .A(signal_2117), .B(cell_1893_and_out[0]), .Z(
        signal_2161) );
  XOR2_X1 cell_1893_U2 ( .A(signal_3555), .B(signal_3546), .Z(
        cell_1893_and_in[1]) );
  XOR2_X1 cell_1893_U1 ( .A(signal_2117), .B(signal_2108), .Z(
        cell_1893_and_in[0]) );
  XOR2_X1 cell_1893_a_HPC2_and_U14 ( .A(Fresh[179]), .B(cell_1893_and_in[0]), 
        .Z(cell_1893_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1893_a_HPC2_and_U13 ( .A(Fresh[179]), .B(cell_1893_and_in[1]), 
        .Z(cell_1893_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1893_a_HPC2_and_U12 ( .A1(cell_1893_a_HPC2_and_a_reg[1]), .A2(
        cell_1893_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1893_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1893_a_HPC2_and_U11 ( .A1(cell_1893_a_HPC2_and_a_reg[0]), .A2(
        cell_1893_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1893_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1893_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1893_a_HPC2_and_n9), 
        .ZN(cell_1893_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1893_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1893_a_HPC2_and_n9), 
        .ZN(cell_1893_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1893_a_HPC2_and_U8 ( .A(Fresh[179]), .ZN(cell_1893_a_HPC2_and_n9) );
  AND2_X1 cell_1893_a_HPC2_and_U7 ( .A1(cell_1893_and_in[1]), .A2(n451), .ZN(
        cell_1893_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1893_a_HPC2_and_U6 ( .A1(cell_1893_and_in[0]), .A2(n437), .ZN(
        cell_1893_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1893_a_HPC2_and_U5 ( .A(cell_1893_a_HPC2_and_n8), .B(
        cell_1893_a_HPC2_and_z_1__1_), .ZN(cell_1893_and_out[1]) );
  XNOR2_X1 cell_1893_a_HPC2_and_U4 ( .A(
        cell_1893_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1893_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1893_a_HPC2_and_n8) );
  XNOR2_X1 cell_1893_a_HPC2_and_U3 ( .A(cell_1893_a_HPC2_and_n7), .B(
        cell_1893_a_HPC2_and_z_0__0_), .ZN(cell_1893_and_out[0]) );
  XNOR2_X1 cell_1893_a_HPC2_and_U2 ( .A(
        cell_1893_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1893_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1893_a_HPC2_and_n7) );
  DFF_X1 cell_1893_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1893_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1893_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1893_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1893_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1893_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1893_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1893_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1893_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1893_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1894_U4 ( .A(signal_3409), .B(cell_1894_and_out[1]), .Z(
        signal_3672) );
  XOR2_X1 cell_1894_U3 ( .A(signal_1995), .B(cell_1894_and_out[0]), .Z(
        signal_2162) );
  XOR2_X1 cell_1894_U2 ( .A(signal_3409), .B(signal_3578), .Z(
        cell_1894_and_in[1]) );
  XOR2_X1 cell_1894_U1 ( .A(signal_1995), .B(signal_2140), .Z(
        cell_1894_and_in[0]) );
  XOR2_X1 cell_1894_a_HPC2_and_U14 ( .A(Fresh[180]), .B(cell_1894_and_in[0]), 
        .Z(cell_1894_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1894_a_HPC2_and_U13 ( .A(Fresh[180]), .B(cell_1894_and_in[1]), 
        .Z(cell_1894_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1894_a_HPC2_and_U12 ( .A1(cell_1894_a_HPC2_and_a_reg[1]), .A2(
        cell_1894_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1894_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1894_a_HPC2_and_U11 ( .A1(cell_1894_a_HPC2_and_a_reg[0]), .A2(
        cell_1894_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1894_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1894_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1894_a_HPC2_and_n9), 
        .ZN(cell_1894_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1894_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1894_a_HPC2_and_n9), 
        .ZN(cell_1894_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1894_a_HPC2_and_U8 ( .A(Fresh[180]), .ZN(cell_1894_a_HPC2_and_n9) );
  AND2_X1 cell_1894_a_HPC2_and_U7 ( .A1(cell_1894_and_in[1]), .A2(n443), .ZN(
        cell_1894_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1894_a_HPC2_and_U6 ( .A1(cell_1894_and_in[0]), .A2(n429), .ZN(
        cell_1894_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1894_a_HPC2_and_U5 ( .A(cell_1894_a_HPC2_and_n8), .B(
        cell_1894_a_HPC2_and_z_1__1_), .ZN(cell_1894_and_out[1]) );
  XNOR2_X1 cell_1894_a_HPC2_and_U4 ( .A(
        cell_1894_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1894_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1894_a_HPC2_and_n8) );
  XNOR2_X1 cell_1894_a_HPC2_and_U3 ( .A(cell_1894_a_HPC2_and_n7), .B(
        cell_1894_a_HPC2_and_z_0__0_), .ZN(cell_1894_and_out[0]) );
  XNOR2_X1 cell_1894_a_HPC2_and_U2 ( .A(
        cell_1894_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1894_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1894_a_HPC2_and_n7) );
  DFF_X1 cell_1894_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1894_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1894_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1894_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1894_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1894_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1894_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1894_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1894_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1894_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1895_U4 ( .A(signal_3477), .B(cell_1895_and_out[1]), .Z(
        signal_3673) );
  XOR2_X1 cell_1895_U3 ( .A(signal_2039), .B(cell_1895_and_out[0]), .Z(
        signal_2163) );
  XOR2_X1 cell_1895_U2 ( .A(signal_3477), .B(signal_3495), .Z(
        cell_1895_and_in[1]) );
  XOR2_X1 cell_1895_U1 ( .A(signal_2039), .B(signal_2057), .Z(
        cell_1895_and_in[0]) );
  XOR2_X1 cell_1895_a_HPC2_and_U14 ( .A(Fresh[181]), .B(cell_1895_and_in[0]), 
        .Z(cell_1895_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1895_a_HPC2_and_U13 ( .A(Fresh[181]), .B(cell_1895_and_in[1]), 
        .Z(cell_1895_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1895_a_HPC2_and_U12 ( .A1(cell_1895_a_HPC2_and_a_reg[1]), .A2(
        cell_1895_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1895_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1895_a_HPC2_and_U11 ( .A1(cell_1895_a_HPC2_and_a_reg[0]), .A2(
        cell_1895_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1895_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1895_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1895_a_HPC2_and_n9), 
        .ZN(cell_1895_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1895_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1895_a_HPC2_and_n9), 
        .ZN(cell_1895_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1895_a_HPC2_and_U8 ( .A(Fresh[181]), .ZN(cell_1895_a_HPC2_and_n9) );
  AND2_X1 cell_1895_a_HPC2_and_U7 ( .A1(cell_1895_and_in[1]), .A2(n443), .ZN(
        cell_1895_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1895_a_HPC2_and_U6 ( .A1(cell_1895_and_in[0]), .A2(n429), .ZN(
        cell_1895_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1895_a_HPC2_and_U5 ( .A(cell_1895_a_HPC2_and_n8), .B(
        cell_1895_a_HPC2_and_z_1__1_), .ZN(cell_1895_and_out[1]) );
  XNOR2_X1 cell_1895_a_HPC2_and_U4 ( .A(
        cell_1895_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1895_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1895_a_HPC2_and_n8) );
  XNOR2_X1 cell_1895_a_HPC2_and_U3 ( .A(cell_1895_a_HPC2_and_n7), .B(
        cell_1895_a_HPC2_and_z_0__0_), .ZN(cell_1895_and_out[0]) );
  XNOR2_X1 cell_1895_a_HPC2_and_U2 ( .A(
        cell_1895_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1895_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1895_a_HPC2_and_n7) );
  DFF_X1 cell_1895_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1895_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1895_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1895_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1895_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1895_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1895_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1895_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1895_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1895_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1896_U4 ( .A(signal_3403), .B(cell_1896_and_out[1]), .Z(
        signal_3674) );
  XOR2_X1 cell_1896_U3 ( .A(signal_1989), .B(cell_1896_and_out[0]), .Z(
        signal_2164) );
  XOR2_X1 cell_1896_U2 ( .A(signal_3403), .B(signal_3582), .Z(
        cell_1896_and_in[1]) );
  XOR2_X1 cell_1896_U1 ( .A(signal_1989), .B(signal_2144), .Z(
        cell_1896_and_in[0]) );
  XOR2_X1 cell_1896_a_HPC2_and_U14 ( .A(Fresh[182]), .B(cell_1896_and_in[0]), 
        .Z(cell_1896_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1896_a_HPC2_and_U13 ( .A(Fresh[182]), .B(cell_1896_and_in[1]), 
        .Z(cell_1896_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1896_a_HPC2_and_U12 ( .A1(cell_1896_a_HPC2_and_a_reg[1]), .A2(
        cell_1896_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1896_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1896_a_HPC2_and_U11 ( .A1(cell_1896_a_HPC2_and_a_reg[0]), .A2(
        cell_1896_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1896_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1896_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1896_a_HPC2_and_n9), 
        .ZN(cell_1896_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1896_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1896_a_HPC2_and_n9), 
        .ZN(cell_1896_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1896_a_HPC2_and_U8 ( .A(Fresh[182]), .ZN(cell_1896_a_HPC2_and_n9) );
  AND2_X1 cell_1896_a_HPC2_and_U7 ( .A1(cell_1896_and_in[1]), .A2(n451), .ZN(
        cell_1896_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1896_a_HPC2_and_U6 ( .A1(cell_1896_and_in[0]), .A2(n437), .ZN(
        cell_1896_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1896_a_HPC2_and_U5 ( .A(cell_1896_a_HPC2_and_n8), .B(
        cell_1896_a_HPC2_and_z_1__1_), .ZN(cell_1896_and_out[1]) );
  XNOR2_X1 cell_1896_a_HPC2_and_U4 ( .A(
        cell_1896_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1896_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1896_a_HPC2_and_n8) );
  XNOR2_X1 cell_1896_a_HPC2_and_U3 ( .A(cell_1896_a_HPC2_and_n7), .B(
        cell_1896_a_HPC2_and_z_0__0_), .ZN(cell_1896_and_out[0]) );
  XNOR2_X1 cell_1896_a_HPC2_and_U2 ( .A(
        cell_1896_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1896_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1896_a_HPC2_and_n7) );
  DFF_X1 cell_1896_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1896_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1896_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1896_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1896_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1896_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1896_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1896_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1896_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1896_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1897_U4 ( .A(signal_3573), .B(cell_1897_and_out[1]), .Z(
        signal_3675) );
  XOR2_X1 cell_1897_U3 ( .A(signal_2135), .B(cell_1897_and_out[0]), .Z(
        signal_2165) );
  XOR2_X1 cell_1897_U2 ( .A(signal_3573), .B(signal_3567), .Z(
        cell_1897_and_in[1]) );
  XOR2_X1 cell_1897_U1 ( .A(signal_2135), .B(signal_2129), .Z(
        cell_1897_and_in[0]) );
  XOR2_X1 cell_1897_a_HPC2_and_U14 ( .A(Fresh[183]), .B(cell_1897_and_in[0]), 
        .Z(cell_1897_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1897_a_HPC2_and_U13 ( .A(Fresh[183]), .B(cell_1897_and_in[1]), 
        .Z(cell_1897_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1897_a_HPC2_and_U12 ( .A1(cell_1897_a_HPC2_and_a_reg[1]), .A2(
        cell_1897_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1897_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1897_a_HPC2_and_U11 ( .A1(cell_1897_a_HPC2_and_a_reg[0]), .A2(
        cell_1897_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1897_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1897_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1897_a_HPC2_and_n9), 
        .ZN(cell_1897_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1897_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1897_a_HPC2_and_n9), 
        .ZN(cell_1897_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1897_a_HPC2_and_U8 ( .A(Fresh[183]), .ZN(cell_1897_a_HPC2_and_n9) );
  AND2_X1 cell_1897_a_HPC2_and_U7 ( .A1(cell_1897_and_in[1]), .A2(n443), .ZN(
        cell_1897_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1897_a_HPC2_and_U6 ( .A1(cell_1897_and_in[0]), .A2(n429), .ZN(
        cell_1897_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1897_a_HPC2_and_U5 ( .A(cell_1897_a_HPC2_and_n8), .B(
        cell_1897_a_HPC2_and_z_1__1_), .ZN(cell_1897_and_out[1]) );
  XNOR2_X1 cell_1897_a_HPC2_and_U4 ( .A(
        cell_1897_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1897_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1897_a_HPC2_and_n8) );
  XNOR2_X1 cell_1897_a_HPC2_and_U3 ( .A(cell_1897_a_HPC2_and_n7), .B(
        cell_1897_a_HPC2_and_z_0__0_), .ZN(cell_1897_and_out[0]) );
  XNOR2_X1 cell_1897_a_HPC2_and_U2 ( .A(
        cell_1897_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1897_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1897_a_HPC2_and_n7) );
  DFF_X1 cell_1897_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1897_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1897_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1897_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1897_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1897_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1897_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1897_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1897_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1897_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1898_U4 ( .A(signal_3495), .B(cell_1898_and_out[1]), .Z(
        signal_3676) );
  XOR2_X1 cell_1898_U3 ( .A(signal_2057), .B(cell_1898_and_out[0]), .Z(
        signal_2166) );
  XOR2_X1 cell_1898_U2 ( .A(signal_3495), .B(signal_3470), .Z(
        cell_1898_and_in[1]) );
  XOR2_X1 cell_1898_U1 ( .A(signal_2057), .B(signal_2032), .Z(
        cell_1898_and_in[0]) );
  XOR2_X1 cell_1898_a_HPC2_and_U14 ( .A(Fresh[184]), .B(cell_1898_and_in[0]), 
        .Z(cell_1898_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1898_a_HPC2_and_U13 ( .A(Fresh[184]), .B(cell_1898_and_in[1]), 
        .Z(cell_1898_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1898_a_HPC2_and_U12 ( .A1(cell_1898_a_HPC2_and_a_reg[1]), .A2(
        cell_1898_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1898_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1898_a_HPC2_and_U11 ( .A1(cell_1898_a_HPC2_and_a_reg[0]), .A2(
        cell_1898_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1898_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1898_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1898_a_HPC2_and_n9), 
        .ZN(cell_1898_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1898_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1898_a_HPC2_and_n9), 
        .ZN(cell_1898_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1898_a_HPC2_and_U8 ( .A(Fresh[184]), .ZN(cell_1898_a_HPC2_and_n9) );
  AND2_X1 cell_1898_a_HPC2_and_U7 ( .A1(cell_1898_and_in[1]), .A2(n443), .ZN(
        cell_1898_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1898_a_HPC2_and_U6 ( .A1(cell_1898_and_in[0]), .A2(n429), .ZN(
        cell_1898_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1898_a_HPC2_and_U5 ( .A(cell_1898_a_HPC2_and_n8), .B(
        cell_1898_a_HPC2_and_z_1__1_), .ZN(cell_1898_and_out[1]) );
  XNOR2_X1 cell_1898_a_HPC2_and_U4 ( .A(
        cell_1898_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1898_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1898_a_HPC2_and_n8) );
  XNOR2_X1 cell_1898_a_HPC2_and_U3 ( .A(cell_1898_a_HPC2_and_n7), .B(
        cell_1898_a_HPC2_and_z_0__0_), .ZN(cell_1898_and_out[0]) );
  XNOR2_X1 cell_1898_a_HPC2_and_U2 ( .A(
        cell_1898_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1898_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1898_a_HPC2_and_n7) );
  DFF_X1 cell_1898_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1898_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1898_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1898_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1898_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1898_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1898_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1898_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1898_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1898_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1899_U4 ( .A(signal_3408), .B(cell_1899_and_out[1]), .Z(
        signal_3677) );
  XOR2_X1 cell_1899_U3 ( .A(signal_1994), .B(cell_1899_and_out[0]), .Z(
        signal_2167) );
  XOR2_X1 cell_1899_U2 ( .A(signal_3408), .B(signal_3529), .Z(
        cell_1899_and_in[1]) );
  XOR2_X1 cell_1899_U1 ( .A(signal_1994), .B(signal_2091), .Z(
        cell_1899_and_in[0]) );
  XOR2_X1 cell_1899_a_HPC2_and_U14 ( .A(Fresh[185]), .B(cell_1899_and_in[0]), 
        .Z(cell_1899_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1899_a_HPC2_and_U13 ( .A(Fresh[185]), .B(cell_1899_and_in[1]), 
        .Z(cell_1899_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1899_a_HPC2_and_U12 ( .A1(cell_1899_a_HPC2_and_a_reg[1]), .A2(
        cell_1899_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1899_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1899_a_HPC2_and_U11 ( .A1(cell_1899_a_HPC2_and_a_reg[0]), .A2(
        cell_1899_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1899_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1899_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1899_a_HPC2_and_n9), 
        .ZN(cell_1899_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1899_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1899_a_HPC2_and_n9), 
        .ZN(cell_1899_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1899_a_HPC2_and_U8 ( .A(Fresh[185]), .ZN(cell_1899_a_HPC2_and_n9) );
  AND2_X1 cell_1899_a_HPC2_and_U7 ( .A1(cell_1899_and_in[1]), .A2(n443), .ZN(
        cell_1899_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1899_a_HPC2_and_U6 ( .A1(cell_1899_and_in[0]), .A2(n429), .ZN(
        cell_1899_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1899_a_HPC2_and_U5 ( .A(cell_1899_a_HPC2_and_n8), .B(
        cell_1899_a_HPC2_and_z_1__1_), .ZN(cell_1899_and_out[1]) );
  XNOR2_X1 cell_1899_a_HPC2_and_U4 ( .A(
        cell_1899_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1899_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1899_a_HPC2_and_n8) );
  XNOR2_X1 cell_1899_a_HPC2_and_U3 ( .A(cell_1899_a_HPC2_and_n7), .B(
        cell_1899_a_HPC2_and_z_0__0_), .ZN(cell_1899_and_out[0]) );
  XNOR2_X1 cell_1899_a_HPC2_and_U2 ( .A(
        cell_1899_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1899_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1899_a_HPC2_and_n7) );
  DFF_X1 cell_1899_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1899_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1899_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1899_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1899_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1899_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1899_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1899_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1899_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1899_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1900_U4 ( .A(signal_3530), .B(cell_1900_and_out[1]), .Z(
        signal_3678) );
  XOR2_X1 cell_1900_U3 ( .A(signal_2092), .B(cell_1900_and_out[0]), .Z(
        signal_2168) );
  XOR2_X1 cell_1900_U2 ( .A(signal_3530), .B(signal_3525), .Z(
        cell_1900_and_in[1]) );
  XOR2_X1 cell_1900_U1 ( .A(signal_2092), .B(signal_2087), .Z(
        cell_1900_and_in[0]) );
  XOR2_X1 cell_1900_a_HPC2_and_U14 ( .A(Fresh[186]), .B(cell_1900_and_in[0]), 
        .Z(cell_1900_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1900_a_HPC2_and_U13 ( .A(Fresh[186]), .B(cell_1900_and_in[1]), 
        .Z(cell_1900_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1900_a_HPC2_and_U12 ( .A1(cell_1900_a_HPC2_and_a_reg[1]), .A2(
        cell_1900_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1900_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1900_a_HPC2_and_U11 ( .A1(cell_1900_a_HPC2_and_a_reg[0]), .A2(
        cell_1900_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1900_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1900_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1900_a_HPC2_and_n9), 
        .ZN(cell_1900_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1900_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1900_a_HPC2_and_n9), 
        .ZN(cell_1900_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1900_a_HPC2_and_U8 ( .A(Fresh[186]), .ZN(cell_1900_a_HPC2_and_n9) );
  AND2_X1 cell_1900_a_HPC2_and_U7 ( .A1(cell_1900_and_in[1]), .A2(n454), .ZN(
        cell_1900_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1900_a_HPC2_and_U6 ( .A1(cell_1900_and_in[0]), .A2(n440), .ZN(
        cell_1900_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1900_a_HPC2_and_U5 ( .A(cell_1900_a_HPC2_and_n8), .B(
        cell_1900_a_HPC2_and_z_1__1_), .ZN(cell_1900_and_out[1]) );
  XNOR2_X1 cell_1900_a_HPC2_and_U4 ( .A(
        cell_1900_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1900_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1900_a_HPC2_and_n8) );
  XNOR2_X1 cell_1900_a_HPC2_and_U3 ( .A(cell_1900_a_HPC2_and_n7), .B(
        cell_1900_a_HPC2_and_z_0__0_), .ZN(cell_1900_and_out[0]) );
  XNOR2_X1 cell_1900_a_HPC2_and_U2 ( .A(
        cell_1900_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1900_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1900_a_HPC2_and_n7) );
  DFF_X1 cell_1900_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1900_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1900_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1900_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1900_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1900_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1900_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1900_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1900_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1900_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1901_U4 ( .A(signal_3544), .B(cell_1901_and_out[1]), .Z(
        signal_3679) );
  XOR2_X1 cell_1901_U3 ( .A(signal_2106), .B(cell_1901_and_out[0]), .Z(
        signal_2169) );
  XOR2_X1 cell_1901_U2 ( .A(signal_3544), .B(signal_3574), .Z(
        cell_1901_and_in[1]) );
  XOR2_X1 cell_1901_U1 ( .A(signal_2106), .B(signal_2136), .Z(
        cell_1901_and_in[0]) );
  XOR2_X1 cell_1901_a_HPC2_and_U14 ( .A(Fresh[187]), .B(cell_1901_and_in[0]), 
        .Z(cell_1901_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1901_a_HPC2_and_U13 ( .A(Fresh[187]), .B(cell_1901_and_in[1]), 
        .Z(cell_1901_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1901_a_HPC2_and_U12 ( .A1(cell_1901_a_HPC2_and_a_reg[1]), .A2(
        cell_1901_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1901_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1901_a_HPC2_and_U11 ( .A1(cell_1901_a_HPC2_and_a_reg[0]), .A2(
        cell_1901_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1901_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1901_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1901_a_HPC2_and_n9), 
        .ZN(cell_1901_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1901_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1901_a_HPC2_and_n9), 
        .ZN(cell_1901_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1901_a_HPC2_and_U8 ( .A(Fresh[187]), .ZN(cell_1901_a_HPC2_and_n9) );
  AND2_X1 cell_1901_a_HPC2_and_U7 ( .A1(cell_1901_and_in[1]), .A2(n451), .ZN(
        cell_1901_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1901_a_HPC2_and_U6 ( .A1(cell_1901_and_in[0]), .A2(n437), .ZN(
        cell_1901_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1901_a_HPC2_and_U5 ( .A(cell_1901_a_HPC2_and_n8), .B(
        cell_1901_a_HPC2_and_z_1__1_), .ZN(cell_1901_and_out[1]) );
  XNOR2_X1 cell_1901_a_HPC2_and_U4 ( .A(
        cell_1901_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1901_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1901_a_HPC2_and_n8) );
  XNOR2_X1 cell_1901_a_HPC2_and_U3 ( .A(cell_1901_a_HPC2_and_n7), .B(
        cell_1901_a_HPC2_and_z_0__0_), .ZN(cell_1901_and_out[0]) );
  XNOR2_X1 cell_1901_a_HPC2_and_U2 ( .A(
        cell_1901_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1901_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1901_a_HPC2_and_n7) );
  DFF_X1 cell_1901_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1901_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1901_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1901_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1901_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1901_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1901_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1901_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1901_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1901_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1902_U4 ( .A(signal_3529), .B(cell_1902_and_out[1]), .Z(
        signal_3680) );
  XOR2_X1 cell_1902_U3 ( .A(signal_2091), .B(cell_1902_and_out[0]), .Z(
        signal_2170) );
  XOR2_X1 cell_1902_U2 ( .A(signal_3529), .B(signal_3458), .Z(
        cell_1902_and_in[1]) );
  XOR2_X1 cell_1902_U1 ( .A(signal_2091), .B(signal_2020), .Z(
        cell_1902_and_in[0]) );
  XOR2_X1 cell_1902_a_HPC2_and_U14 ( .A(Fresh[188]), .B(cell_1902_and_in[0]), 
        .Z(cell_1902_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1902_a_HPC2_and_U13 ( .A(Fresh[188]), .B(cell_1902_and_in[1]), 
        .Z(cell_1902_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1902_a_HPC2_and_U12 ( .A1(cell_1902_a_HPC2_and_a_reg[1]), .A2(
        cell_1902_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1902_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1902_a_HPC2_and_U11 ( .A1(cell_1902_a_HPC2_and_a_reg[0]), .A2(
        cell_1902_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1902_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1902_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1902_a_HPC2_and_n9), 
        .ZN(cell_1902_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1902_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1902_a_HPC2_and_n9), 
        .ZN(cell_1902_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1902_a_HPC2_and_U8 ( .A(Fresh[188]), .ZN(cell_1902_a_HPC2_and_n9) );
  AND2_X1 cell_1902_a_HPC2_and_U7 ( .A1(cell_1902_and_in[1]), .A2(n451), .ZN(
        cell_1902_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1902_a_HPC2_and_U6 ( .A1(cell_1902_and_in[0]), .A2(n437), .ZN(
        cell_1902_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1902_a_HPC2_and_U5 ( .A(cell_1902_a_HPC2_and_n8), .B(
        cell_1902_a_HPC2_and_z_1__1_), .ZN(cell_1902_and_out[1]) );
  XNOR2_X1 cell_1902_a_HPC2_and_U4 ( .A(
        cell_1902_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1902_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1902_a_HPC2_and_n8) );
  XNOR2_X1 cell_1902_a_HPC2_and_U3 ( .A(cell_1902_a_HPC2_and_n7), .B(
        cell_1902_a_HPC2_and_z_0__0_), .ZN(cell_1902_and_out[0]) );
  XNOR2_X1 cell_1902_a_HPC2_and_U2 ( .A(
        cell_1902_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1902_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1902_a_HPC2_and_n7) );
  DFF_X1 cell_1902_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1902_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1902_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1902_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1902_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1902_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1902_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1902_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1902_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1902_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1903_U4 ( .A(signal_3563), .B(cell_1903_and_out[1]), .Z(
        signal_3681) );
  XOR2_X1 cell_1903_U3 ( .A(signal_2125), .B(cell_1903_and_out[0]), .Z(
        signal_2171) );
  XOR2_X1 cell_1903_U2 ( .A(signal_3563), .B(signal_3547), .Z(
        cell_1903_and_in[1]) );
  XOR2_X1 cell_1903_U1 ( .A(signal_2125), .B(signal_2109), .Z(
        cell_1903_and_in[0]) );
  XOR2_X1 cell_1903_a_HPC2_and_U14 ( .A(Fresh[189]), .B(cell_1903_and_in[0]), 
        .Z(cell_1903_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1903_a_HPC2_and_U13 ( .A(Fresh[189]), .B(cell_1903_and_in[1]), 
        .Z(cell_1903_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1903_a_HPC2_and_U12 ( .A1(cell_1903_a_HPC2_and_a_reg[1]), .A2(
        cell_1903_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1903_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1903_a_HPC2_and_U11 ( .A1(cell_1903_a_HPC2_and_a_reg[0]), .A2(
        cell_1903_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1903_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1903_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1903_a_HPC2_and_n9), 
        .ZN(cell_1903_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1903_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1903_a_HPC2_and_n9), 
        .ZN(cell_1903_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1903_a_HPC2_and_U8 ( .A(Fresh[189]), .ZN(cell_1903_a_HPC2_and_n9) );
  AND2_X1 cell_1903_a_HPC2_and_U7 ( .A1(cell_1903_and_in[1]), .A2(n453), .ZN(
        cell_1903_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1903_a_HPC2_and_U6 ( .A1(cell_1903_and_in[0]), .A2(n439), .ZN(
        cell_1903_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1903_a_HPC2_and_U5 ( .A(cell_1903_a_HPC2_and_n8), .B(
        cell_1903_a_HPC2_and_z_1__1_), .ZN(cell_1903_and_out[1]) );
  XNOR2_X1 cell_1903_a_HPC2_and_U4 ( .A(
        cell_1903_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1903_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1903_a_HPC2_and_n8) );
  XNOR2_X1 cell_1903_a_HPC2_and_U3 ( .A(cell_1903_a_HPC2_and_n7), .B(
        cell_1903_a_HPC2_and_z_0__0_), .ZN(cell_1903_and_out[0]) );
  XNOR2_X1 cell_1903_a_HPC2_and_U2 ( .A(
        cell_1903_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1903_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1903_a_HPC2_and_n7) );
  DFF_X1 cell_1903_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1903_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1903_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1903_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1903_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1903_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1903_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1903_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1903_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1903_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1904_U4 ( .A(signal_3507), .B(cell_1904_and_out[1]), .Z(
        signal_3682) );
  XOR2_X1 cell_1904_U3 ( .A(signal_2069), .B(cell_1904_and_out[0]), .Z(
        signal_2172) );
  XOR2_X1 cell_1904_U2 ( .A(signal_3507), .B(signal_3484), .Z(
        cell_1904_and_in[1]) );
  XOR2_X1 cell_1904_U1 ( .A(signal_2069), .B(signal_2046), .Z(
        cell_1904_and_in[0]) );
  XOR2_X1 cell_1904_a_HPC2_and_U14 ( .A(Fresh[190]), .B(cell_1904_and_in[0]), 
        .Z(cell_1904_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1904_a_HPC2_and_U13 ( .A(Fresh[190]), .B(cell_1904_and_in[1]), 
        .Z(cell_1904_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1904_a_HPC2_and_U12 ( .A1(cell_1904_a_HPC2_and_a_reg[1]), .A2(
        cell_1904_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1904_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1904_a_HPC2_and_U11 ( .A1(cell_1904_a_HPC2_and_a_reg[0]), .A2(
        cell_1904_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1904_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1904_a_HPC2_and_U10 ( .A1(n455), .A2(cell_1904_a_HPC2_and_n9), 
        .ZN(cell_1904_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1904_a_HPC2_and_U9 ( .A1(n441), .A2(cell_1904_a_HPC2_and_n9), 
        .ZN(cell_1904_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1904_a_HPC2_and_U8 ( .A(Fresh[190]), .ZN(cell_1904_a_HPC2_and_n9) );
  AND2_X1 cell_1904_a_HPC2_and_U7 ( .A1(cell_1904_and_in[1]), .A2(n455), .ZN(
        cell_1904_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1904_a_HPC2_and_U6 ( .A1(cell_1904_and_in[0]), .A2(n441), .ZN(
        cell_1904_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1904_a_HPC2_and_U5 ( .A(cell_1904_a_HPC2_and_n8), .B(
        cell_1904_a_HPC2_and_z_1__1_), .ZN(cell_1904_and_out[1]) );
  XNOR2_X1 cell_1904_a_HPC2_and_U4 ( .A(
        cell_1904_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1904_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1904_a_HPC2_and_n8) );
  XNOR2_X1 cell_1904_a_HPC2_and_U3 ( .A(cell_1904_a_HPC2_and_n7), .B(
        cell_1904_a_HPC2_and_z_0__0_), .ZN(cell_1904_and_out[0]) );
  XNOR2_X1 cell_1904_a_HPC2_and_U2 ( .A(
        cell_1904_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1904_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1904_a_HPC2_and_n7) );
  DFF_X1 cell_1904_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1904_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1904_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_1904_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1904_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1904_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_1904_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1904_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1904_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1904_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1905_U4 ( .A(signal_3576), .B(cell_1905_and_out[1]), .Z(
        signal_3683) );
  XOR2_X1 cell_1905_U3 ( .A(signal_2138), .B(cell_1905_and_out[0]), .Z(
        signal_2173) );
  XOR2_X1 cell_1905_U2 ( .A(signal_3576), .B(signal_3480), .Z(
        cell_1905_and_in[1]) );
  XOR2_X1 cell_1905_U1 ( .A(signal_2138), .B(signal_2042), .Z(
        cell_1905_and_in[0]) );
  XOR2_X1 cell_1905_a_HPC2_and_U14 ( .A(Fresh[191]), .B(cell_1905_and_in[0]), 
        .Z(cell_1905_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1905_a_HPC2_and_U13 ( .A(Fresh[191]), .B(cell_1905_and_in[1]), 
        .Z(cell_1905_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1905_a_HPC2_and_U12 ( .A1(cell_1905_a_HPC2_and_a_reg[1]), .A2(
        cell_1905_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1905_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1905_a_HPC2_and_U11 ( .A1(cell_1905_a_HPC2_and_a_reg[0]), .A2(
        cell_1905_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1905_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1905_a_HPC2_and_U10 ( .A1(n455), .A2(cell_1905_a_HPC2_and_n9), 
        .ZN(cell_1905_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1905_a_HPC2_and_U9 ( .A1(n441), .A2(cell_1905_a_HPC2_and_n9), 
        .ZN(cell_1905_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1905_a_HPC2_and_U8 ( .A(Fresh[191]), .ZN(cell_1905_a_HPC2_and_n9) );
  AND2_X1 cell_1905_a_HPC2_and_U7 ( .A1(cell_1905_and_in[1]), .A2(n455), .ZN(
        cell_1905_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1905_a_HPC2_and_U6 ( .A1(cell_1905_and_in[0]), .A2(n441), .ZN(
        cell_1905_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1905_a_HPC2_and_U5 ( .A(cell_1905_a_HPC2_and_n8), .B(
        cell_1905_a_HPC2_and_z_1__1_), .ZN(cell_1905_and_out[1]) );
  XNOR2_X1 cell_1905_a_HPC2_and_U4 ( .A(
        cell_1905_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1905_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1905_a_HPC2_and_n8) );
  XNOR2_X1 cell_1905_a_HPC2_and_U3 ( .A(cell_1905_a_HPC2_and_n7), .B(
        cell_1905_a_HPC2_and_z_0__0_), .ZN(cell_1905_and_out[0]) );
  XNOR2_X1 cell_1905_a_HPC2_and_U2 ( .A(
        cell_1905_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1905_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1905_a_HPC2_and_n7) );
  DFF_X1 cell_1905_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1905_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1905_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_1905_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1905_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1905_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_1905_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1905_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1905_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1905_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1906_U4 ( .A(signal_3538), .B(cell_1906_and_out[1]), .Z(
        signal_3684) );
  XOR2_X1 cell_1906_U3 ( .A(signal_2100), .B(cell_1906_and_out[0]), .Z(
        signal_2174) );
  XOR2_X1 cell_1906_U2 ( .A(signal_3538), .B(signal_3542), .Z(
        cell_1906_and_in[1]) );
  XOR2_X1 cell_1906_U1 ( .A(signal_2100), .B(signal_2104), .Z(
        cell_1906_and_in[0]) );
  XOR2_X1 cell_1906_a_HPC2_and_U14 ( .A(Fresh[192]), .B(cell_1906_and_in[0]), 
        .Z(cell_1906_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1906_a_HPC2_and_U13 ( .A(Fresh[192]), .B(cell_1906_and_in[1]), 
        .Z(cell_1906_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1906_a_HPC2_and_U12 ( .A1(cell_1906_a_HPC2_and_a_reg[1]), .A2(
        cell_1906_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1906_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1906_a_HPC2_and_U11 ( .A1(cell_1906_a_HPC2_and_a_reg[0]), .A2(
        cell_1906_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1906_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1906_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1906_a_HPC2_and_n9), 
        .ZN(cell_1906_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1906_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1906_a_HPC2_and_n9), 
        .ZN(cell_1906_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1906_a_HPC2_and_U8 ( .A(Fresh[192]), .ZN(cell_1906_a_HPC2_and_n9) );
  AND2_X1 cell_1906_a_HPC2_and_U7 ( .A1(cell_1906_and_in[1]), .A2(n452), .ZN(
        cell_1906_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1906_a_HPC2_and_U6 ( .A1(cell_1906_and_in[0]), .A2(n438), .ZN(
        cell_1906_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1906_a_HPC2_and_U5 ( .A(cell_1906_a_HPC2_and_n8), .B(
        cell_1906_a_HPC2_and_z_1__1_), .ZN(cell_1906_and_out[1]) );
  XNOR2_X1 cell_1906_a_HPC2_and_U4 ( .A(
        cell_1906_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1906_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1906_a_HPC2_and_n8) );
  XNOR2_X1 cell_1906_a_HPC2_and_U3 ( .A(cell_1906_a_HPC2_and_n7), .B(
        cell_1906_a_HPC2_and_z_0__0_), .ZN(cell_1906_and_out[0]) );
  XNOR2_X1 cell_1906_a_HPC2_and_U2 ( .A(
        cell_1906_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1906_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1906_a_HPC2_and_n7) );
  DFF_X1 cell_1906_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1906_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1906_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1906_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1906_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1906_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1906_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1906_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1906_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1906_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1907_U4 ( .A(signal_3567), .B(cell_1907_and_out[1]), .Z(
        signal_3685) );
  XOR2_X1 cell_1907_U3 ( .A(signal_2129), .B(cell_1907_and_out[0]), .Z(
        signal_2175) );
  XOR2_X1 cell_1907_U2 ( .A(signal_3567), .B(signal_3474), .Z(
        cell_1907_and_in[1]) );
  XOR2_X1 cell_1907_U1 ( .A(signal_2129), .B(signal_2036), .Z(
        cell_1907_and_in[0]) );
  XOR2_X1 cell_1907_a_HPC2_and_U14 ( .A(Fresh[193]), .B(cell_1907_and_in[0]), 
        .Z(cell_1907_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1907_a_HPC2_and_U13 ( .A(Fresh[193]), .B(cell_1907_and_in[1]), 
        .Z(cell_1907_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1907_a_HPC2_and_U12 ( .A1(cell_1907_a_HPC2_and_a_reg[1]), .A2(
        cell_1907_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1907_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1907_a_HPC2_and_U11 ( .A1(cell_1907_a_HPC2_and_a_reg[0]), .A2(
        cell_1907_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1907_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1907_a_HPC2_and_U10 ( .A1(n455), .A2(cell_1907_a_HPC2_and_n9), 
        .ZN(cell_1907_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1907_a_HPC2_and_U9 ( .A1(n441), .A2(cell_1907_a_HPC2_and_n9), 
        .ZN(cell_1907_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1907_a_HPC2_and_U8 ( .A(Fresh[193]), .ZN(cell_1907_a_HPC2_and_n9) );
  AND2_X1 cell_1907_a_HPC2_and_U7 ( .A1(cell_1907_and_in[1]), .A2(n455), .ZN(
        cell_1907_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1907_a_HPC2_and_U6 ( .A1(cell_1907_and_in[0]), .A2(n441), .ZN(
        cell_1907_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1907_a_HPC2_and_U5 ( .A(cell_1907_a_HPC2_and_n8), .B(
        cell_1907_a_HPC2_and_z_1__1_), .ZN(cell_1907_and_out[1]) );
  XNOR2_X1 cell_1907_a_HPC2_and_U4 ( .A(
        cell_1907_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1907_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1907_a_HPC2_and_n8) );
  XNOR2_X1 cell_1907_a_HPC2_and_U3 ( .A(cell_1907_a_HPC2_and_n7), .B(
        cell_1907_a_HPC2_and_z_0__0_), .ZN(cell_1907_and_out[0]) );
  XNOR2_X1 cell_1907_a_HPC2_and_U2 ( .A(
        cell_1907_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1907_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1907_a_HPC2_and_n7) );
  DFF_X1 cell_1907_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1907_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1907_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_1907_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1907_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1907_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_1907_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1907_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1907_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1907_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1908_U4 ( .A(signal_3557), .B(cell_1908_and_out[1]), .Z(
        signal_3686) );
  XOR2_X1 cell_1908_U3 ( .A(signal_2119), .B(cell_1908_and_out[0]), .Z(
        signal_2176) );
  XOR2_X1 cell_1908_U2 ( .A(signal_3557), .B(signal_3586), .Z(
        cell_1908_and_in[1]) );
  XOR2_X1 cell_1908_U1 ( .A(signal_2119), .B(signal_2148), .Z(
        cell_1908_and_in[0]) );
  XOR2_X1 cell_1908_a_HPC2_and_U14 ( .A(Fresh[194]), .B(cell_1908_and_in[0]), 
        .Z(cell_1908_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1908_a_HPC2_and_U13 ( .A(Fresh[194]), .B(cell_1908_and_in[1]), 
        .Z(cell_1908_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1908_a_HPC2_and_U12 ( .A1(cell_1908_a_HPC2_and_a_reg[1]), .A2(
        cell_1908_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1908_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1908_a_HPC2_and_U11 ( .A1(cell_1908_a_HPC2_and_a_reg[0]), .A2(
        cell_1908_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1908_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1908_a_HPC2_and_U10 ( .A1(n455), .A2(cell_1908_a_HPC2_and_n9), 
        .ZN(cell_1908_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1908_a_HPC2_and_U9 ( .A1(n441), .A2(cell_1908_a_HPC2_and_n9), 
        .ZN(cell_1908_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1908_a_HPC2_and_U8 ( .A(Fresh[194]), .ZN(cell_1908_a_HPC2_and_n9) );
  AND2_X1 cell_1908_a_HPC2_and_U7 ( .A1(cell_1908_and_in[1]), .A2(n455), .ZN(
        cell_1908_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1908_a_HPC2_and_U6 ( .A1(cell_1908_and_in[0]), .A2(n441), .ZN(
        cell_1908_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1908_a_HPC2_and_U5 ( .A(cell_1908_a_HPC2_and_n8), .B(
        cell_1908_a_HPC2_and_z_1__1_), .ZN(cell_1908_and_out[1]) );
  XNOR2_X1 cell_1908_a_HPC2_and_U4 ( .A(
        cell_1908_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1908_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1908_a_HPC2_and_n8) );
  XNOR2_X1 cell_1908_a_HPC2_and_U3 ( .A(cell_1908_a_HPC2_and_n7), .B(
        cell_1908_a_HPC2_and_z_0__0_), .ZN(cell_1908_and_out[0]) );
  XNOR2_X1 cell_1908_a_HPC2_and_U2 ( .A(
        cell_1908_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1908_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1908_a_HPC2_and_n7) );
  DFF_X1 cell_1908_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1908_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1908_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_1908_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1908_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1908_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_1908_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1908_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1908_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1908_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1909_U4 ( .A(signal_3537), .B(cell_1909_and_out[1]), .Z(
        signal_3687) );
  XOR2_X1 cell_1909_U3 ( .A(signal_2099), .B(cell_1909_and_out[0]), .Z(
        signal_2177) );
  XOR2_X1 cell_1909_U2 ( .A(signal_3537), .B(signal_3472), .Z(
        cell_1909_and_in[1]) );
  XOR2_X1 cell_1909_U1 ( .A(signal_2099), .B(signal_2034), .Z(
        cell_1909_and_in[0]) );
  XOR2_X1 cell_1909_a_HPC2_and_U14 ( .A(Fresh[195]), .B(cell_1909_and_in[0]), 
        .Z(cell_1909_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1909_a_HPC2_and_U13 ( .A(Fresh[195]), .B(cell_1909_and_in[1]), 
        .Z(cell_1909_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1909_a_HPC2_and_U12 ( .A1(cell_1909_a_HPC2_and_a_reg[1]), .A2(
        cell_1909_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1909_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1909_a_HPC2_and_U11 ( .A1(cell_1909_a_HPC2_and_a_reg[0]), .A2(
        cell_1909_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1909_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1909_a_HPC2_and_U10 ( .A1(n455), .A2(cell_1909_a_HPC2_and_n9), 
        .ZN(cell_1909_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1909_a_HPC2_and_U9 ( .A1(n441), .A2(cell_1909_a_HPC2_and_n9), 
        .ZN(cell_1909_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1909_a_HPC2_and_U8 ( .A(Fresh[195]), .ZN(cell_1909_a_HPC2_and_n9) );
  AND2_X1 cell_1909_a_HPC2_and_U7 ( .A1(cell_1909_and_in[1]), .A2(n455), .ZN(
        cell_1909_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1909_a_HPC2_and_U6 ( .A1(cell_1909_and_in[0]), .A2(n441), .ZN(
        cell_1909_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1909_a_HPC2_and_U5 ( .A(cell_1909_a_HPC2_and_n8), .B(
        cell_1909_a_HPC2_and_z_1__1_), .ZN(cell_1909_and_out[1]) );
  XNOR2_X1 cell_1909_a_HPC2_and_U4 ( .A(
        cell_1909_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1909_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1909_a_HPC2_and_n8) );
  XNOR2_X1 cell_1909_a_HPC2_and_U3 ( .A(cell_1909_a_HPC2_and_n7), .B(
        cell_1909_a_HPC2_and_z_0__0_), .ZN(cell_1909_and_out[0]) );
  XNOR2_X1 cell_1909_a_HPC2_and_U2 ( .A(
        cell_1909_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1909_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1909_a_HPC2_and_n7) );
  DFF_X1 cell_1909_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1909_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1909_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_1909_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1909_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1909_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_1909_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1909_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1909_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1909_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1910_U4 ( .A(signal_3423), .B(cell_1910_and_out[1]), .Z(
        signal_3688) );
  XOR2_X1 cell_1910_U3 ( .A(signal_2009), .B(cell_1910_and_out[0]), .Z(
        signal_2178) );
  XOR2_X1 cell_1910_U2 ( .A(signal_3423), .B(signal_3485), .Z(
        cell_1910_and_in[1]) );
  XOR2_X1 cell_1910_U1 ( .A(signal_2009), .B(signal_2047), .Z(
        cell_1910_and_in[0]) );
  XOR2_X1 cell_1910_a_HPC2_and_U14 ( .A(Fresh[196]), .B(cell_1910_and_in[0]), 
        .Z(cell_1910_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1910_a_HPC2_and_U13 ( .A(Fresh[196]), .B(cell_1910_and_in[1]), 
        .Z(cell_1910_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1910_a_HPC2_and_U12 ( .A1(cell_1910_a_HPC2_and_a_reg[1]), .A2(
        cell_1910_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1910_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1910_a_HPC2_and_U11 ( .A1(cell_1910_a_HPC2_and_a_reg[0]), .A2(
        cell_1910_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1910_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1910_a_HPC2_and_U10 ( .A1(signal_3235), .A2(
        cell_1910_a_HPC2_and_n9), .ZN(cell_1910_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1910_a_HPC2_and_U9 ( .A1(signal_1514), .A2(
        cell_1910_a_HPC2_and_n9), .ZN(cell_1910_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1910_a_HPC2_and_U8 ( .A(Fresh[196]), .ZN(cell_1910_a_HPC2_and_n9) );
  AND2_X1 cell_1910_a_HPC2_and_U7 ( .A1(cell_1910_and_in[1]), .A2(signal_3235), 
        .ZN(cell_1910_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1910_a_HPC2_and_U6 ( .A1(cell_1910_and_in[0]), .A2(signal_1514), 
        .ZN(cell_1910_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1910_a_HPC2_and_U5 ( .A(cell_1910_a_HPC2_and_n8), .B(
        cell_1910_a_HPC2_and_z_1__1_), .ZN(cell_1910_and_out[1]) );
  XNOR2_X1 cell_1910_a_HPC2_and_U4 ( .A(
        cell_1910_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1910_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1910_a_HPC2_and_n8) );
  XNOR2_X1 cell_1910_a_HPC2_and_U3 ( .A(cell_1910_a_HPC2_and_n7), .B(
        cell_1910_a_HPC2_and_z_0__0_), .ZN(cell_1910_and_out[0]) );
  XNOR2_X1 cell_1910_a_HPC2_and_U2 ( .A(
        cell_1910_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1910_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1910_a_HPC2_and_n7) );
  DFF_X1 cell_1910_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1910_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1910_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1514), 
        .CK(clk), .Q(cell_1910_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1910_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1910_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3235), 
        .CK(clk), .Q(cell_1910_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1910_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1910_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1910_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1911_U4 ( .A(signal_3259), .B(cell_1911_and_out[1]), .Z(
        signal_3689) );
  XOR2_X1 cell_1911_U3 ( .A(signal_1985), .B(cell_1911_and_out[0]), .Z(
        signal_2179) );
  XOR2_X1 cell_1911_U2 ( .A(signal_3259), .B(signal_3560), .Z(
        cell_1911_and_in[1]) );
  XOR2_X1 cell_1911_U1 ( .A(signal_1985), .B(signal_2122), .Z(
        cell_1911_and_in[0]) );
  XOR2_X1 cell_1911_a_HPC2_and_U14 ( .A(Fresh[197]), .B(cell_1911_and_in[0]), 
        .Z(cell_1911_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1911_a_HPC2_and_U13 ( .A(Fresh[197]), .B(cell_1911_and_in[1]), 
        .Z(cell_1911_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1911_a_HPC2_and_U12 ( .A1(cell_1911_a_HPC2_and_a_reg[1]), .A2(
        cell_1911_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1911_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1911_a_HPC2_and_U11 ( .A1(cell_1911_a_HPC2_and_a_reg[0]), .A2(
        cell_1911_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1911_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1911_a_HPC2_and_U10 ( .A1(signal_3235), .A2(
        cell_1911_a_HPC2_and_n9), .ZN(cell_1911_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1911_a_HPC2_and_U9 ( .A1(signal_1514), .A2(
        cell_1911_a_HPC2_and_n9), .ZN(cell_1911_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1911_a_HPC2_and_U8 ( .A(Fresh[197]), .ZN(cell_1911_a_HPC2_and_n9) );
  AND2_X1 cell_1911_a_HPC2_and_U7 ( .A1(cell_1911_and_in[1]), .A2(signal_3235), 
        .ZN(cell_1911_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1911_a_HPC2_and_U6 ( .A1(cell_1911_and_in[0]), .A2(signal_1514), 
        .ZN(cell_1911_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1911_a_HPC2_and_U5 ( .A(cell_1911_a_HPC2_and_n8), .B(
        cell_1911_a_HPC2_and_z_1__1_), .ZN(cell_1911_and_out[1]) );
  XNOR2_X1 cell_1911_a_HPC2_and_U4 ( .A(
        cell_1911_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1911_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1911_a_HPC2_and_n8) );
  XNOR2_X1 cell_1911_a_HPC2_and_U3 ( .A(cell_1911_a_HPC2_and_n7), .B(
        cell_1911_a_HPC2_and_z_0__0_), .ZN(cell_1911_and_out[0]) );
  XNOR2_X1 cell_1911_a_HPC2_and_U2 ( .A(
        cell_1911_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1911_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1911_a_HPC2_and_n7) );
  DFF_X1 cell_1911_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1911_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1911_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1514), 
        .CK(clk), .Q(cell_1911_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1911_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1911_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3235), 
        .CK(clk), .Q(cell_1911_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1911_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1911_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1911_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1912_U4 ( .A(signal_3433), .B(cell_1912_and_out[1]), .Z(
        signal_3690) );
  XOR2_X1 cell_1912_U3 ( .A(signal_2019), .B(cell_1912_and_out[0]), .Z(
        signal_2180) );
  XOR2_X1 cell_1912_U2 ( .A(signal_3433), .B(signal_3588), .Z(
        cell_1912_and_in[1]) );
  XOR2_X1 cell_1912_U1 ( .A(signal_2019), .B(signal_2150), .Z(
        cell_1912_and_in[0]) );
  XOR2_X1 cell_1912_a_HPC2_and_U14 ( .A(Fresh[198]), .B(cell_1912_and_in[0]), 
        .Z(cell_1912_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1912_a_HPC2_and_U13 ( .A(Fresh[198]), .B(cell_1912_and_in[1]), 
        .Z(cell_1912_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1912_a_HPC2_and_U12 ( .A1(cell_1912_a_HPC2_and_a_reg[1]), .A2(
        cell_1912_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1912_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1912_a_HPC2_and_U11 ( .A1(cell_1912_a_HPC2_and_a_reg[0]), .A2(
        cell_1912_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1912_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1912_a_HPC2_and_U10 ( .A1(signal_3235), .A2(
        cell_1912_a_HPC2_and_n9), .ZN(cell_1912_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1912_a_HPC2_and_U9 ( .A1(signal_1514), .A2(
        cell_1912_a_HPC2_and_n9), .ZN(cell_1912_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1912_a_HPC2_and_U8 ( .A(Fresh[198]), .ZN(cell_1912_a_HPC2_and_n9) );
  AND2_X1 cell_1912_a_HPC2_and_U7 ( .A1(cell_1912_and_in[1]), .A2(signal_3235), 
        .ZN(cell_1912_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1912_a_HPC2_and_U6 ( .A1(cell_1912_and_in[0]), .A2(signal_1514), 
        .ZN(cell_1912_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1912_a_HPC2_and_U5 ( .A(cell_1912_a_HPC2_and_n8), .B(
        cell_1912_a_HPC2_and_z_1__1_), .ZN(cell_1912_and_out[1]) );
  XNOR2_X1 cell_1912_a_HPC2_and_U4 ( .A(
        cell_1912_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1912_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1912_a_HPC2_and_n8) );
  XNOR2_X1 cell_1912_a_HPC2_and_U3 ( .A(cell_1912_a_HPC2_and_n7), .B(
        cell_1912_a_HPC2_and_z_0__0_), .ZN(cell_1912_and_out[0]) );
  XNOR2_X1 cell_1912_a_HPC2_and_U2 ( .A(
        cell_1912_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1912_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1912_a_HPC2_and_n7) );
  DFF_X1 cell_1912_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1912_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1912_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1514), 
        .CK(clk), .Q(cell_1912_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1912_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1912_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3235), 
        .CK(clk), .Q(cell_1912_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1912_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1912_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1912_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1913_U4 ( .A(signal_3539), .B(cell_1913_and_out[1]), .Z(
        signal_3691) );
  XOR2_X1 cell_1913_U3 ( .A(signal_2101), .B(cell_1913_and_out[0]), .Z(
        signal_2181) );
  XOR2_X1 cell_1913_U2 ( .A(signal_3539), .B(signal_3588), .Z(
        cell_1913_and_in[1]) );
  XOR2_X1 cell_1913_U1 ( .A(signal_2101), .B(signal_2150), .Z(
        cell_1913_and_in[0]) );
  XOR2_X1 cell_1913_a_HPC2_and_U14 ( .A(Fresh[199]), .B(cell_1913_and_in[0]), 
        .Z(cell_1913_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1913_a_HPC2_and_U13 ( .A(Fresh[199]), .B(cell_1913_and_in[1]), 
        .Z(cell_1913_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1913_a_HPC2_and_U12 ( .A1(cell_1913_a_HPC2_and_a_reg[1]), .A2(
        cell_1913_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1913_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1913_a_HPC2_and_U11 ( .A1(cell_1913_a_HPC2_and_a_reg[0]), .A2(
        cell_1913_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1913_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1913_a_HPC2_and_U10 ( .A1(n455), .A2(cell_1913_a_HPC2_and_n9), 
        .ZN(cell_1913_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1913_a_HPC2_and_U9 ( .A1(n441), .A2(cell_1913_a_HPC2_and_n9), 
        .ZN(cell_1913_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1913_a_HPC2_and_U8 ( .A(Fresh[199]), .ZN(cell_1913_a_HPC2_and_n9) );
  AND2_X1 cell_1913_a_HPC2_and_U7 ( .A1(cell_1913_and_in[1]), .A2(n455), .ZN(
        cell_1913_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1913_a_HPC2_and_U6 ( .A1(cell_1913_and_in[0]), .A2(n441), .ZN(
        cell_1913_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1913_a_HPC2_and_U5 ( .A(cell_1913_a_HPC2_and_n8), .B(
        cell_1913_a_HPC2_and_z_1__1_), .ZN(cell_1913_and_out[1]) );
  XNOR2_X1 cell_1913_a_HPC2_and_U4 ( .A(
        cell_1913_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1913_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1913_a_HPC2_and_n8) );
  XNOR2_X1 cell_1913_a_HPC2_and_U3 ( .A(cell_1913_a_HPC2_and_n7), .B(
        cell_1913_a_HPC2_and_z_0__0_), .ZN(cell_1913_and_out[0]) );
  XNOR2_X1 cell_1913_a_HPC2_and_U2 ( .A(
        cell_1913_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1913_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1913_a_HPC2_and_n7) );
  DFF_X1 cell_1913_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1913_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1913_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_1913_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1913_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1913_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_1913_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1913_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1913_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1913_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1914_U4 ( .A(signal_3540), .B(cell_1914_and_out[1]), .Z(
        signal_3692) );
  XOR2_X1 cell_1914_U3 ( .A(signal_2102), .B(cell_1914_and_out[0]), .Z(
        signal_2182) );
  XOR2_X1 cell_1914_U2 ( .A(signal_3540), .B(signal_3494), .Z(
        cell_1914_and_in[1]) );
  XOR2_X1 cell_1914_U1 ( .A(signal_2102), .B(signal_2056), .Z(
        cell_1914_and_in[0]) );
  XOR2_X1 cell_1914_a_HPC2_and_U14 ( .A(Fresh[200]), .B(cell_1914_and_in[0]), 
        .Z(cell_1914_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1914_a_HPC2_and_U13 ( .A(Fresh[200]), .B(cell_1914_and_in[1]), 
        .Z(cell_1914_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1914_a_HPC2_and_U12 ( .A1(cell_1914_a_HPC2_and_a_reg[1]), .A2(
        cell_1914_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1914_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1914_a_HPC2_and_U11 ( .A1(cell_1914_a_HPC2_and_a_reg[0]), .A2(
        cell_1914_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1914_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1914_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1914_a_HPC2_and_n9), 
        .ZN(cell_1914_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1914_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1914_a_HPC2_and_n9), 
        .ZN(cell_1914_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1914_a_HPC2_and_U8 ( .A(Fresh[200]), .ZN(cell_1914_a_HPC2_and_n9) );
  AND2_X1 cell_1914_a_HPC2_and_U7 ( .A1(cell_1914_and_in[1]), .A2(n449), .ZN(
        cell_1914_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1914_a_HPC2_and_U6 ( .A1(cell_1914_and_in[0]), .A2(n435), .ZN(
        cell_1914_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1914_a_HPC2_and_U5 ( .A(cell_1914_a_HPC2_and_n8), .B(
        cell_1914_a_HPC2_and_z_1__1_), .ZN(cell_1914_and_out[1]) );
  XNOR2_X1 cell_1914_a_HPC2_and_U4 ( .A(
        cell_1914_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1914_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1914_a_HPC2_and_n8) );
  XNOR2_X1 cell_1914_a_HPC2_and_U3 ( .A(cell_1914_a_HPC2_and_n7), .B(
        cell_1914_a_HPC2_and_z_0__0_), .ZN(cell_1914_and_out[0]) );
  XNOR2_X1 cell_1914_a_HPC2_and_U2 ( .A(
        cell_1914_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1914_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1914_a_HPC2_and_n7) );
  DFF_X1 cell_1914_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1914_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1914_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1914_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1914_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1914_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1914_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1914_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1914_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1914_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1915_U4 ( .A(signal_3483), .B(cell_1915_and_out[1]), .Z(
        signal_3693) );
  XOR2_X1 cell_1915_U3 ( .A(signal_2045), .B(cell_1915_and_out[0]), .Z(
        signal_2183) );
  XOR2_X1 cell_1915_U2 ( .A(signal_3483), .B(signal_3470), .Z(
        cell_1915_and_in[1]) );
  XOR2_X1 cell_1915_U1 ( .A(signal_2045), .B(signal_2032), .Z(
        cell_1915_and_in[0]) );
  XOR2_X1 cell_1915_a_HPC2_and_U14 ( .A(Fresh[201]), .B(cell_1915_and_in[0]), 
        .Z(cell_1915_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1915_a_HPC2_and_U13 ( .A(Fresh[201]), .B(cell_1915_and_in[1]), 
        .Z(cell_1915_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1915_a_HPC2_and_U12 ( .A1(cell_1915_a_HPC2_and_a_reg[1]), .A2(
        cell_1915_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1915_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1915_a_HPC2_and_U11 ( .A1(cell_1915_a_HPC2_and_a_reg[0]), .A2(
        cell_1915_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1915_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1915_a_HPC2_and_U10 ( .A1(signal_3235), .A2(
        cell_1915_a_HPC2_and_n9), .ZN(cell_1915_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1915_a_HPC2_and_U9 ( .A1(signal_1514), .A2(
        cell_1915_a_HPC2_and_n9), .ZN(cell_1915_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1915_a_HPC2_and_U8 ( .A(Fresh[201]), .ZN(cell_1915_a_HPC2_and_n9) );
  AND2_X1 cell_1915_a_HPC2_and_U7 ( .A1(cell_1915_and_in[1]), .A2(signal_3235), 
        .ZN(cell_1915_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1915_a_HPC2_and_U6 ( .A1(cell_1915_and_in[0]), .A2(signal_1514), 
        .ZN(cell_1915_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1915_a_HPC2_and_U5 ( .A(cell_1915_a_HPC2_and_n8), .B(
        cell_1915_a_HPC2_and_z_1__1_), .ZN(cell_1915_and_out[1]) );
  XNOR2_X1 cell_1915_a_HPC2_and_U4 ( .A(
        cell_1915_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1915_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1915_a_HPC2_and_n8) );
  XNOR2_X1 cell_1915_a_HPC2_and_U3 ( .A(cell_1915_a_HPC2_and_n7), .B(
        cell_1915_a_HPC2_and_z_0__0_), .ZN(cell_1915_and_out[0]) );
  XNOR2_X1 cell_1915_a_HPC2_and_U2 ( .A(
        cell_1915_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1915_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1915_a_HPC2_and_n7) );
  DFF_X1 cell_1915_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1915_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1915_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1514), 
        .CK(clk), .Q(cell_1915_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1915_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1915_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3235), 
        .CK(clk), .Q(cell_1915_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1915_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1915_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1915_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1916_U4 ( .A(signal_3536), .B(cell_1916_and_out[1]), .Z(
        signal_3694) );
  XOR2_X1 cell_1916_U3 ( .A(signal_2098), .B(cell_1916_and_out[0]), .Z(
        signal_2184) );
  XOR2_X1 cell_1916_U2 ( .A(signal_3536), .B(signal_3528), .Z(
        cell_1916_and_in[1]) );
  XOR2_X1 cell_1916_U1 ( .A(signal_2098), .B(signal_2090), .Z(
        cell_1916_and_in[0]) );
  XOR2_X1 cell_1916_a_HPC2_and_U14 ( .A(Fresh[202]), .B(cell_1916_and_in[0]), 
        .Z(cell_1916_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1916_a_HPC2_and_U13 ( .A(Fresh[202]), .B(cell_1916_and_in[1]), 
        .Z(cell_1916_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1916_a_HPC2_and_U12 ( .A1(cell_1916_a_HPC2_and_a_reg[1]), .A2(
        cell_1916_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1916_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1916_a_HPC2_and_U11 ( .A1(cell_1916_a_HPC2_and_a_reg[0]), .A2(
        cell_1916_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1916_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1916_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1916_a_HPC2_and_n9), 
        .ZN(cell_1916_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1916_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1916_a_HPC2_and_n9), 
        .ZN(cell_1916_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1916_a_HPC2_and_U8 ( .A(Fresh[202]), .ZN(cell_1916_a_HPC2_and_n9) );
  AND2_X1 cell_1916_a_HPC2_and_U7 ( .A1(cell_1916_and_in[1]), .A2(n443), .ZN(
        cell_1916_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1916_a_HPC2_and_U6 ( .A1(cell_1916_and_in[0]), .A2(n429), .ZN(
        cell_1916_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1916_a_HPC2_and_U5 ( .A(cell_1916_a_HPC2_and_n8), .B(
        cell_1916_a_HPC2_and_z_1__1_), .ZN(cell_1916_and_out[1]) );
  XNOR2_X1 cell_1916_a_HPC2_and_U4 ( .A(
        cell_1916_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1916_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1916_a_HPC2_and_n8) );
  XNOR2_X1 cell_1916_a_HPC2_and_U3 ( .A(cell_1916_a_HPC2_and_n7), .B(
        cell_1916_a_HPC2_and_z_0__0_), .ZN(cell_1916_and_out[0]) );
  XNOR2_X1 cell_1916_a_HPC2_and_U2 ( .A(
        cell_1916_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1916_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1916_a_HPC2_and_n7) );
  DFF_X1 cell_1916_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1916_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1916_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1916_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1916_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1916_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1916_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1916_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1916_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1916_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1917_U4 ( .A(signal_3533), .B(cell_1917_and_out[1]), .Z(
        signal_3695) );
  XOR2_X1 cell_1917_U3 ( .A(signal_2095), .B(cell_1917_and_out[0]), .Z(
        signal_2185) );
  XOR2_X1 cell_1917_U2 ( .A(signal_3533), .B(signal_3479), .Z(
        cell_1917_and_in[1]) );
  XOR2_X1 cell_1917_U1 ( .A(signal_2095), .B(signal_2041), .Z(
        cell_1917_and_in[0]) );
  XOR2_X1 cell_1917_a_HPC2_and_U14 ( .A(Fresh[203]), .B(cell_1917_and_in[0]), 
        .Z(cell_1917_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1917_a_HPC2_and_U13 ( .A(Fresh[203]), .B(cell_1917_and_in[1]), 
        .Z(cell_1917_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1917_a_HPC2_and_U12 ( .A1(cell_1917_a_HPC2_and_a_reg[1]), .A2(
        cell_1917_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1917_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1917_a_HPC2_and_U11 ( .A1(cell_1917_a_HPC2_and_a_reg[0]), .A2(
        cell_1917_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1917_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1917_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1917_a_HPC2_and_n9), 
        .ZN(cell_1917_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1917_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1917_a_HPC2_and_n9), 
        .ZN(cell_1917_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1917_a_HPC2_and_U8 ( .A(Fresh[203]), .ZN(cell_1917_a_HPC2_and_n9) );
  AND2_X1 cell_1917_a_HPC2_and_U7 ( .A1(cell_1917_and_in[1]), .A2(n452), .ZN(
        cell_1917_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1917_a_HPC2_and_U6 ( .A1(cell_1917_and_in[0]), .A2(n438), .ZN(
        cell_1917_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1917_a_HPC2_and_U5 ( .A(cell_1917_a_HPC2_and_n8), .B(
        cell_1917_a_HPC2_and_z_1__1_), .ZN(cell_1917_and_out[1]) );
  XNOR2_X1 cell_1917_a_HPC2_and_U4 ( .A(
        cell_1917_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1917_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1917_a_HPC2_and_n8) );
  XNOR2_X1 cell_1917_a_HPC2_and_U3 ( .A(cell_1917_a_HPC2_and_n7), .B(
        cell_1917_a_HPC2_and_z_0__0_), .ZN(cell_1917_and_out[0]) );
  XNOR2_X1 cell_1917_a_HPC2_and_U2 ( .A(
        cell_1917_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1917_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1917_a_HPC2_and_n7) );
  DFF_X1 cell_1917_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1917_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1917_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1917_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1917_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1917_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1917_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1917_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1917_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1917_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1918_U4 ( .A(signal_3580), .B(cell_1918_and_out[1]), .Z(
        signal_3696) );
  XOR2_X1 cell_1918_U3 ( .A(signal_2142), .B(cell_1918_and_out[0]), .Z(
        signal_2186) );
  XOR2_X1 cell_1918_U2 ( .A(signal_3580), .B(signal_3508), .Z(
        cell_1918_and_in[1]) );
  XOR2_X1 cell_1918_U1 ( .A(signal_2142), .B(signal_2070), .Z(
        cell_1918_and_in[0]) );
  XOR2_X1 cell_1918_a_HPC2_and_U14 ( .A(Fresh[204]), .B(cell_1918_and_in[0]), 
        .Z(cell_1918_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1918_a_HPC2_and_U13 ( .A(Fresh[204]), .B(cell_1918_and_in[1]), 
        .Z(cell_1918_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1918_a_HPC2_and_U12 ( .A1(cell_1918_a_HPC2_and_a_reg[1]), .A2(
        cell_1918_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1918_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1918_a_HPC2_and_U11 ( .A1(cell_1918_a_HPC2_and_a_reg[0]), .A2(
        cell_1918_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1918_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1918_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1918_a_HPC2_and_n9), 
        .ZN(cell_1918_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1918_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1918_a_HPC2_and_n9), 
        .ZN(cell_1918_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1918_a_HPC2_and_U8 ( .A(Fresh[204]), .ZN(cell_1918_a_HPC2_and_n9) );
  AND2_X1 cell_1918_a_HPC2_and_U7 ( .A1(cell_1918_and_in[1]), .A2(n444), .ZN(
        cell_1918_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1918_a_HPC2_and_U6 ( .A1(cell_1918_and_in[0]), .A2(n430), .ZN(
        cell_1918_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1918_a_HPC2_and_U5 ( .A(cell_1918_a_HPC2_and_n8), .B(
        cell_1918_a_HPC2_and_z_1__1_), .ZN(cell_1918_and_out[1]) );
  XNOR2_X1 cell_1918_a_HPC2_and_U4 ( .A(
        cell_1918_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1918_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1918_a_HPC2_and_n8) );
  XNOR2_X1 cell_1918_a_HPC2_and_U3 ( .A(cell_1918_a_HPC2_and_n7), .B(
        cell_1918_a_HPC2_and_z_0__0_), .ZN(cell_1918_and_out[0]) );
  XNOR2_X1 cell_1918_a_HPC2_and_U2 ( .A(
        cell_1918_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1918_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1918_a_HPC2_and_n7) );
  DFF_X1 cell_1918_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1918_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1918_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1918_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1918_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1918_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1918_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1918_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1918_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1918_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1919_U4 ( .A(signal_3508), .B(cell_1919_and_out[1]), .Z(
        signal_3697) );
  XOR2_X1 cell_1919_U3 ( .A(signal_2070), .B(cell_1919_and_out[0]), .Z(
        signal_2187) );
  XOR2_X1 cell_1919_U2 ( .A(signal_3508), .B(signal_3570), .Z(
        cell_1919_and_in[1]) );
  XOR2_X1 cell_1919_U1 ( .A(signal_2070), .B(signal_2132), .Z(
        cell_1919_and_in[0]) );
  XOR2_X1 cell_1919_a_HPC2_and_U14 ( .A(Fresh[205]), .B(cell_1919_and_in[0]), 
        .Z(cell_1919_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1919_a_HPC2_and_U13 ( .A(Fresh[205]), .B(cell_1919_and_in[1]), 
        .Z(cell_1919_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1919_a_HPC2_and_U12 ( .A1(cell_1919_a_HPC2_and_a_reg[1]), .A2(
        cell_1919_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1919_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1919_a_HPC2_and_U11 ( .A1(cell_1919_a_HPC2_and_a_reg[0]), .A2(
        cell_1919_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1919_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1919_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1919_a_HPC2_and_n9), 
        .ZN(cell_1919_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1919_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1919_a_HPC2_and_n9), 
        .ZN(cell_1919_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1919_a_HPC2_and_U8 ( .A(Fresh[205]), .ZN(cell_1919_a_HPC2_and_n9) );
  AND2_X1 cell_1919_a_HPC2_and_U7 ( .A1(cell_1919_and_in[1]), .A2(n452), .ZN(
        cell_1919_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1919_a_HPC2_and_U6 ( .A1(cell_1919_and_in[0]), .A2(n438), .ZN(
        cell_1919_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1919_a_HPC2_and_U5 ( .A(cell_1919_a_HPC2_and_n8), .B(
        cell_1919_a_HPC2_and_z_1__1_), .ZN(cell_1919_and_out[1]) );
  XNOR2_X1 cell_1919_a_HPC2_and_U4 ( .A(
        cell_1919_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1919_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1919_a_HPC2_and_n8) );
  XNOR2_X1 cell_1919_a_HPC2_and_U3 ( .A(cell_1919_a_HPC2_and_n7), .B(
        cell_1919_a_HPC2_and_z_0__0_), .ZN(cell_1919_and_out[0]) );
  XNOR2_X1 cell_1919_a_HPC2_and_U2 ( .A(
        cell_1919_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1919_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1919_a_HPC2_and_n7) );
  DFF_X1 cell_1919_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1919_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1919_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1919_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1919_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1919_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1919_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1919_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1919_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1919_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1920_U4 ( .A(signal_3534), .B(cell_1920_and_out[1]), .Z(
        signal_3698) );
  XOR2_X1 cell_1920_U3 ( .A(signal_2096), .B(cell_1920_and_out[0]), .Z(
        signal_2188) );
  XOR2_X1 cell_1920_U2 ( .A(signal_3534), .B(signal_3465), .Z(
        cell_1920_and_in[1]) );
  XOR2_X1 cell_1920_U1 ( .A(signal_2096), .B(signal_2027), .Z(
        cell_1920_and_in[0]) );
  XOR2_X1 cell_1920_a_HPC2_and_U14 ( .A(Fresh[206]), .B(cell_1920_and_in[0]), 
        .Z(cell_1920_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1920_a_HPC2_and_U13 ( .A(Fresh[206]), .B(cell_1920_and_in[1]), 
        .Z(cell_1920_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1920_a_HPC2_and_U12 ( .A1(cell_1920_a_HPC2_and_a_reg[1]), .A2(
        cell_1920_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1920_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1920_a_HPC2_and_U11 ( .A1(cell_1920_a_HPC2_and_a_reg[0]), .A2(
        cell_1920_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1920_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1920_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1920_a_HPC2_and_n9), 
        .ZN(cell_1920_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1920_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1920_a_HPC2_and_n9), 
        .ZN(cell_1920_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1920_a_HPC2_and_U8 ( .A(Fresh[206]), .ZN(cell_1920_a_HPC2_and_n9) );
  AND2_X1 cell_1920_a_HPC2_and_U7 ( .A1(cell_1920_and_in[1]), .A2(n445), .ZN(
        cell_1920_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1920_a_HPC2_and_U6 ( .A1(cell_1920_and_in[0]), .A2(n431), .ZN(
        cell_1920_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1920_a_HPC2_and_U5 ( .A(cell_1920_a_HPC2_and_n8), .B(
        cell_1920_a_HPC2_and_z_1__1_), .ZN(cell_1920_and_out[1]) );
  XNOR2_X1 cell_1920_a_HPC2_and_U4 ( .A(
        cell_1920_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1920_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1920_a_HPC2_and_n8) );
  XNOR2_X1 cell_1920_a_HPC2_and_U3 ( .A(cell_1920_a_HPC2_and_n7), .B(
        cell_1920_a_HPC2_and_z_0__0_), .ZN(cell_1920_and_out[0]) );
  XNOR2_X1 cell_1920_a_HPC2_and_U2 ( .A(
        cell_1920_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1920_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1920_a_HPC2_and_n7) );
  DFF_X1 cell_1920_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1920_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1920_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1920_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1920_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1920_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1920_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1920_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1920_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1920_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1921_U4 ( .A(signal_3539), .B(cell_1921_and_out[1]), .Z(
        signal_3699) );
  XOR2_X1 cell_1921_U3 ( .A(signal_2101), .B(cell_1921_and_out[0]), .Z(
        signal_2189) );
  XOR2_X1 cell_1921_U2 ( .A(signal_3539), .B(signal_3477), .Z(
        cell_1921_and_in[1]) );
  XOR2_X1 cell_1921_U1 ( .A(signal_2101), .B(signal_2039), .Z(
        cell_1921_and_in[0]) );
  XOR2_X1 cell_1921_a_HPC2_and_U14 ( .A(Fresh[207]), .B(cell_1921_and_in[0]), 
        .Z(cell_1921_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1921_a_HPC2_and_U13 ( .A(Fresh[207]), .B(cell_1921_and_in[1]), 
        .Z(cell_1921_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1921_a_HPC2_and_U12 ( .A1(cell_1921_a_HPC2_and_a_reg[1]), .A2(
        cell_1921_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1921_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1921_a_HPC2_and_U11 ( .A1(cell_1921_a_HPC2_and_a_reg[0]), .A2(
        cell_1921_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1921_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1921_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1921_a_HPC2_and_n9), 
        .ZN(cell_1921_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1921_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1921_a_HPC2_and_n9), 
        .ZN(cell_1921_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1921_a_HPC2_and_U8 ( .A(Fresh[207]), .ZN(cell_1921_a_HPC2_and_n9) );
  AND2_X1 cell_1921_a_HPC2_and_U7 ( .A1(cell_1921_and_in[1]), .A2(n446), .ZN(
        cell_1921_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1921_a_HPC2_and_U6 ( .A1(cell_1921_and_in[0]), .A2(n432), .ZN(
        cell_1921_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1921_a_HPC2_and_U5 ( .A(cell_1921_a_HPC2_and_n8), .B(
        cell_1921_a_HPC2_and_z_1__1_), .ZN(cell_1921_and_out[1]) );
  XNOR2_X1 cell_1921_a_HPC2_and_U4 ( .A(
        cell_1921_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1921_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1921_a_HPC2_and_n8) );
  XNOR2_X1 cell_1921_a_HPC2_and_U3 ( .A(cell_1921_a_HPC2_and_n7), .B(
        cell_1921_a_HPC2_and_z_0__0_), .ZN(cell_1921_and_out[0]) );
  XNOR2_X1 cell_1921_a_HPC2_and_U2 ( .A(
        cell_1921_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1921_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1921_a_HPC2_and_n7) );
  DFF_X1 cell_1921_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1921_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1921_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1921_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1921_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1921_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1921_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1921_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1921_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1921_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1922_U4 ( .A(signal_3548), .B(cell_1922_and_out[1]), .Z(
        signal_3700) );
  XOR2_X1 cell_1922_U3 ( .A(signal_2110), .B(cell_1922_and_out[0]), .Z(
        signal_2190) );
  XOR2_X1 cell_1922_U2 ( .A(signal_3548), .B(signal_3566), .Z(
        cell_1922_and_in[1]) );
  XOR2_X1 cell_1922_U1 ( .A(signal_2110), .B(signal_2128), .Z(
        cell_1922_and_in[0]) );
  XOR2_X1 cell_1922_a_HPC2_and_U14 ( .A(Fresh[208]), .B(cell_1922_and_in[0]), 
        .Z(cell_1922_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1922_a_HPC2_and_U13 ( .A(Fresh[208]), .B(cell_1922_and_in[1]), 
        .Z(cell_1922_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1922_a_HPC2_and_U12 ( .A1(cell_1922_a_HPC2_and_a_reg[1]), .A2(
        cell_1922_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1922_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1922_a_HPC2_and_U11 ( .A1(cell_1922_a_HPC2_and_a_reg[0]), .A2(
        cell_1922_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1922_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1922_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1922_a_HPC2_and_n9), 
        .ZN(cell_1922_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1922_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1922_a_HPC2_and_n9), 
        .ZN(cell_1922_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1922_a_HPC2_and_U8 ( .A(Fresh[208]), .ZN(cell_1922_a_HPC2_and_n9) );
  AND2_X1 cell_1922_a_HPC2_and_U7 ( .A1(cell_1922_and_in[1]), .A2(n447), .ZN(
        cell_1922_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1922_a_HPC2_and_U6 ( .A1(cell_1922_and_in[0]), .A2(n433), .ZN(
        cell_1922_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1922_a_HPC2_and_U5 ( .A(cell_1922_a_HPC2_and_n8), .B(
        cell_1922_a_HPC2_and_z_1__1_), .ZN(cell_1922_and_out[1]) );
  XNOR2_X1 cell_1922_a_HPC2_and_U4 ( .A(
        cell_1922_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1922_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1922_a_HPC2_and_n8) );
  XNOR2_X1 cell_1922_a_HPC2_and_U3 ( .A(cell_1922_a_HPC2_and_n7), .B(
        cell_1922_a_HPC2_and_z_0__0_), .ZN(cell_1922_and_out[0]) );
  XNOR2_X1 cell_1922_a_HPC2_and_U2 ( .A(
        cell_1922_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1922_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1922_a_HPC2_and_n7) );
  DFF_X1 cell_1922_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1922_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1922_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1922_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1922_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1922_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1922_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1922_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1922_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1922_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1923_U4 ( .A(signal_3499), .B(cell_1923_and_out[1]), .Z(
        signal_3701) );
  XOR2_X1 cell_1923_U3 ( .A(signal_2061), .B(cell_1923_and_out[0]), .Z(
        signal_2191) );
  XOR2_X1 cell_1923_U2 ( .A(signal_3499), .B(signal_3514), .Z(
        cell_1923_and_in[1]) );
  XOR2_X1 cell_1923_U1 ( .A(signal_2061), .B(signal_2076), .Z(
        cell_1923_and_in[0]) );
  XOR2_X1 cell_1923_a_HPC2_and_U14 ( .A(Fresh[209]), .B(cell_1923_and_in[0]), 
        .Z(cell_1923_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1923_a_HPC2_and_U13 ( .A(Fresh[209]), .B(cell_1923_and_in[1]), 
        .Z(cell_1923_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1923_a_HPC2_and_U12 ( .A1(cell_1923_a_HPC2_and_a_reg[1]), .A2(
        cell_1923_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1923_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1923_a_HPC2_and_U11 ( .A1(cell_1923_a_HPC2_and_a_reg[0]), .A2(
        cell_1923_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1923_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1923_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1923_a_HPC2_and_n9), 
        .ZN(cell_1923_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1923_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1923_a_HPC2_and_n9), 
        .ZN(cell_1923_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1923_a_HPC2_and_U8 ( .A(Fresh[209]), .ZN(cell_1923_a_HPC2_and_n9) );
  AND2_X1 cell_1923_a_HPC2_and_U7 ( .A1(cell_1923_and_in[1]), .A2(n452), .ZN(
        cell_1923_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1923_a_HPC2_and_U6 ( .A1(cell_1923_and_in[0]), .A2(n438), .ZN(
        cell_1923_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1923_a_HPC2_and_U5 ( .A(cell_1923_a_HPC2_and_n8), .B(
        cell_1923_a_HPC2_and_z_1__1_), .ZN(cell_1923_and_out[1]) );
  XNOR2_X1 cell_1923_a_HPC2_and_U4 ( .A(
        cell_1923_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1923_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1923_a_HPC2_and_n8) );
  XNOR2_X1 cell_1923_a_HPC2_and_U3 ( .A(cell_1923_a_HPC2_and_n7), .B(
        cell_1923_a_HPC2_and_z_0__0_), .ZN(cell_1923_and_out[0]) );
  XNOR2_X1 cell_1923_a_HPC2_and_U2 ( .A(
        cell_1923_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1923_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1923_a_HPC2_and_n7) );
  DFF_X1 cell_1923_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1923_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1923_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1923_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1923_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1923_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1923_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1923_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1923_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1923_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1924_U4 ( .A(signal_3498), .B(cell_1924_and_out[1]), .Z(
        signal_3702) );
  XOR2_X1 cell_1924_U3 ( .A(signal_2060), .B(cell_1924_and_out[0]), .Z(
        signal_2192) );
  XOR2_X1 cell_1924_U2 ( .A(signal_3498), .B(signal_3491), .Z(
        cell_1924_and_in[1]) );
  XOR2_X1 cell_1924_U1 ( .A(signal_2060), .B(signal_2053), .Z(
        cell_1924_and_in[0]) );
  XOR2_X1 cell_1924_a_HPC2_and_U14 ( .A(Fresh[210]), .B(cell_1924_and_in[0]), 
        .Z(cell_1924_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1924_a_HPC2_and_U13 ( .A(Fresh[210]), .B(cell_1924_and_in[1]), 
        .Z(cell_1924_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1924_a_HPC2_and_U12 ( .A1(cell_1924_a_HPC2_and_a_reg[1]), .A2(
        cell_1924_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1924_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1924_a_HPC2_and_U11 ( .A1(cell_1924_a_HPC2_and_a_reg[0]), .A2(
        cell_1924_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1924_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1924_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1924_a_HPC2_and_n9), 
        .ZN(cell_1924_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1924_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1924_a_HPC2_and_n9), 
        .ZN(cell_1924_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1924_a_HPC2_and_U8 ( .A(Fresh[210]), .ZN(cell_1924_a_HPC2_and_n9) );
  AND2_X1 cell_1924_a_HPC2_and_U7 ( .A1(cell_1924_and_in[1]), .A2(n448), .ZN(
        cell_1924_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1924_a_HPC2_and_U6 ( .A1(cell_1924_and_in[0]), .A2(n434), .ZN(
        cell_1924_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1924_a_HPC2_and_U5 ( .A(cell_1924_a_HPC2_and_n8), .B(
        cell_1924_a_HPC2_and_z_1__1_), .ZN(cell_1924_and_out[1]) );
  XNOR2_X1 cell_1924_a_HPC2_and_U4 ( .A(
        cell_1924_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1924_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1924_a_HPC2_and_n8) );
  XNOR2_X1 cell_1924_a_HPC2_and_U3 ( .A(cell_1924_a_HPC2_and_n7), .B(
        cell_1924_a_HPC2_and_z_0__0_), .ZN(cell_1924_and_out[0]) );
  XNOR2_X1 cell_1924_a_HPC2_and_U2 ( .A(
        cell_1924_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1924_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1924_a_HPC2_and_n7) );
  DFF_X1 cell_1924_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1924_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1924_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1924_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1924_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1924_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1924_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1924_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1924_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1924_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1925_U4 ( .A(n383), .B(cell_1925_and_out[1]), .Z(signal_3703)
         );
  XOR2_X1 cell_1925_U3 ( .A(n382), .B(cell_1925_and_out[0]), .Z(signal_2193)
         );
  XOR2_X1 cell_1925_U2 ( .A(n383), .B(signal_3472), .Z(cell_1925_and_in[1]) );
  XOR2_X1 cell_1925_U1 ( .A(n382), .B(signal_2034), .Z(cell_1925_and_in[0]) );
  XOR2_X1 cell_1925_a_HPC2_and_U14 ( .A(Fresh[211]), .B(cell_1925_and_in[0]), 
        .Z(cell_1925_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1925_a_HPC2_and_U13 ( .A(Fresh[211]), .B(cell_1925_and_in[1]), 
        .Z(cell_1925_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1925_a_HPC2_and_U12 ( .A1(cell_1925_a_HPC2_and_a_reg[1]), .A2(
        cell_1925_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1925_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1925_a_HPC2_and_U11 ( .A1(cell_1925_a_HPC2_and_a_reg[0]), .A2(
        cell_1925_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1925_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1925_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1925_a_HPC2_and_n9), 
        .ZN(cell_1925_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1925_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1925_a_HPC2_and_n9), 
        .ZN(cell_1925_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1925_a_HPC2_and_U8 ( .A(Fresh[211]), .ZN(cell_1925_a_HPC2_and_n9) );
  AND2_X1 cell_1925_a_HPC2_and_U7 ( .A1(cell_1925_and_in[1]), .A2(n452), .ZN(
        cell_1925_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1925_a_HPC2_and_U6 ( .A1(cell_1925_and_in[0]), .A2(n438), .ZN(
        cell_1925_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1925_a_HPC2_and_U5 ( .A(cell_1925_a_HPC2_and_n8), .B(
        cell_1925_a_HPC2_and_z_1__1_), .ZN(cell_1925_and_out[1]) );
  XNOR2_X1 cell_1925_a_HPC2_and_U4 ( .A(
        cell_1925_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1925_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1925_a_HPC2_and_n8) );
  XNOR2_X1 cell_1925_a_HPC2_and_U3 ( .A(cell_1925_a_HPC2_and_n7), .B(
        cell_1925_a_HPC2_and_z_0__0_), .ZN(cell_1925_and_out[0]) );
  XNOR2_X1 cell_1925_a_HPC2_and_U2 ( .A(
        cell_1925_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1925_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1925_a_HPC2_and_n7) );
  DFF_X1 cell_1925_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1925_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1925_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1925_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1925_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1925_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1925_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1925_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1925_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1925_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1926_U4 ( .A(signal_3475), .B(cell_1926_and_out[1]), .Z(
        signal_3704) );
  XOR2_X1 cell_1926_U3 ( .A(signal_2037), .B(cell_1926_and_out[0]), .Z(
        signal_2194) );
  XOR2_X1 cell_1926_U2 ( .A(signal_3475), .B(signal_3544), .Z(
        cell_1926_and_in[1]) );
  XOR2_X1 cell_1926_U1 ( .A(signal_2037), .B(signal_2106), .Z(
        cell_1926_and_in[0]) );
  XOR2_X1 cell_1926_a_HPC2_and_U14 ( .A(Fresh[212]), .B(cell_1926_and_in[0]), 
        .Z(cell_1926_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1926_a_HPC2_and_U13 ( .A(Fresh[212]), .B(cell_1926_and_in[1]), 
        .Z(cell_1926_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1926_a_HPC2_and_U12 ( .A1(cell_1926_a_HPC2_and_a_reg[1]), .A2(
        cell_1926_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1926_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1926_a_HPC2_and_U11 ( .A1(cell_1926_a_HPC2_and_a_reg[0]), .A2(
        cell_1926_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1926_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1926_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1926_a_HPC2_and_n9), 
        .ZN(cell_1926_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1926_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1926_a_HPC2_and_n9), 
        .ZN(cell_1926_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1926_a_HPC2_and_U8 ( .A(Fresh[212]), .ZN(cell_1926_a_HPC2_and_n9) );
  AND2_X1 cell_1926_a_HPC2_and_U7 ( .A1(cell_1926_and_in[1]), .A2(n451), .ZN(
        cell_1926_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1926_a_HPC2_and_U6 ( .A1(cell_1926_and_in[0]), .A2(n437), .ZN(
        cell_1926_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1926_a_HPC2_and_U5 ( .A(cell_1926_a_HPC2_and_n8), .B(
        cell_1926_a_HPC2_and_z_1__1_), .ZN(cell_1926_and_out[1]) );
  XNOR2_X1 cell_1926_a_HPC2_and_U4 ( .A(
        cell_1926_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1926_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1926_a_HPC2_and_n8) );
  XNOR2_X1 cell_1926_a_HPC2_and_U3 ( .A(cell_1926_a_HPC2_and_n7), .B(
        cell_1926_a_HPC2_and_z_0__0_), .ZN(cell_1926_and_out[0]) );
  XNOR2_X1 cell_1926_a_HPC2_and_U2 ( .A(
        cell_1926_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1926_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1926_a_HPC2_and_n7) );
  DFF_X1 cell_1926_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1926_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1926_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1926_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1926_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1926_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1926_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1926_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1926_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1926_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1927_U4 ( .A(signal_3482), .B(cell_1927_and_out[1]), .Z(
        signal_3705) );
  XOR2_X1 cell_1927_U3 ( .A(signal_2044), .B(cell_1927_and_out[0]), .Z(
        signal_2195) );
  XOR2_X1 cell_1927_U2 ( .A(signal_3482), .B(signal_3507), .Z(
        cell_1927_and_in[1]) );
  XOR2_X1 cell_1927_U1 ( .A(signal_2044), .B(signal_2069), .Z(
        cell_1927_and_in[0]) );
  XOR2_X1 cell_1927_a_HPC2_and_U14 ( .A(Fresh[213]), .B(cell_1927_and_in[0]), 
        .Z(cell_1927_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1927_a_HPC2_and_U13 ( .A(Fresh[213]), .B(cell_1927_and_in[1]), 
        .Z(cell_1927_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1927_a_HPC2_and_U12 ( .A1(cell_1927_a_HPC2_and_a_reg[1]), .A2(
        cell_1927_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1927_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1927_a_HPC2_and_U11 ( .A1(cell_1927_a_HPC2_and_a_reg[0]), .A2(
        cell_1927_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1927_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1927_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1927_a_HPC2_and_n9), 
        .ZN(cell_1927_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1927_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1927_a_HPC2_and_n9), 
        .ZN(cell_1927_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1927_a_HPC2_and_U8 ( .A(Fresh[213]), .ZN(cell_1927_a_HPC2_and_n9) );
  AND2_X1 cell_1927_a_HPC2_and_U7 ( .A1(cell_1927_and_in[1]), .A2(n444), .ZN(
        cell_1927_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1927_a_HPC2_and_U6 ( .A1(cell_1927_and_in[0]), .A2(n430), .ZN(
        cell_1927_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1927_a_HPC2_and_U5 ( .A(cell_1927_a_HPC2_and_n8), .B(
        cell_1927_a_HPC2_and_z_1__1_), .ZN(cell_1927_and_out[1]) );
  XNOR2_X1 cell_1927_a_HPC2_and_U4 ( .A(
        cell_1927_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1927_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1927_a_HPC2_and_n8) );
  XNOR2_X1 cell_1927_a_HPC2_and_U3 ( .A(cell_1927_a_HPC2_and_n7), .B(
        cell_1927_a_HPC2_and_z_0__0_), .ZN(cell_1927_and_out[0]) );
  XNOR2_X1 cell_1927_a_HPC2_and_U2 ( .A(
        cell_1927_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1927_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1927_a_HPC2_and_n7) );
  DFF_X1 cell_1927_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1927_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1927_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1927_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1927_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1927_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1927_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1927_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1927_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1927_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1928_U4 ( .A(signal_3547), .B(cell_1928_and_out[1]), .Z(
        signal_3706) );
  XOR2_X1 cell_1928_U3 ( .A(signal_2109), .B(cell_1928_and_out[0]), .Z(
        signal_2196) );
  XOR2_X1 cell_1928_U2 ( .A(signal_3547), .B(signal_3413), .Z(
        cell_1928_and_in[1]) );
  XOR2_X1 cell_1928_U1 ( .A(signal_2109), .B(signal_1999), .Z(
        cell_1928_and_in[0]) );
  XOR2_X1 cell_1928_a_HPC2_and_U14 ( .A(Fresh[214]), .B(cell_1928_and_in[0]), 
        .Z(cell_1928_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1928_a_HPC2_and_U13 ( .A(Fresh[214]), .B(cell_1928_and_in[1]), 
        .Z(cell_1928_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1928_a_HPC2_and_U12 ( .A1(cell_1928_a_HPC2_and_a_reg[1]), .A2(
        cell_1928_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1928_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1928_a_HPC2_and_U11 ( .A1(cell_1928_a_HPC2_and_a_reg[0]), .A2(
        cell_1928_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1928_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1928_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1928_a_HPC2_and_n9), 
        .ZN(cell_1928_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1928_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1928_a_HPC2_and_n9), 
        .ZN(cell_1928_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1928_a_HPC2_and_U8 ( .A(Fresh[214]), .ZN(cell_1928_a_HPC2_and_n9) );
  AND2_X1 cell_1928_a_HPC2_and_U7 ( .A1(cell_1928_and_in[1]), .A2(n444), .ZN(
        cell_1928_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1928_a_HPC2_and_U6 ( .A1(cell_1928_and_in[0]), .A2(n430), .ZN(
        cell_1928_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1928_a_HPC2_and_U5 ( .A(cell_1928_a_HPC2_and_n8), .B(
        cell_1928_a_HPC2_and_z_1__1_), .ZN(cell_1928_and_out[1]) );
  XNOR2_X1 cell_1928_a_HPC2_and_U4 ( .A(
        cell_1928_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1928_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1928_a_HPC2_and_n8) );
  XNOR2_X1 cell_1928_a_HPC2_and_U3 ( .A(cell_1928_a_HPC2_and_n7), .B(
        cell_1928_a_HPC2_and_z_0__0_), .ZN(cell_1928_and_out[0]) );
  XNOR2_X1 cell_1928_a_HPC2_and_U2 ( .A(
        cell_1928_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1928_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1928_a_HPC2_and_n7) );
  DFF_X1 cell_1928_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1928_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1928_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1928_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1928_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1928_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1928_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1928_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1928_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1928_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1929_U4 ( .A(signal_3463), .B(cell_1929_and_out[1]), .Z(
        signal_3707) );
  XOR2_X1 cell_1929_U3 ( .A(signal_2025), .B(cell_1929_and_out[0]), .Z(
        signal_2197) );
  XOR2_X1 cell_1929_U2 ( .A(signal_3463), .B(signal_3580), .Z(
        cell_1929_and_in[1]) );
  XOR2_X1 cell_1929_U1 ( .A(signal_2025), .B(signal_2142), .Z(
        cell_1929_and_in[0]) );
  XOR2_X1 cell_1929_a_HPC2_and_U14 ( .A(Fresh[215]), .B(cell_1929_and_in[0]), 
        .Z(cell_1929_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1929_a_HPC2_and_U13 ( .A(Fresh[215]), .B(cell_1929_and_in[1]), 
        .Z(cell_1929_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1929_a_HPC2_and_U12 ( .A1(cell_1929_a_HPC2_and_a_reg[1]), .A2(
        cell_1929_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1929_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1929_a_HPC2_and_U11 ( .A1(cell_1929_a_HPC2_and_a_reg[0]), .A2(
        cell_1929_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1929_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1929_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1929_a_HPC2_and_n9), 
        .ZN(cell_1929_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1929_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1929_a_HPC2_and_n9), 
        .ZN(cell_1929_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1929_a_HPC2_and_U8 ( .A(Fresh[215]), .ZN(cell_1929_a_HPC2_and_n9) );
  AND2_X1 cell_1929_a_HPC2_and_U7 ( .A1(cell_1929_and_in[1]), .A2(n444), .ZN(
        cell_1929_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1929_a_HPC2_and_U6 ( .A1(cell_1929_and_in[0]), .A2(n430), .ZN(
        cell_1929_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1929_a_HPC2_and_U5 ( .A(cell_1929_a_HPC2_and_n8), .B(
        cell_1929_a_HPC2_and_z_1__1_), .ZN(cell_1929_and_out[1]) );
  XNOR2_X1 cell_1929_a_HPC2_and_U4 ( .A(
        cell_1929_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1929_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1929_a_HPC2_and_n8) );
  XNOR2_X1 cell_1929_a_HPC2_and_U3 ( .A(cell_1929_a_HPC2_and_n7), .B(
        cell_1929_a_HPC2_and_z_0__0_), .ZN(cell_1929_and_out[0]) );
  XNOR2_X1 cell_1929_a_HPC2_and_U2 ( .A(
        cell_1929_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1929_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1929_a_HPC2_and_n7) );
  DFF_X1 cell_1929_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1929_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1929_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1929_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1929_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1929_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1929_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1929_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1929_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1929_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1930_U4 ( .A(signal_3564), .B(cell_1930_and_out[1]), .Z(
        signal_3708) );
  XOR2_X1 cell_1930_U3 ( .A(signal_2126), .B(cell_1930_and_out[0]), .Z(
        signal_2198) );
  XOR2_X1 cell_1930_U2 ( .A(signal_3564), .B(signal_3502), .Z(
        cell_1930_and_in[1]) );
  XOR2_X1 cell_1930_U1 ( .A(signal_2126), .B(signal_2064), .Z(
        cell_1930_and_in[0]) );
  XOR2_X1 cell_1930_a_HPC2_and_U14 ( .A(Fresh[216]), .B(cell_1930_and_in[0]), 
        .Z(cell_1930_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1930_a_HPC2_and_U13 ( .A(Fresh[216]), .B(cell_1930_and_in[1]), 
        .Z(cell_1930_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1930_a_HPC2_and_U12 ( .A1(cell_1930_a_HPC2_and_a_reg[1]), .A2(
        cell_1930_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1930_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1930_a_HPC2_and_U11 ( .A1(cell_1930_a_HPC2_and_a_reg[0]), .A2(
        cell_1930_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1930_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1930_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1930_a_HPC2_and_n9), 
        .ZN(cell_1930_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1930_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1930_a_HPC2_and_n9), 
        .ZN(cell_1930_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1930_a_HPC2_and_U8 ( .A(Fresh[216]), .ZN(cell_1930_a_HPC2_and_n9) );
  AND2_X1 cell_1930_a_HPC2_and_U7 ( .A1(cell_1930_and_in[1]), .A2(n452), .ZN(
        cell_1930_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1930_a_HPC2_and_U6 ( .A1(cell_1930_and_in[0]), .A2(n438), .ZN(
        cell_1930_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1930_a_HPC2_and_U5 ( .A(cell_1930_a_HPC2_and_n8), .B(
        cell_1930_a_HPC2_and_z_1__1_), .ZN(cell_1930_and_out[1]) );
  XNOR2_X1 cell_1930_a_HPC2_and_U4 ( .A(
        cell_1930_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1930_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1930_a_HPC2_and_n8) );
  XNOR2_X1 cell_1930_a_HPC2_and_U3 ( .A(cell_1930_a_HPC2_and_n7), .B(
        cell_1930_a_HPC2_and_z_0__0_), .ZN(cell_1930_and_out[0]) );
  XNOR2_X1 cell_1930_a_HPC2_and_U2 ( .A(
        cell_1930_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1930_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1930_a_HPC2_and_n7) );
  DFF_X1 cell_1930_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1930_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1930_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1930_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1930_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1930_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1930_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1930_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1930_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1930_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1931_U4 ( .A(signal_3478), .B(cell_1931_and_out[1]), .Z(
        signal_3709) );
  XOR2_X1 cell_1931_U3 ( .A(signal_2040), .B(cell_1931_and_out[0]), .Z(
        signal_2199) );
  XOR2_X1 cell_1931_U2 ( .A(signal_3478), .B(signal_3543), .Z(
        cell_1931_and_in[1]) );
  XOR2_X1 cell_1931_U1 ( .A(signal_2040), .B(signal_2105), .Z(
        cell_1931_and_in[0]) );
  XOR2_X1 cell_1931_a_HPC2_and_U14 ( .A(Fresh[217]), .B(cell_1931_and_in[0]), 
        .Z(cell_1931_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1931_a_HPC2_and_U13 ( .A(Fresh[217]), .B(cell_1931_and_in[1]), 
        .Z(cell_1931_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1931_a_HPC2_and_U12 ( .A1(cell_1931_a_HPC2_and_a_reg[1]), .A2(
        cell_1931_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1931_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1931_a_HPC2_and_U11 ( .A1(cell_1931_a_HPC2_and_a_reg[0]), .A2(
        cell_1931_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1931_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1931_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1931_a_HPC2_and_n9), 
        .ZN(cell_1931_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1931_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1931_a_HPC2_and_n9), 
        .ZN(cell_1931_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1931_a_HPC2_and_U8 ( .A(Fresh[217]), .ZN(cell_1931_a_HPC2_and_n9) );
  AND2_X1 cell_1931_a_HPC2_and_U7 ( .A1(cell_1931_and_in[1]), .A2(n452), .ZN(
        cell_1931_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1931_a_HPC2_and_U6 ( .A1(cell_1931_and_in[0]), .A2(n438), .ZN(
        cell_1931_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1931_a_HPC2_and_U5 ( .A(cell_1931_a_HPC2_and_n8), .B(
        cell_1931_a_HPC2_and_z_1__1_), .ZN(cell_1931_and_out[1]) );
  XNOR2_X1 cell_1931_a_HPC2_and_U4 ( .A(
        cell_1931_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1931_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1931_a_HPC2_and_n8) );
  XNOR2_X1 cell_1931_a_HPC2_and_U3 ( .A(cell_1931_a_HPC2_and_n7), .B(
        cell_1931_a_HPC2_and_z_0__0_), .ZN(cell_1931_and_out[0]) );
  XNOR2_X1 cell_1931_a_HPC2_and_U2 ( .A(
        cell_1931_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1931_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1931_a_HPC2_and_n7) );
  DFF_X1 cell_1931_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1931_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1931_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1931_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1931_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1931_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1931_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1931_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1931_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1931_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1932_U4 ( .A(signal_3565), .B(cell_1932_and_out[1]), .Z(
        signal_3710) );
  XOR2_X1 cell_1932_U3 ( .A(signal_2127), .B(cell_1932_and_out[0]), .Z(
        signal_2200) );
  XOR2_X1 cell_1932_U2 ( .A(signal_3565), .B(signal_3402), .Z(
        cell_1932_and_in[1]) );
  XOR2_X1 cell_1932_U1 ( .A(signal_2127), .B(signal_1988), .Z(
        cell_1932_and_in[0]) );
  XOR2_X1 cell_1932_a_HPC2_and_U14 ( .A(Fresh[218]), .B(cell_1932_and_in[0]), 
        .Z(cell_1932_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1932_a_HPC2_and_U13 ( .A(Fresh[218]), .B(cell_1932_and_in[1]), 
        .Z(cell_1932_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1932_a_HPC2_and_U12 ( .A1(cell_1932_a_HPC2_and_a_reg[1]), .A2(
        cell_1932_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1932_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1932_a_HPC2_and_U11 ( .A1(cell_1932_a_HPC2_and_a_reg[0]), .A2(
        cell_1932_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1932_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1932_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1932_a_HPC2_and_n9), 
        .ZN(cell_1932_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1932_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1932_a_HPC2_and_n9), 
        .ZN(cell_1932_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1932_a_HPC2_and_U8 ( .A(Fresh[218]), .ZN(cell_1932_a_HPC2_and_n9) );
  AND2_X1 cell_1932_a_HPC2_and_U7 ( .A1(cell_1932_and_in[1]), .A2(n452), .ZN(
        cell_1932_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1932_a_HPC2_and_U6 ( .A1(cell_1932_and_in[0]), .A2(n438), .ZN(
        cell_1932_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1932_a_HPC2_and_U5 ( .A(cell_1932_a_HPC2_and_n8), .B(
        cell_1932_a_HPC2_and_z_1__1_), .ZN(cell_1932_and_out[1]) );
  XNOR2_X1 cell_1932_a_HPC2_and_U4 ( .A(
        cell_1932_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1932_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1932_a_HPC2_and_n8) );
  XNOR2_X1 cell_1932_a_HPC2_and_U3 ( .A(cell_1932_a_HPC2_and_n7), .B(
        cell_1932_a_HPC2_and_z_0__0_), .ZN(cell_1932_and_out[0]) );
  XNOR2_X1 cell_1932_a_HPC2_and_U2 ( .A(
        cell_1932_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1932_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1932_a_HPC2_and_n7) );
  DFF_X1 cell_1932_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1932_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1932_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1932_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1932_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1932_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1932_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1932_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1932_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1932_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1933_U4 ( .A(signal_3405), .B(cell_1933_and_out[1]), .Z(
        signal_3711) );
  XOR2_X1 cell_1933_U3 ( .A(signal_1991), .B(cell_1933_and_out[0]), .Z(
        signal_2201) );
  XOR2_X1 cell_1933_U2 ( .A(signal_3405), .B(signal_3579), .Z(
        cell_1933_and_in[1]) );
  XOR2_X1 cell_1933_U1 ( .A(signal_1991), .B(signal_2141), .Z(
        cell_1933_and_in[0]) );
  XOR2_X1 cell_1933_a_HPC2_and_U14 ( .A(Fresh[219]), .B(cell_1933_and_in[0]), 
        .Z(cell_1933_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1933_a_HPC2_and_U13 ( .A(Fresh[219]), .B(cell_1933_and_in[1]), 
        .Z(cell_1933_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1933_a_HPC2_and_U12 ( .A1(cell_1933_a_HPC2_and_a_reg[1]), .A2(
        cell_1933_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1933_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1933_a_HPC2_and_U11 ( .A1(cell_1933_a_HPC2_and_a_reg[0]), .A2(
        cell_1933_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1933_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1933_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1933_a_HPC2_and_n9), 
        .ZN(cell_1933_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1933_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1933_a_HPC2_and_n9), 
        .ZN(cell_1933_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1933_a_HPC2_and_U8 ( .A(Fresh[219]), .ZN(cell_1933_a_HPC2_and_n9) );
  AND2_X1 cell_1933_a_HPC2_and_U7 ( .A1(cell_1933_and_in[1]), .A2(n453), .ZN(
        cell_1933_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1933_a_HPC2_and_U6 ( .A1(cell_1933_and_in[0]), .A2(n439), .ZN(
        cell_1933_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1933_a_HPC2_and_U5 ( .A(cell_1933_a_HPC2_and_n8), .B(
        cell_1933_a_HPC2_and_z_1__1_), .ZN(cell_1933_and_out[1]) );
  XNOR2_X1 cell_1933_a_HPC2_and_U4 ( .A(
        cell_1933_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1933_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1933_a_HPC2_and_n8) );
  XNOR2_X1 cell_1933_a_HPC2_and_U3 ( .A(cell_1933_a_HPC2_and_n7), .B(
        cell_1933_a_HPC2_and_z_0__0_), .ZN(cell_1933_and_out[0]) );
  XNOR2_X1 cell_1933_a_HPC2_and_U2 ( .A(
        cell_1933_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1933_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1933_a_HPC2_and_n7) );
  DFF_X1 cell_1933_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1933_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1933_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1933_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1933_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1933_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1933_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1933_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1933_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1933_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1934_U4 ( .A(signal_3506), .B(cell_1934_and_out[1]), .Z(
        signal_3712) );
  XOR2_X1 cell_1934_U3 ( .A(signal_2068), .B(cell_1934_and_out[0]), .Z(
        signal_2202) );
  XOR2_X1 cell_1934_U2 ( .A(signal_3506), .B(signal_3541), .Z(
        cell_1934_and_in[1]) );
  XOR2_X1 cell_1934_U1 ( .A(signal_2068), .B(signal_2103), .Z(
        cell_1934_and_in[0]) );
  XOR2_X1 cell_1934_a_HPC2_and_U14 ( .A(Fresh[220]), .B(cell_1934_and_in[0]), 
        .Z(cell_1934_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1934_a_HPC2_and_U13 ( .A(Fresh[220]), .B(cell_1934_and_in[1]), 
        .Z(cell_1934_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1934_a_HPC2_and_U12 ( .A1(cell_1934_a_HPC2_and_a_reg[1]), .A2(
        cell_1934_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1934_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1934_a_HPC2_and_U11 ( .A1(cell_1934_a_HPC2_and_a_reg[0]), .A2(
        cell_1934_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1934_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1934_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1934_a_HPC2_and_n9), 
        .ZN(cell_1934_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1934_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1934_a_HPC2_and_n9), 
        .ZN(cell_1934_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1934_a_HPC2_and_U8 ( .A(Fresh[220]), .ZN(cell_1934_a_HPC2_and_n9) );
  AND2_X1 cell_1934_a_HPC2_and_U7 ( .A1(cell_1934_and_in[1]), .A2(n444), .ZN(
        cell_1934_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1934_a_HPC2_and_U6 ( .A1(cell_1934_and_in[0]), .A2(n430), .ZN(
        cell_1934_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1934_a_HPC2_and_U5 ( .A(cell_1934_a_HPC2_and_n8), .B(
        cell_1934_a_HPC2_and_z_1__1_), .ZN(cell_1934_and_out[1]) );
  XNOR2_X1 cell_1934_a_HPC2_and_U4 ( .A(
        cell_1934_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1934_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1934_a_HPC2_and_n8) );
  XNOR2_X1 cell_1934_a_HPC2_and_U3 ( .A(cell_1934_a_HPC2_and_n7), .B(
        cell_1934_a_HPC2_and_z_0__0_), .ZN(cell_1934_and_out[0]) );
  XNOR2_X1 cell_1934_a_HPC2_and_U2 ( .A(
        cell_1934_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1934_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1934_a_HPC2_and_n7) );
  DFF_X1 cell_1934_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1934_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1934_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1934_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1934_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1934_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1934_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1934_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1934_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1934_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1935_U4 ( .A(signal_3486), .B(cell_1935_and_out[1]), .Z(
        signal_3713) );
  XOR2_X1 cell_1935_U3 ( .A(signal_2048), .B(cell_1935_and_out[0]), .Z(
        signal_2203) );
  XOR2_X1 cell_1935_U2 ( .A(signal_3486), .B(signal_3506), .Z(
        cell_1935_and_in[1]) );
  XOR2_X1 cell_1935_U1 ( .A(signal_2048), .B(signal_2068), .Z(
        cell_1935_and_in[0]) );
  XOR2_X1 cell_1935_a_HPC2_and_U14 ( .A(Fresh[221]), .B(cell_1935_and_in[0]), 
        .Z(cell_1935_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1935_a_HPC2_and_U13 ( .A(Fresh[221]), .B(cell_1935_and_in[1]), 
        .Z(cell_1935_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1935_a_HPC2_and_U12 ( .A1(cell_1935_a_HPC2_and_a_reg[1]), .A2(
        cell_1935_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1935_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1935_a_HPC2_and_U11 ( .A1(cell_1935_a_HPC2_and_a_reg[0]), .A2(
        cell_1935_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1935_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1935_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1935_a_HPC2_and_n9), 
        .ZN(cell_1935_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1935_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1935_a_HPC2_and_n9), 
        .ZN(cell_1935_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1935_a_HPC2_and_U8 ( .A(Fresh[221]), .ZN(cell_1935_a_HPC2_and_n9) );
  AND2_X1 cell_1935_a_HPC2_and_U7 ( .A1(cell_1935_and_in[1]), .A2(n444), .ZN(
        cell_1935_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1935_a_HPC2_and_U6 ( .A1(cell_1935_and_in[0]), .A2(n430), .ZN(
        cell_1935_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1935_a_HPC2_and_U5 ( .A(cell_1935_a_HPC2_and_n8), .B(
        cell_1935_a_HPC2_and_z_1__1_), .ZN(cell_1935_and_out[1]) );
  XNOR2_X1 cell_1935_a_HPC2_and_U4 ( .A(
        cell_1935_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1935_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1935_a_HPC2_and_n8) );
  XNOR2_X1 cell_1935_a_HPC2_and_U3 ( .A(cell_1935_a_HPC2_and_n7), .B(
        cell_1935_a_HPC2_and_z_0__0_), .ZN(cell_1935_and_out[0]) );
  XNOR2_X1 cell_1935_a_HPC2_and_U2 ( .A(
        cell_1935_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1935_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1935_a_HPC2_and_n7) );
  DFF_X1 cell_1935_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1935_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1935_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1935_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1935_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1935_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1935_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1935_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1935_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1935_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1936_U4 ( .A(signal_3590), .B(cell_1936_and_out[1]), .Z(
        signal_3714) );
  XOR2_X1 cell_1936_U3 ( .A(signal_2152), .B(cell_1936_and_out[0]), .Z(
        signal_2204) );
  XOR2_X1 cell_1936_U2 ( .A(signal_3590), .B(signal_3464), .Z(
        cell_1936_and_in[1]) );
  XOR2_X1 cell_1936_U1 ( .A(signal_2152), .B(signal_2026), .Z(
        cell_1936_and_in[0]) );
  XOR2_X1 cell_1936_a_HPC2_and_U14 ( .A(Fresh[222]), .B(cell_1936_and_in[0]), 
        .Z(cell_1936_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1936_a_HPC2_and_U13 ( .A(Fresh[222]), .B(cell_1936_and_in[1]), 
        .Z(cell_1936_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1936_a_HPC2_and_U12 ( .A1(cell_1936_a_HPC2_and_a_reg[1]), .A2(
        cell_1936_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1936_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1936_a_HPC2_and_U11 ( .A1(cell_1936_a_HPC2_and_a_reg[0]), .A2(
        cell_1936_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1936_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1936_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1936_a_HPC2_and_n9), 
        .ZN(cell_1936_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1936_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1936_a_HPC2_and_n9), 
        .ZN(cell_1936_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1936_a_HPC2_and_U8 ( .A(Fresh[222]), .ZN(cell_1936_a_HPC2_and_n9) );
  AND2_X1 cell_1936_a_HPC2_and_U7 ( .A1(cell_1936_and_in[1]), .A2(n444), .ZN(
        cell_1936_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1936_a_HPC2_and_U6 ( .A1(cell_1936_and_in[0]), .A2(n430), .ZN(
        cell_1936_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1936_a_HPC2_and_U5 ( .A(cell_1936_a_HPC2_and_n8), .B(
        cell_1936_a_HPC2_and_z_1__1_), .ZN(cell_1936_and_out[1]) );
  XNOR2_X1 cell_1936_a_HPC2_and_U4 ( .A(
        cell_1936_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1936_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1936_a_HPC2_and_n8) );
  XNOR2_X1 cell_1936_a_HPC2_and_U3 ( .A(cell_1936_a_HPC2_and_n7), .B(
        cell_1936_a_HPC2_and_z_0__0_), .ZN(cell_1936_and_out[0]) );
  XNOR2_X1 cell_1936_a_HPC2_and_U2 ( .A(
        cell_1936_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1936_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1936_a_HPC2_and_n7) );
  DFF_X1 cell_1936_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1936_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1936_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1936_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1936_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1936_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1936_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1936_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1936_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1936_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1937_U4 ( .A(signal_3513), .B(cell_1937_and_out[1]), .Z(
        signal_3715) );
  XOR2_X1 cell_1937_U3 ( .A(signal_2075), .B(cell_1937_and_out[0]), .Z(
        signal_2205) );
  XOR2_X1 cell_1937_U2 ( .A(signal_3513), .B(signal_3568), .Z(
        cell_1937_and_in[1]) );
  XOR2_X1 cell_1937_U1 ( .A(signal_2075), .B(signal_2130), .Z(
        cell_1937_and_in[0]) );
  XOR2_X1 cell_1937_a_HPC2_and_U14 ( .A(Fresh[223]), .B(cell_1937_and_in[0]), 
        .Z(cell_1937_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1937_a_HPC2_and_U13 ( .A(Fresh[223]), .B(cell_1937_and_in[1]), 
        .Z(cell_1937_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1937_a_HPC2_and_U12 ( .A1(cell_1937_a_HPC2_and_a_reg[1]), .A2(
        cell_1937_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1937_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1937_a_HPC2_and_U11 ( .A1(cell_1937_a_HPC2_and_a_reg[0]), .A2(
        cell_1937_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1937_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1937_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1937_a_HPC2_and_n9), 
        .ZN(cell_1937_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1937_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1937_a_HPC2_and_n9), 
        .ZN(cell_1937_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1937_a_HPC2_and_U8 ( .A(Fresh[223]), .ZN(cell_1937_a_HPC2_and_n9) );
  AND2_X1 cell_1937_a_HPC2_and_U7 ( .A1(cell_1937_and_in[1]), .A2(n453), .ZN(
        cell_1937_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1937_a_HPC2_and_U6 ( .A1(cell_1937_and_in[0]), .A2(n439), .ZN(
        cell_1937_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1937_a_HPC2_and_U5 ( .A(cell_1937_a_HPC2_and_n8), .B(
        cell_1937_a_HPC2_and_z_1__1_), .ZN(cell_1937_and_out[1]) );
  XNOR2_X1 cell_1937_a_HPC2_and_U4 ( .A(
        cell_1937_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1937_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1937_a_HPC2_and_n8) );
  XNOR2_X1 cell_1937_a_HPC2_and_U3 ( .A(cell_1937_a_HPC2_and_n7), .B(
        cell_1937_a_HPC2_and_z_0__0_), .ZN(cell_1937_and_out[0]) );
  XNOR2_X1 cell_1937_a_HPC2_and_U2 ( .A(
        cell_1937_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1937_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1937_a_HPC2_and_n7) );
  DFF_X1 cell_1937_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1937_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1937_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1937_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1937_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1937_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1937_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1937_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1937_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1937_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1938_U4 ( .A(signal_3466), .B(cell_1938_and_out[1]), .Z(
        signal_3716) );
  XOR2_X1 cell_1938_U3 ( .A(signal_2028), .B(cell_1938_and_out[0]), .Z(
        signal_2206) );
  XOR2_X1 cell_1938_U2 ( .A(signal_3466), .B(signal_3577), .Z(
        cell_1938_and_in[1]) );
  XOR2_X1 cell_1938_U1 ( .A(signal_2028), .B(signal_2139), .Z(
        cell_1938_and_in[0]) );
  XOR2_X1 cell_1938_a_HPC2_and_U14 ( .A(Fresh[224]), .B(cell_1938_and_in[0]), 
        .Z(cell_1938_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1938_a_HPC2_and_U13 ( .A(Fresh[224]), .B(cell_1938_and_in[1]), 
        .Z(cell_1938_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1938_a_HPC2_and_U12 ( .A1(cell_1938_a_HPC2_and_a_reg[1]), .A2(
        cell_1938_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1938_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1938_a_HPC2_and_U11 ( .A1(cell_1938_a_HPC2_and_a_reg[0]), .A2(
        cell_1938_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1938_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1938_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1938_a_HPC2_and_n9), 
        .ZN(cell_1938_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1938_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1938_a_HPC2_and_n9), 
        .ZN(cell_1938_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1938_a_HPC2_and_U8 ( .A(Fresh[224]), .ZN(cell_1938_a_HPC2_and_n9) );
  AND2_X1 cell_1938_a_HPC2_and_U7 ( .A1(cell_1938_and_in[1]), .A2(n453), .ZN(
        cell_1938_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1938_a_HPC2_and_U6 ( .A1(cell_1938_and_in[0]), .A2(n439), .ZN(
        cell_1938_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1938_a_HPC2_and_U5 ( .A(cell_1938_a_HPC2_and_n8), .B(
        cell_1938_a_HPC2_and_z_1__1_), .ZN(cell_1938_and_out[1]) );
  XNOR2_X1 cell_1938_a_HPC2_and_U4 ( .A(
        cell_1938_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1938_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1938_a_HPC2_and_n8) );
  XNOR2_X1 cell_1938_a_HPC2_and_U3 ( .A(cell_1938_a_HPC2_and_n7), .B(
        cell_1938_a_HPC2_and_z_0__0_), .ZN(cell_1938_and_out[0]) );
  XNOR2_X1 cell_1938_a_HPC2_and_U2 ( .A(
        cell_1938_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1938_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1938_a_HPC2_and_n7) );
  DFF_X1 cell_1938_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1938_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1938_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1938_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1938_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1938_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1938_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1938_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1938_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1938_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1939_U4 ( .A(signal_3523), .B(cell_1939_and_out[1]), .Z(
        signal_3717) );
  XOR2_X1 cell_1939_U3 ( .A(signal_2085), .B(cell_1939_and_out[0]), .Z(
        signal_2207) );
  XOR2_X1 cell_1939_U2 ( .A(signal_3523), .B(signal_3585), .Z(
        cell_1939_and_in[1]) );
  XOR2_X1 cell_1939_U1 ( .A(signal_2085), .B(signal_2147), .Z(
        cell_1939_and_in[0]) );
  XOR2_X1 cell_1939_a_HPC2_and_U14 ( .A(Fresh[225]), .B(cell_1939_and_in[0]), 
        .Z(cell_1939_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1939_a_HPC2_and_U13 ( .A(Fresh[225]), .B(cell_1939_and_in[1]), 
        .Z(cell_1939_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1939_a_HPC2_and_U12 ( .A1(cell_1939_a_HPC2_and_a_reg[1]), .A2(
        cell_1939_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1939_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1939_a_HPC2_and_U11 ( .A1(cell_1939_a_HPC2_and_a_reg[0]), .A2(
        cell_1939_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1939_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1939_a_HPC2_and_U10 ( .A1(n444), .A2(cell_1939_a_HPC2_and_n9), 
        .ZN(cell_1939_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1939_a_HPC2_and_U9 ( .A1(n430), .A2(cell_1939_a_HPC2_and_n9), 
        .ZN(cell_1939_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1939_a_HPC2_and_U8 ( .A(Fresh[225]), .ZN(cell_1939_a_HPC2_and_n9) );
  AND2_X1 cell_1939_a_HPC2_and_U7 ( .A1(cell_1939_and_in[1]), .A2(n444), .ZN(
        cell_1939_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1939_a_HPC2_and_U6 ( .A1(cell_1939_and_in[0]), .A2(n430), .ZN(
        cell_1939_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1939_a_HPC2_and_U5 ( .A(cell_1939_a_HPC2_and_n8), .B(
        cell_1939_a_HPC2_and_z_1__1_), .ZN(cell_1939_and_out[1]) );
  XNOR2_X1 cell_1939_a_HPC2_and_U4 ( .A(
        cell_1939_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1939_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1939_a_HPC2_and_n8) );
  XNOR2_X1 cell_1939_a_HPC2_and_U3 ( .A(cell_1939_a_HPC2_and_n7), .B(
        cell_1939_a_HPC2_and_z_0__0_), .ZN(cell_1939_and_out[0]) );
  XNOR2_X1 cell_1939_a_HPC2_and_U2 ( .A(
        cell_1939_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1939_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1939_a_HPC2_and_n7) );
  DFF_X1 cell_1939_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1939_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1939_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_1939_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1939_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1939_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_1939_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1939_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1939_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1939_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1940_U4 ( .A(signal_3534), .B(cell_1940_and_out[1]), .Z(
        signal_3718) );
  XOR2_X1 cell_1940_U3 ( .A(signal_2096), .B(cell_1940_and_out[0]), .Z(
        signal_2208) );
  XOR2_X1 cell_1940_U2 ( .A(signal_3534), .B(signal_3528), .Z(
        cell_1940_and_in[1]) );
  XOR2_X1 cell_1940_U1 ( .A(signal_2096), .B(signal_2090), .Z(
        cell_1940_and_in[0]) );
  XOR2_X1 cell_1940_a_HPC2_and_U14 ( .A(Fresh[226]), .B(cell_1940_and_in[0]), 
        .Z(cell_1940_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1940_a_HPC2_and_U13 ( .A(Fresh[226]), .B(cell_1940_and_in[1]), 
        .Z(cell_1940_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1940_a_HPC2_and_U12 ( .A1(cell_1940_a_HPC2_and_a_reg[1]), .A2(
        cell_1940_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1940_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1940_a_HPC2_and_U11 ( .A1(cell_1940_a_HPC2_and_a_reg[0]), .A2(
        cell_1940_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1940_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1940_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1940_a_HPC2_and_n9), 
        .ZN(cell_1940_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1940_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1940_a_HPC2_and_n9), 
        .ZN(cell_1940_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1940_a_HPC2_and_U8 ( .A(Fresh[226]), .ZN(cell_1940_a_HPC2_and_n9) );
  AND2_X1 cell_1940_a_HPC2_and_U7 ( .A1(cell_1940_and_in[1]), .A2(n445), .ZN(
        cell_1940_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1940_a_HPC2_and_U6 ( .A1(cell_1940_and_in[0]), .A2(n431), .ZN(
        cell_1940_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1940_a_HPC2_and_U5 ( .A(cell_1940_a_HPC2_and_n8), .B(
        cell_1940_a_HPC2_and_z_1__1_), .ZN(cell_1940_and_out[1]) );
  XNOR2_X1 cell_1940_a_HPC2_and_U4 ( .A(
        cell_1940_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1940_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1940_a_HPC2_and_n8) );
  XNOR2_X1 cell_1940_a_HPC2_and_U3 ( .A(cell_1940_a_HPC2_and_n7), .B(
        cell_1940_a_HPC2_and_z_0__0_), .ZN(cell_1940_and_out[0]) );
  XNOR2_X1 cell_1940_a_HPC2_and_U2 ( .A(
        cell_1940_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1940_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1940_a_HPC2_and_n7) );
  DFF_X1 cell_1940_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1940_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1940_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1940_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1940_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1940_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1940_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1940_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1940_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1940_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1941_U4 ( .A(signal_3545), .B(cell_1941_and_out[1]), .Z(
        signal_3719) );
  XOR2_X1 cell_1941_U3 ( .A(signal_2107), .B(cell_1941_and_out[0]), .Z(
        signal_2209) );
  XOR2_X1 cell_1941_U2 ( .A(signal_3545), .B(n379), .Z(cell_1941_and_in[1]) );
  XOR2_X1 cell_1941_U1 ( .A(signal_2107), .B(n377), .Z(cell_1941_and_in[0]) );
  XOR2_X1 cell_1941_a_HPC2_and_U14 ( .A(Fresh[227]), .B(cell_1941_and_in[0]), 
        .Z(cell_1941_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1941_a_HPC2_and_U13 ( .A(Fresh[227]), .B(cell_1941_and_in[1]), 
        .Z(cell_1941_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1941_a_HPC2_and_U12 ( .A1(cell_1941_a_HPC2_and_a_reg[1]), .A2(
        cell_1941_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1941_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1941_a_HPC2_and_U11 ( .A1(cell_1941_a_HPC2_and_a_reg[0]), .A2(
        cell_1941_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1941_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1941_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1941_a_HPC2_and_n9), 
        .ZN(cell_1941_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1941_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1941_a_HPC2_and_n9), 
        .ZN(cell_1941_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1941_a_HPC2_and_U8 ( .A(Fresh[227]), .ZN(cell_1941_a_HPC2_and_n9) );
  AND2_X1 cell_1941_a_HPC2_and_U7 ( .A1(cell_1941_and_in[1]), .A2(n445), .ZN(
        cell_1941_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1941_a_HPC2_and_U6 ( .A1(cell_1941_and_in[0]), .A2(n431), .ZN(
        cell_1941_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1941_a_HPC2_and_U5 ( .A(cell_1941_a_HPC2_and_n8), .B(
        cell_1941_a_HPC2_and_z_1__1_), .ZN(cell_1941_and_out[1]) );
  XNOR2_X1 cell_1941_a_HPC2_and_U4 ( .A(
        cell_1941_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1941_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1941_a_HPC2_and_n8) );
  XNOR2_X1 cell_1941_a_HPC2_and_U3 ( .A(cell_1941_a_HPC2_and_n7), .B(
        cell_1941_a_HPC2_and_z_0__0_), .ZN(cell_1941_and_out[0]) );
  XNOR2_X1 cell_1941_a_HPC2_and_U2 ( .A(
        cell_1941_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1941_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1941_a_HPC2_and_n7) );
  DFF_X1 cell_1941_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1941_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1941_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1941_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1941_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1941_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1941_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1941_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1941_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1941_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1942_U4 ( .A(signal_3500), .B(cell_1942_and_out[1]), .Z(
        signal_3720) );
  XOR2_X1 cell_1942_U3 ( .A(signal_2062), .B(cell_1942_and_out[0]), .Z(
        signal_2210) );
  XOR2_X1 cell_1942_U2 ( .A(signal_3500), .B(signal_3565), .Z(
        cell_1942_and_in[1]) );
  XOR2_X1 cell_1942_U1 ( .A(signal_2062), .B(signal_2127), .Z(
        cell_1942_and_in[0]) );
  XOR2_X1 cell_1942_a_HPC2_and_U14 ( .A(Fresh[228]), .B(cell_1942_and_in[0]), 
        .Z(cell_1942_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1942_a_HPC2_and_U13 ( .A(Fresh[228]), .B(cell_1942_and_in[1]), 
        .Z(cell_1942_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1942_a_HPC2_and_U12 ( .A1(cell_1942_a_HPC2_and_a_reg[1]), .A2(
        cell_1942_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1942_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1942_a_HPC2_and_U11 ( .A1(cell_1942_a_HPC2_and_a_reg[0]), .A2(
        cell_1942_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1942_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1942_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1942_a_HPC2_and_n9), 
        .ZN(cell_1942_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1942_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1942_a_HPC2_and_n9), 
        .ZN(cell_1942_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1942_a_HPC2_and_U8 ( .A(Fresh[228]), .ZN(cell_1942_a_HPC2_and_n9) );
  AND2_X1 cell_1942_a_HPC2_and_U7 ( .A1(cell_1942_and_in[1]), .A2(n445), .ZN(
        cell_1942_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1942_a_HPC2_and_U6 ( .A1(cell_1942_and_in[0]), .A2(n431), .ZN(
        cell_1942_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1942_a_HPC2_and_U5 ( .A(cell_1942_a_HPC2_and_n8), .B(
        cell_1942_a_HPC2_and_z_1__1_), .ZN(cell_1942_and_out[1]) );
  XNOR2_X1 cell_1942_a_HPC2_and_U4 ( .A(
        cell_1942_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1942_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1942_a_HPC2_and_n8) );
  XNOR2_X1 cell_1942_a_HPC2_and_U3 ( .A(cell_1942_a_HPC2_and_n7), .B(
        cell_1942_a_HPC2_and_z_0__0_), .ZN(cell_1942_and_out[0]) );
  XNOR2_X1 cell_1942_a_HPC2_and_U2 ( .A(
        cell_1942_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1942_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1942_a_HPC2_and_n7) );
  DFF_X1 cell_1942_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1942_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1942_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1942_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1942_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1942_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1942_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1942_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1942_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1942_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1943_U4 ( .A(signal_3489), .B(cell_1943_and_out[1]), .Z(
        signal_3721) );
  XOR2_X1 cell_1943_U3 ( .A(signal_2051), .B(cell_1943_and_out[0]), .Z(
        signal_2211) );
  XOR2_X1 cell_1943_U2 ( .A(signal_3489), .B(signal_3512), .Z(
        cell_1943_and_in[1]) );
  XOR2_X1 cell_1943_U1 ( .A(signal_2051), .B(signal_2074), .Z(
        cell_1943_and_in[0]) );
  XOR2_X1 cell_1943_a_HPC2_and_U14 ( .A(Fresh[229]), .B(cell_1943_and_in[0]), 
        .Z(cell_1943_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1943_a_HPC2_and_U13 ( .A(Fresh[229]), .B(cell_1943_and_in[1]), 
        .Z(cell_1943_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1943_a_HPC2_and_U12 ( .A1(cell_1943_a_HPC2_and_a_reg[1]), .A2(
        cell_1943_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1943_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1943_a_HPC2_and_U11 ( .A1(cell_1943_a_HPC2_and_a_reg[0]), .A2(
        cell_1943_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1943_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1943_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1943_a_HPC2_and_n9), 
        .ZN(cell_1943_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1943_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1943_a_HPC2_and_n9), 
        .ZN(cell_1943_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1943_a_HPC2_and_U8 ( .A(Fresh[229]), .ZN(cell_1943_a_HPC2_and_n9) );
  AND2_X1 cell_1943_a_HPC2_and_U7 ( .A1(cell_1943_and_in[1]), .A2(n445), .ZN(
        cell_1943_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1943_a_HPC2_and_U6 ( .A1(cell_1943_and_in[0]), .A2(n431), .ZN(
        cell_1943_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1943_a_HPC2_and_U5 ( .A(cell_1943_a_HPC2_and_n8), .B(
        cell_1943_a_HPC2_and_z_1__1_), .ZN(cell_1943_and_out[1]) );
  XNOR2_X1 cell_1943_a_HPC2_and_U4 ( .A(
        cell_1943_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1943_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1943_a_HPC2_and_n8) );
  XNOR2_X1 cell_1943_a_HPC2_and_U3 ( .A(cell_1943_a_HPC2_and_n7), .B(
        cell_1943_a_HPC2_and_z_0__0_), .ZN(cell_1943_and_out[0]) );
  XNOR2_X1 cell_1943_a_HPC2_and_U2 ( .A(
        cell_1943_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1943_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1943_a_HPC2_and_n7) );
  DFF_X1 cell_1943_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1943_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1943_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1943_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1943_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1943_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1943_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1943_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1943_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1943_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1944_U4 ( .A(signal_3507), .B(cell_1944_and_out[1]), .Z(
        signal_3722) );
  XOR2_X1 cell_1944_U3 ( .A(signal_2069), .B(cell_1944_and_out[0]), .Z(
        signal_2212) );
  XOR2_X1 cell_1944_U2 ( .A(signal_3507), .B(signal_3428), .Z(
        cell_1944_and_in[1]) );
  XOR2_X1 cell_1944_U1 ( .A(signal_2069), .B(signal_2014), .Z(
        cell_1944_and_in[0]) );
  XOR2_X1 cell_1944_a_HPC2_and_U14 ( .A(Fresh[230]), .B(cell_1944_and_in[0]), 
        .Z(cell_1944_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1944_a_HPC2_and_U13 ( .A(Fresh[230]), .B(cell_1944_and_in[1]), 
        .Z(cell_1944_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1944_a_HPC2_and_U12 ( .A1(cell_1944_a_HPC2_and_a_reg[1]), .A2(
        cell_1944_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1944_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1944_a_HPC2_and_U11 ( .A1(cell_1944_a_HPC2_and_a_reg[0]), .A2(
        cell_1944_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1944_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1944_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1944_a_HPC2_and_n9), 
        .ZN(cell_1944_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1944_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1944_a_HPC2_and_n9), 
        .ZN(cell_1944_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1944_a_HPC2_and_U8 ( .A(Fresh[230]), .ZN(cell_1944_a_HPC2_and_n9) );
  AND2_X1 cell_1944_a_HPC2_and_U7 ( .A1(cell_1944_and_in[1]), .A2(n445), .ZN(
        cell_1944_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1944_a_HPC2_and_U6 ( .A1(cell_1944_and_in[0]), .A2(n431), .ZN(
        cell_1944_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1944_a_HPC2_and_U5 ( .A(cell_1944_a_HPC2_and_n8), .B(
        cell_1944_a_HPC2_and_z_1__1_), .ZN(cell_1944_and_out[1]) );
  XNOR2_X1 cell_1944_a_HPC2_and_U4 ( .A(
        cell_1944_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1944_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1944_a_HPC2_and_n8) );
  XNOR2_X1 cell_1944_a_HPC2_and_U3 ( .A(cell_1944_a_HPC2_and_n7), .B(
        cell_1944_a_HPC2_and_z_0__0_), .ZN(cell_1944_and_out[0]) );
  XNOR2_X1 cell_1944_a_HPC2_and_U2 ( .A(
        cell_1944_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1944_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1944_a_HPC2_and_n7) );
  DFF_X1 cell_1944_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1944_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1944_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1944_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1944_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1944_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1944_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1944_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1944_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1944_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1945_U4 ( .A(signal_3519), .B(cell_1945_and_out[1]), .Z(
        signal_3723) );
  XOR2_X1 cell_1945_U3 ( .A(signal_2081), .B(cell_1945_and_out[0]), .Z(
        signal_2213) );
  XOR2_X1 cell_1945_U2 ( .A(signal_3519), .B(signal_3419), .Z(
        cell_1945_and_in[1]) );
  XOR2_X1 cell_1945_U1 ( .A(signal_2081), .B(signal_2005), .Z(
        cell_1945_and_in[0]) );
  XOR2_X1 cell_1945_a_HPC2_and_U14 ( .A(Fresh[231]), .B(cell_1945_and_in[0]), 
        .Z(cell_1945_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1945_a_HPC2_and_U13 ( .A(Fresh[231]), .B(cell_1945_and_in[1]), 
        .Z(cell_1945_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1945_a_HPC2_and_U12 ( .A1(cell_1945_a_HPC2_and_a_reg[1]), .A2(
        cell_1945_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1945_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1945_a_HPC2_and_U11 ( .A1(cell_1945_a_HPC2_and_a_reg[0]), .A2(
        cell_1945_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1945_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1945_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1945_a_HPC2_and_n9), 
        .ZN(cell_1945_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1945_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1945_a_HPC2_and_n9), 
        .ZN(cell_1945_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1945_a_HPC2_and_U8 ( .A(Fresh[231]), .ZN(cell_1945_a_HPC2_and_n9) );
  AND2_X1 cell_1945_a_HPC2_and_U7 ( .A1(cell_1945_and_in[1]), .A2(n453), .ZN(
        cell_1945_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1945_a_HPC2_and_U6 ( .A1(cell_1945_and_in[0]), .A2(n439), .ZN(
        cell_1945_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1945_a_HPC2_and_U5 ( .A(cell_1945_a_HPC2_and_n8), .B(
        cell_1945_a_HPC2_and_z_1__1_), .ZN(cell_1945_and_out[1]) );
  XNOR2_X1 cell_1945_a_HPC2_and_U4 ( .A(
        cell_1945_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1945_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1945_a_HPC2_and_n8) );
  XNOR2_X1 cell_1945_a_HPC2_and_U3 ( .A(cell_1945_a_HPC2_and_n7), .B(
        cell_1945_a_HPC2_and_z_0__0_), .ZN(cell_1945_and_out[0]) );
  XNOR2_X1 cell_1945_a_HPC2_and_U2 ( .A(
        cell_1945_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1945_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1945_a_HPC2_and_n7) );
  DFF_X1 cell_1945_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1945_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1945_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1945_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1945_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1945_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1945_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1945_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1945_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1945_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1946_U4 ( .A(1'b0), .B(cell_1946_and_out[1]), .Z(signal_3724)
         );
  XOR2_X1 cell_1946_U3 ( .A(1'b1), .B(cell_1946_and_out[0]), .Z(signal_2214)
         );
  XOR2_X1 cell_1946_U2 ( .A(1'b0), .B(signal_3571), .Z(cell_1946_and_in[1]) );
  XOR2_X1 cell_1946_U1 ( .A(1'b1), .B(signal_2133), .Z(cell_1946_and_in[0]) );
  XOR2_X1 cell_1946_a_HPC2_and_U14 ( .A(Fresh[232]), .B(cell_1946_and_in[0]), 
        .Z(cell_1946_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1946_a_HPC2_and_U13 ( .A(Fresh[232]), .B(cell_1946_and_in[1]), 
        .Z(cell_1946_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1946_a_HPC2_and_U12 ( .A1(cell_1946_a_HPC2_and_a_reg[1]), .A2(
        cell_1946_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1946_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1946_a_HPC2_and_U11 ( .A1(cell_1946_a_HPC2_and_a_reg[0]), .A2(
        cell_1946_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1946_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1946_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1946_a_HPC2_and_n9), 
        .ZN(cell_1946_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1946_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1946_a_HPC2_and_n9), 
        .ZN(cell_1946_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1946_a_HPC2_and_U8 ( .A(Fresh[232]), .ZN(cell_1946_a_HPC2_and_n9) );
  AND2_X1 cell_1946_a_HPC2_and_U7 ( .A1(cell_1946_and_in[1]), .A2(n453), .ZN(
        cell_1946_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1946_a_HPC2_and_U6 ( .A1(cell_1946_and_in[0]), .A2(n439), .ZN(
        cell_1946_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1946_a_HPC2_and_U5 ( .A(cell_1946_a_HPC2_and_n8), .B(
        cell_1946_a_HPC2_and_z_1__1_), .ZN(cell_1946_and_out[1]) );
  XNOR2_X1 cell_1946_a_HPC2_and_U4 ( .A(
        cell_1946_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1946_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1946_a_HPC2_and_n8) );
  XNOR2_X1 cell_1946_a_HPC2_and_U3 ( .A(cell_1946_a_HPC2_and_n7), .B(
        cell_1946_a_HPC2_and_z_0__0_), .ZN(cell_1946_and_out[0]) );
  XNOR2_X1 cell_1946_a_HPC2_and_U2 ( .A(
        cell_1946_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1946_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1946_a_HPC2_and_n7) );
  DFF_X1 cell_1946_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1946_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1946_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1946_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1946_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1946_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1946_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1946_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1946_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1946_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1947_U4 ( .A(signal_3497), .B(cell_1947_and_out[1]), .Z(
        signal_3725) );
  XOR2_X1 cell_1947_U3 ( .A(signal_2059), .B(cell_1947_and_out[0]), .Z(
        signal_2215) );
  XOR2_X1 cell_1947_U2 ( .A(signal_3497), .B(signal_3260), .Z(
        cell_1947_and_in[1]) );
  XOR2_X1 cell_1947_U1 ( .A(signal_2059), .B(signal_1986), .Z(
        cell_1947_and_in[0]) );
  XOR2_X1 cell_1947_a_HPC2_and_U14 ( .A(Fresh[233]), .B(cell_1947_and_in[0]), 
        .Z(cell_1947_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1947_a_HPC2_and_U13 ( .A(Fresh[233]), .B(cell_1947_and_in[1]), 
        .Z(cell_1947_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1947_a_HPC2_and_U12 ( .A1(cell_1947_a_HPC2_and_a_reg[1]), .A2(
        cell_1947_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1947_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1947_a_HPC2_and_U11 ( .A1(cell_1947_a_HPC2_and_a_reg[0]), .A2(
        cell_1947_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1947_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1947_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1947_a_HPC2_and_n9), 
        .ZN(cell_1947_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1947_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1947_a_HPC2_and_n9), 
        .ZN(cell_1947_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1947_a_HPC2_and_U8 ( .A(Fresh[233]), .ZN(cell_1947_a_HPC2_and_n9) );
  AND2_X1 cell_1947_a_HPC2_and_U7 ( .A1(cell_1947_and_in[1]), .A2(n453), .ZN(
        cell_1947_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1947_a_HPC2_and_U6 ( .A1(cell_1947_and_in[0]), .A2(n439), .ZN(
        cell_1947_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1947_a_HPC2_and_U5 ( .A(cell_1947_a_HPC2_and_n8), .B(
        cell_1947_a_HPC2_and_z_1__1_), .ZN(cell_1947_and_out[1]) );
  XNOR2_X1 cell_1947_a_HPC2_and_U4 ( .A(
        cell_1947_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1947_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1947_a_HPC2_and_n8) );
  XNOR2_X1 cell_1947_a_HPC2_and_U3 ( .A(cell_1947_a_HPC2_and_n7), .B(
        cell_1947_a_HPC2_and_z_0__0_), .ZN(cell_1947_and_out[0]) );
  XNOR2_X1 cell_1947_a_HPC2_and_U2 ( .A(
        cell_1947_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1947_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1947_a_HPC2_and_n7) );
  DFF_X1 cell_1947_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1947_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1947_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1947_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1947_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1947_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1947_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1947_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1947_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1947_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1948_U4 ( .A(signal_3476), .B(cell_1948_and_out[1]), .Z(
        signal_3726) );
  XOR2_X1 cell_1948_U3 ( .A(signal_2038), .B(cell_1948_and_out[0]), .Z(
        signal_2216) );
  XOR2_X1 cell_1948_U2 ( .A(signal_3476), .B(signal_3258), .Z(
        cell_1948_and_in[1]) );
  XOR2_X1 cell_1948_U1 ( .A(signal_2038), .B(signal_1984), .Z(
        cell_1948_and_in[0]) );
  XOR2_X1 cell_1948_a_HPC2_and_U14 ( .A(Fresh[234]), .B(cell_1948_and_in[0]), 
        .Z(cell_1948_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1948_a_HPC2_and_U13 ( .A(Fresh[234]), .B(cell_1948_and_in[1]), 
        .Z(cell_1948_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1948_a_HPC2_and_U12 ( .A1(cell_1948_a_HPC2_and_a_reg[1]), .A2(
        cell_1948_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1948_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1948_a_HPC2_and_U11 ( .A1(cell_1948_a_HPC2_and_a_reg[0]), .A2(
        cell_1948_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1948_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1948_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1948_a_HPC2_and_n9), 
        .ZN(cell_1948_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1948_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1948_a_HPC2_and_n9), 
        .ZN(cell_1948_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1948_a_HPC2_and_U8 ( .A(Fresh[234]), .ZN(cell_1948_a_HPC2_and_n9) );
  AND2_X1 cell_1948_a_HPC2_and_U7 ( .A1(cell_1948_and_in[1]), .A2(n445), .ZN(
        cell_1948_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1948_a_HPC2_and_U6 ( .A1(cell_1948_and_in[0]), .A2(n431), .ZN(
        cell_1948_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1948_a_HPC2_and_U5 ( .A(cell_1948_a_HPC2_and_n8), .B(
        cell_1948_a_HPC2_and_z_1__1_), .ZN(cell_1948_and_out[1]) );
  XNOR2_X1 cell_1948_a_HPC2_and_U4 ( .A(
        cell_1948_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1948_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1948_a_HPC2_and_n8) );
  XNOR2_X1 cell_1948_a_HPC2_and_U3 ( .A(cell_1948_a_HPC2_and_n7), .B(
        cell_1948_a_HPC2_and_z_0__0_), .ZN(cell_1948_and_out[0]) );
  XNOR2_X1 cell_1948_a_HPC2_and_U2 ( .A(
        cell_1948_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1948_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1948_a_HPC2_and_n7) );
  DFF_X1 cell_1948_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1948_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1948_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1948_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1948_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1948_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1948_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1948_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1948_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1948_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1949_U4 ( .A(signal_3511), .B(cell_1949_and_out[1]), .Z(
        signal_3727) );
  XOR2_X1 cell_1949_U3 ( .A(signal_2073), .B(cell_1949_and_out[0]), .Z(
        signal_2217) );
  XOR2_X1 cell_1949_U2 ( .A(signal_3511), .B(signal_3560), .Z(
        cell_1949_and_in[1]) );
  XOR2_X1 cell_1949_U1 ( .A(signal_2073), .B(signal_2122), .Z(
        cell_1949_and_in[0]) );
  XOR2_X1 cell_1949_a_HPC2_and_U14 ( .A(Fresh[235]), .B(cell_1949_and_in[0]), 
        .Z(cell_1949_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1949_a_HPC2_and_U13 ( .A(Fresh[235]), .B(cell_1949_and_in[1]), 
        .Z(cell_1949_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1949_a_HPC2_and_U12 ( .A1(cell_1949_a_HPC2_and_a_reg[1]), .A2(
        cell_1949_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1949_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1949_a_HPC2_and_U11 ( .A1(cell_1949_a_HPC2_and_a_reg[0]), .A2(
        cell_1949_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1949_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1949_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1949_a_HPC2_and_n9), 
        .ZN(cell_1949_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1949_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1949_a_HPC2_and_n9), 
        .ZN(cell_1949_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1949_a_HPC2_and_U8 ( .A(Fresh[235]), .ZN(cell_1949_a_HPC2_and_n9) );
  AND2_X1 cell_1949_a_HPC2_and_U7 ( .A1(cell_1949_and_in[1]), .A2(n445), .ZN(
        cell_1949_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1949_a_HPC2_and_U6 ( .A1(cell_1949_and_in[0]), .A2(n431), .ZN(
        cell_1949_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1949_a_HPC2_and_U5 ( .A(cell_1949_a_HPC2_and_n8), .B(
        cell_1949_a_HPC2_and_z_1__1_), .ZN(cell_1949_and_out[1]) );
  XNOR2_X1 cell_1949_a_HPC2_and_U4 ( .A(
        cell_1949_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1949_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1949_a_HPC2_and_n8) );
  XNOR2_X1 cell_1949_a_HPC2_and_U3 ( .A(cell_1949_a_HPC2_and_n7), .B(
        cell_1949_a_HPC2_and_z_0__0_), .ZN(cell_1949_and_out[0]) );
  XNOR2_X1 cell_1949_a_HPC2_and_U2 ( .A(
        cell_1949_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1949_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1949_a_HPC2_and_n7) );
  DFF_X1 cell_1949_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1949_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1949_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1949_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1949_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1949_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1949_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1949_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1949_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1949_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1950_U4 ( .A(signal_3259), .B(cell_1950_and_out[1]), .Z(
        signal_3728) );
  XOR2_X1 cell_1950_U3 ( .A(signal_1985), .B(cell_1950_and_out[0]), .Z(
        signal_2218) );
  XOR2_X1 cell_1950_U2 ( .A(signal_3259), .B(signal_3509), .Z(
        cell_1950_and_in[1]) );
  XOR2_X1 cell_1950_U1 ( .A(signal_1985), .B(signal_2071), .Z(
        cell_1950_and_in[0]) );
  XOR2_X1 cell_1950_a_HPC2_and_U14 ( .A(Fresh[236]), .B(cell_1950_and_in[0]), 
        .Z(cell_1950_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1950_a_HPC2_and_U13 ( .A(Fresh[236]), .B(cell_1950_and_in[1]), 
        .Z(cell_1950_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1950_a_HPC2_and_U12 ( .A1(cell_1950_a_HPC2_and_a_reg[1]), .A2(
        cell_1950_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1950_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1950_a_HPC2_and_U11 ( .A1(cell_1950_a_HPC2_and_a_reg[0]), .A2(
        cell_1950_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1950_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1950_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1950_a_HPC2_and_n9), 
        .ZN(cell_1950_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1950_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1950_a_HPC2_and_n9), 
        .ZN(cell_1950_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1950_a_HPC2_and_U8 ( .A(Fresh[236]), .ZN(cell_1950_a_HPC2_and_n9) );
  AND2_X1 cell_1950_a_HPC2_and_U7 ( .A1(cell_1950_and_in[1]), .A2(n446), .ZN(
        cell_1950_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1950_a_HPC2_and_U6 ( .A1(cell_1950_and_in[0]), .A2(n432), .ZN(
        cell_1950_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1950_a_HPC2_and_U5 ( .A(cell_1950_a_HPC2_and_n8), .B(
        cell_1950_a_HPC2_and_z_1__1_), .ZN(cell_1950_and_out[1]) );
  XNOR2_X1 cell_1950_a_HPC2_and_U4 ( .A(
        cell_1950_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1950_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1950_a_HPC2_and_n8) );
  XNOR2_X1 cell_1950_a_HPC2_and_U3 ( .A(cell_1950_a_HPC2_and_n7), .B(
        cell_1950_a_HPC2_and_z_0__0_), .ZN(cell_1950_and_out[0]) );
  XNOR2_X1 cell_1950_a_HPC2_and_U2 ( .A(
        cell_1950_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1950_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1950_a_HPC2_and_n7) );
  DFF_X1 cell_1950_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1950_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1950_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1950_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1950_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1950_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1950_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1950_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1950_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1950_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1951_U4 ( .A(signal_3564), .B(cell_1951_and_out[1]), .Z(
        signal_3729) );
  XOR2_X1 cell_1951_U3 ( .A(signal_2126), .B(cell_1951_and_out[0]), .Z(
        signal_2219) );
  XOR2_X1 cell_1951_U2 ( .A(signal_3564), .B(signal_3412), .Z(
        cell_1951_and_in[1]) );
  XOR2_X1 cell_1951_U1 ( .A(signal_2126), .B(signal_1998), .Z(
        cell_1951_and_in[0]) );
  XOR2_X1 cell_1951_a_HPC2_and_U14 ( .A(Fresh[237]), .B(cell_1951_and_in[0]), 
        .Z(cell_1951_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1951_a_HPC2_and_U13 ( .A(Fresh[237]), .B(cell_1951_and_in[1]), 
        .Z(cell_1951_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1951_a_HPC2_and_U12 ( .A1(cell_1951_a_HPC2_and_a_reg[1]), .A2(
        cell_1951_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1951_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1951_a_HPC2_and_U11 ( .A1(cell_1951_a_HPC2_and_a_reg[0]), .A2(
        cell_1951_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1951_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1951_a_HPC2_and_U10 ( .A1(n453), .A2(cell_1951_a_HPC2_and_n9), 
        .ZN(cell_1951_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1951_a_HPC2_and_U9 ( .A1(n439), .A2(cell_1951_a_HPC2_and_n9), 
        .ZN(cell_1951_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1951_a_HPC2_and_U8 ( .A(Fresh[237]), .ZN(cell_1951_a_HPC2_and_n9) );
  AND2_X1 cell_1951_a_HPC2_and_U7 ( .A1(cell_1951_and_in[1]), .A2(n453), .ZN(
        cell_1951_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1951_a_HPC2_and_U6 ( .A1(cell_1951_and_in[0]), .A2(n439), .ZN(
        cell_1951_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1951_a_HPC2_and_U5 ( .A(cell_1951_a_HPC2_and_n8), .B(
        cell_1951_a_HPC2_and_z_1__1_), .ZN(cell_1951_and_out[1]) );
  XNOR2_X1 cell_1951_a_HPC2_and_U4 ( .A(
        cell_1951_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1951_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1951_a_HPC2_and_n8) );
  XNOR2_X1 cell_1951_a_HPC2_and_U3 ( .A(cell_1951_a_HPC2_and_n7), .B(
        cell_1951_a_HPC2_and_z_0__0_), .ZN(cell_1951_and_out[0]) );
  XNOR2_X1 cell_1951_a_HPC2_and_U2 ( .A(
        cell_1951_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1951_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1951_a_HPC2_and_n7) );
  DFF_X1 cell_1951_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1951_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1951_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n439), .CK(clk), 
        .Q(cell_1951_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1951_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1951_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n453), .CK(clk), 
        .Q(cell_1951_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1951_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1951_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1951_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1952_U4 ( .A(signal_3557), .B(cell_1952_and_out[1]), .Z(
        signal_3730) );
  XOR2_X1 cell_1952_U3 ( .A(signal_2119), .B(cell_1952_and_out[0]), .Z(
        signal_2220) );
  XOR2_X1 cell_1952_U2 ( .A(signal_3557), .B(signal_3520), .Z(
        cell_1952_and_in[1]) );
  XOR2_X1 cell_1952_U1 ( .A(signal_2119), .B(signal_2082), .Z(
        cell_1952_and_in[0]) );
  XOR2_X1 cell_1952_a_HPC2_and_U14 ( .A(Fresh[238]), .B(cell_1952_and_in[0]), 
        .Z(cell_1952_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1952_a_HPC2_and_U13 ( .A(Fresh[238]), .B(cell_1952_and_in[1]), 
        .Z(cell_1952_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1952_a_HPC2_and_U12 ( .A1(cell_1952_a_HPC2_and_a_reg[1]), .A2(
        cell_1952_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1952_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1952_a_HPC2_and_U11 ( .A1(cell_1952_a_HPC2_and_a_reg[0]), .A2(
        cell_1952_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1952_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1952_a_HPC2_and_U10 ( .A1(n445), .A2(cell_1952_a_HPC2_and_n9), 
        .ZN(cell_1952_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1952_a_HPC2_and_U9 ( .A1(n431), .A2(cell_1952_a_HPC2_and_n9), 
        .ZN(cell_1952_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1952_a_HPC2_and_U8 ( .A(Fresh[238]), .ZN(cell_1952_a_HPC2_and_n9) );
  AND2_X1 cell_1952_a_HPC2_and_U7 ( .A1(cell_1952_and_in[1]), .A2(n445), .ZN(
        cell_1952_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1952_a_HPC2_and_U6 ( .A1(cell_1952_and_in[0]), .A2(n431), .ZN(
        cell_1952_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1952_a_HPC2_and_U5 ( .A(cell_1952_a_HPC2_and_n8), .B(
        cell_1952_a_HPC2_and_z_1__1_), .ZN(cell_1952_and_out[1]) );
  XNOR2_X1 cell_1952_a_HPC2_and_U4 ( .A(
        cell_1952_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1952_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1952_a_HPC2_and_n8) );
  XNOR2_X1 cell_1952_a_HPC2_and_U3 ( .A(cell_1952_a_HPC2_and_n7), .B(
        cell_1952_a_HPC2_and_z_0__0_), .ZN(cell_1952_and_out[0]) );
  XNOR2_X1 cell_1952_a_HPC2_and_U2 ( .A(
        cell_1952_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1952_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1952_a_HPC2_and_n7) );
  DFF_X1 cell_1952_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1952_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1952_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n431), .CK(clk), 
        .Q(cell_1952_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1952_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1952_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n445), .CK(clk), 
        .Q(cell_1952_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1952_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1952_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1952_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1953_U4 ( .A(signal_3497), .B(cell_1953_and_out[1]), .Z(
        signal_3731) );
  XOR2_X1 cell_1953_U3 ( .A(signal_2059), .B(cell_1953_and_out[0]), .Z(
        signal_2221) );
  XOR2_X1 cell_1953_U2 ( .A(signal_3497), .B(signal_3589), .Z(
        cell_1953_and_in[1]) );
  XOR2_X1 cell_1953_U1 ( .A(signal_2059), .B(signal_2151), .Z(
        cell_1953_and_in[0]) );
  XOR2_X1 cell_1953_a_HPC2_and_U14 ( .A(Fresh[239]), .B(cell_1953_and_in[0]), 
        .Z(cell_1953_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1953_a_HPC2_and_U13 ( .A(Fresh[239]), .B(cell_1953_and_in[1]), 
        .Z(cell_1953_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1953_a_HPC2_and_U12 ( .A1(cell_1953_a_HPC2_and_a_reg[1]), .A2(
        cell_1953_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1953_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1953_a_HPC2_and_U11 ( .A1(cell_1953_a_HPC2_and_a_reg[0]), .A2(
        cell_1953_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1953_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1953_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1953_a_HPC2_and_n9), 
        .ZN(cell_1953_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1953_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1953_a_HPC2_and_n9), 
        .ZN(cell_1953_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1953_a_HPC2_and_U8 ( .A(Fresh[239]), .ZN(cell_1953_a_HPC2_and_n9) );
  AND2_X1 cell_1953_a_HPC2_and_U7 ( .A1(cell_1953_and_in[1]), .A2(n446), .ZN(
        cell_1953_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1953_a_HPC2_and_U6 ( .A1(cell_1953_and_in[0]), .A2(n432), .ZN(
        cell_1953_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1953_a_HPC2_and_U5 ( .A(cell_1953_a_HPC2_and_n8), .B(
        cell_1953_a_HPC2_and_z_1__1_), .ZN(cell_1953_and_out[1]) );
  XNOR2_X1 cell_1953_a_HPC2_and_U4 ( .A(
        cell_1953_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1953_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1953_a_HPC2_and_n8) );
  XNOR2_X1 cell_1953_a_HPC2_and_U3 ( .A(cell_1953_a_HPC2_and_n7), .B(
        cell_1953_a_HPC2_and_z_0__0_), .ZN(cell_1953_and_out[0]) );
  XNOR2_X1 cell_1953_a_HPC2_and_U2 ( .A(
        cell_1953_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1953_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1953_a_HPC2_and_n7) );
  DFF_X1 cell_1953_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1953_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1953_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1953_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1953_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1953_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1953_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1953_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1953_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1953_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1954_U4 ( .A(signal_3525), .B(cell_1954_and_out[1]), .Z(
        signal_3732) );
  XOR2_X1 cell_1954_U3 ( .A(signal_2087), .B(cell_1954_and_out[0]), .Z(
        signal_2222) );
  XOR2_X1 cell_1954_U2 ( .A(signal_3525), .B(n371), .Z(cell_1954_and_in[1]) );
  XOR2_X1 cell_1954_U1 ( .A(signal_2087), .B(n369), .Z(cell_1954_and_in[0]) );
  XOR2_X1 cell_1954_a_HPC2_and_U14 ( .A(Fresh[240]), .B(cell_1954_and_in[0]), 
        .Z(cell_1954_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1954_a_HPC2_and_U13 ( .A(Fresh[240]), .B(cell_1954_and_in[1]), 
        .Z(cell_1954_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1954_a_HPC2_and_U12 ( .A1(cell_1954_a_HPC2_and_a_reg[1]), .A2(
        cell_1954_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1954_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1954_a_HPC2_and_U11 ( .A1(cell_1954_a_HPC2_and_a_reg[0]), .A2(
        cell_1954_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1954_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1954_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1954_a_HPC2_and_n9), 
        .ZN(cell_1954_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1954_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1954_a_HPC2_and_n9), 
        .ZN(cell_1954_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1954_a_HPC2_and_U8 ( .A(Fresh[240]), .ZN(cell_1954_a_HPC2_and_n9) );
  AND2_X1 cell_1954_a_HPC2_and_U7 ( .A1(cell_1954_and_in[1]), .A2(n446), .ZN(
        cell_1954_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1954_a_HPC2_and_U6 ( .A1(cell_1954_and_in[0]), .A2(n432), .ZN(
        cell_1954_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1954_a_HPC2_and_U5 ( .A(cell_1954_a_HPC2_and_n8), .B(
        cell_1954_a_HPC2_and_z_1__1_), .ZN(cell_1954_and_out[1]) );
  XNOR2_X1 cell_1954_a_HPC2_and_U4 ( .A(
        cell_1954_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1954_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1954_a_HPC2_and_n8) );
  XNOR2_X1 cell_1954_a_HPC2_and_U3 ( .A(cell_1954_a_HPC2_and_n7), .B(
        cell_1954_a_HPC2_and_z_0__0_), .ZN(cell_1954_and_out[0]) );
  XNOR2_X1 cell_1954_a_HPC2_and_U2 ( .A(
        cell_1954_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1954_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1954_a_HPC2_and_n7) );
  DFF_X1 cell_1954_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1954_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1954_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1954_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1954_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1954_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1954_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1954_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1954_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1954_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1955_U4 ( .A(signal_3533), .B(cell_1955_and_out[1]), .Z(
        signal_3733) );
  XOR2_X1 cell_1955_U3 ( .A(signal_2095), .B(cell_1955_and_out[0]), .Z(
        signal_2223) );
  XOR2_X1 cell_1955_U2 ( .A(signal_3533), .B(signal_3415), .Z(
        cell_1955_and_in[1]) );
  XOR2_X1 cell_1955_U1 ( .A(signal_2095), .B(signal_2001), .Z(
        cell_1955_and_in[0]) );
  XOR2_X1 cell_1955_a_HPC2_and_U14 ( .A(Fresh[241]), .B(cell_1955_and_in[0]), 
        .Z(cell_1955_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1955_a_HPC2_and_U13 ( .A(Fresh[241]), .B(cell_1955_and_in[1]), 
        .Z(cell_1955_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1955_a_HPC2_and_U12 ( .A1(cell_1955_a_HPC2_and_a_reg[1]), .A2(
        cell_1955_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1955_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1955_a_HPC2_and_U11 ( .A1(cell_1955_a_HPC2_and_a_reg[0]), .A2(
        cell_1955_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1955_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1955_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1955_a_HPC2_and_n9), 
        .ZN(cell_1955_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1955_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1955_a_HPC2_and_n9), 
        .ZN(cell_1955_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1955_a_HPC2_and_U8 ( .A(Fresh[241]), .ZN(cell_1955_a_HPC2_and_n9) );
  AND2_X1 cell_1955_a_HPC2_and_U7 ( .A1(cell_1955_and_in[1]), .A2(n446), .ZN(
        cell_1955_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1955_a_HPC2_and_U6 ( .A1(cell_1955_and_in[0]), .A2(n432), .ZN(
        cell_1955_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1955_a_HPC2_and_U5 ( .A(cell_1955_a_HPC2_and_n8), .B(
        cell_1955_a_HPC2_and_z_1__1_), .ZN(cell_1955_and_out[1]) );
  XNOR2_X1 cell_1955_a_HPC2_and_U4 ( .A(
        cell_1955_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1955_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1955_a_HPC2_and_n8) );
  XNOR2_X1 cell_1955_a_HPC2_and_U3 ( .A(cell_1955_a_HPC2_and_n7), .B(
        cell_1955_a_HPC2_and_z_0__0_), .ZN(cell_1955_and_out[0]) );
  XNOR2_X1 cell_1955_a_HPC2_and_U2 ( .A(
        cell_1955_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1955_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1955_a_HPC2_and_n7) );
  DFF_X1 cell_1955_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1955_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1955_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1955_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1955_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1955_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1955_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1955_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1955_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1955_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1956_U4 ( .A(signal_3558), .B(cell_1956_and_out[1]), .Z(
        signal_3734) );
  XOR2_X1 cell_1956_U3 ( .A(signal_2120), .B(cell_1956_and_out[0]), .Z(
        signal_2224) );
  XOR2_X1 cell_1956_U2 ( .A(signal_3558), .B(signal_3551), .Z(
        cell_1956_and_in[1]) );
  XOR2_X1 cell_1956_U1 ( .A(signal_2120), .B(signal_2113), .Z(
        cell_1956_and_in[0]) );
  XOR2_X1 cell_1956_a_HPC2_and_U14 ( .A(Fresh[242]), .B(cell_1956_and_in[0]), 
        .Z(cell_1956_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1956_a_HPC2_and_U13 ( .A(Fresh[242]), .B(cell_1956_and_in[1]), 
        .Z(cell_1956_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1956_a_HPC2_and_U12 ( .A1(cell_1956_a_HPC2_and_a_reg[1]), .A2(
        cell_1956_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1956_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1956_a_HPC2_and_U11 ( .A1(cell_1956_a_HPC2_and_a_reg[0]), .A2(
        cell_1956_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1956_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1956_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1956_a_HPC2_and_n9), 
        .ZN(cell_1956_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1956_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1956_a_HPC2_and_n9), 
        .ZN(cell_1956_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1956_a_HPC2_and_U8 ( .A(Fresh[242]), .ZN(cell_1956_a_HPC2_and_n9) );
  AND2_X1 cell_1956_a_HPC2_and_U7 ( .A1(cell_1956_and_in[1]), .A2(n447), .ZN(
        cell_1956_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1956_a_HPC2_and_U6 ( .A1(cell_1956_and_in[0]), .A2(n433), .ZN(
        cell_1956_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1956_a_HPC2_and_U5 ( .A(cell_1956_a_HPC2_and_n8), .B(
        cell_1956_a_HPC2_and_z_1__1_), .ZN(cell_1956_and_out[1]) );
  XNOR2_X1 cell_1956_a_HPC2_and_U4 ( .A(
        cell_1956_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1956_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1956_a_HPC2_and_n8) );
  XNOR2_X1 cell_1956_a_HPC2_and_U3 ( .A(cell_1956_a_HPC2_and_n7), .B(
        cell_1956_a_HPC2_and_z_0__0_), .ZN(cell_1956_and_out[0]) );
  XNOR2_X1 cell_1956_a_HPC2_and_U2 ( .A(
        cell_1956_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1956_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1956_a_HPC2_and_n7) );
  DFF_X1 cell_1956_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1956_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1956_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1956_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1956_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1956_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1956_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1956_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1956_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1956_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1957_U4 ( .A(signal_3584), .B(cell_1957_and_out[1]), .Z(
        signal_3735) );
  XOR2_X1 cell_1957_U3 ( .A(signal_2146), .B(cell_1957_and_out[0]), .Z(
        signal_2225) );
  XOR2_X1 cell_1957_U2 ( .A(signal_3584), .B(signal_3430), .Z(
        cell_1957_and_in[1]) );
  XOR2_X1 cell_1957_U1 ( .A(signal_2146), .B(signal_2016), .Z(
        cell_1957_and_in[0]) );
  XOR2_X1 cell_1957_a_HPC2_and_U14 ( .A(Fresh[243]), .B(cell_1957_and_in[0]), 
        .Z(cell_1957_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1957_a_HPC2_and_U13 ( .A(Fresh[243]), .B(cell_1957_and_in[1]), 
        .Z(cell_1957_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1957_a_HPC2_and_U12 ( .A1(cell_1957_a_HPC2_and_a_reg[1]), .A2(
        cell_1957_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1957_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1957_a_HPC2_and_U11 ( .A1(cell_1957_a_HPC2_and_a_reg[0]), .A2(
        cell_1957_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1957_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1957_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1957_a_HPC2_and_n9), 
        .ZN(cell_1957_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1957_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1957_a_HPC2_and_n9), 
        .ZN(cell_1957_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1957_a_HPC2_and_U8 ( .A(Fresh[243]), .ZN(cell_1957_a_HPC2_and_n9) );
  AND2_X1 cell_1957_a_HPC2_and_U7 ( .A1(cell_1957_and_in[1]), .A2(n448), .ZN(
        cell_1957_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1957_a_HPC2_and_U6 ( .A1(cell_1957_and_in[0]), .A2(n434), .ZN(
        cell_1957_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1957_a_HPC2_and_U5 ( .A(cell_1957_a_HPC2_and_n8), .B(
        cell_1957_a_HPC2_and_z_1__1_), .ZN(cell_1957_and_out[1]) );
  XNOR2_X1 cell_1957_a_HPC2_and_U4 ( .A(
        cell_1957_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1957_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1957_a_HPC2_and_n8) );
  XNOR2_X1 cell_1957_a_HPC2_and_U3 ( .A(cell_1957_a_HPC2_and_n7), .B(
        cell_1957_a_HPC2_and_z_0__0_), .ZN(cell_1957_and_out[0]) );
  XNOR2_X1 cell_1957_a_HPC2_and_U2 ( .A(
        cell_1957_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1957_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1957_a_HPC2_and_n7) );
  DFF_X1 cell_1957_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1957_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1957_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1957_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1957_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1957_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1957_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1957_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1957_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1957_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1958_U4 ( .A(signal_3474), .B(cell_1958_and_out[1]), .Z(
        signal_3736) );
  XOR2_X1 cell_1958_U3 ( .A(signal_2036), .B(cell_1958_and_out[0]), .Z(
        signal_2226) );
  XOR2_X1 cell_1958_U2 ( .A(signal_3474), .B(signal_3413), .Z(
        cell_1958_and_in[1]) );
  XOR2_X1 cell_1958_U1 ( .A(signal_2036), .B(signal_1999), .Z(
        cell_1958_and_in[0]) );
  XOR2_X1 cell_1958_a_HPC2_and_U14 ( .A(Fresh[244]), .B(cell_1958_and_in[0]), 
        .Z(cell_1958_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1958_a_HPC2_and_U13 ( .A(Fresh[244]), .B(cell_1958_and_in[1]), 
        .Z(cell_1958_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1958_a_HPC2_and_U12 ( .A1(cell_1958_a_HPC2_and_a_reg[1]), .A2(
        cell_1958_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1958_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1958_a_HPC2_and_U11 ( .A1(cell_1958_a_HPC2_and_a_reg[0]), .A2(
        cell_1958_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1958_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1958_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1958_a_HPC2_and_n9), 
        .ZN(cell_1958_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1958_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1958_a_HPC2_and_n9), 
        .ZN(cell_1958_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1958_a_HPC2_and_U8 ( .A(Fresh[244]), .ZN(cell_1958_a_HPC2_and_n9) );
  AND2_X1 cell_1958_a_HPC2_and_U7 ( .A1(cell_1958_and_in[1]), .A2(n446), .ZN(
        cell_1958_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1958_a_HPC2_and_U6 ( .A1(cell_1958_and_in[0]), .A2(n432), .ZN(
        cell_1958_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1958_a_HPC2_and_U5 ( .A(cell_1958_a_HPC2_and_n8), .B(
        cell_1958_a_HPC2_and_z_1__1_), .ZN(cell_1958_and_out[1]) );
  XNOR2_X1 cell_1958_a_HPC2_and_U4 ( .A(
        cell_1958_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1958_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1958_a_HPC2_and_n8) );
  XNOR2_X1 cell_1958_a_HPC2_and_U3 ( .A(cell_1958_a_HPC2_and_n7), .B(
        cell_1958_a_HPC2_and_z_0__0_), .ZN(cell_1958_and_out[0]) );
  XNOR2_X1 cell_1958_a_HPC2_and_U2 ( .A(
        cell_1958_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1958_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1958_a_HPC2_and_n7) );
  DFF_X1 cell_1958_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1958_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1958_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1958_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1958_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1958_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1958_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1958_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1958_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1958_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1959_U4 ( .A(signal_3504), .B(cell_1959_and_out[1]), .Z(
        signal_3737) );
  XOR2_X1 cell_1959_U3 ( .A(signal_2066), .B(cell_1959_and_out[0]), .Z(
        signal_2227) );
  XOR2_X1 cell_1959_U2 ( .A(signal_3504), .B(signal_3480), .Z(
        cell_1959_and_in[1]) );
  XOR2_X1 cell_1959_U1 ( .A(signal_2066), .B(signal_2042), .Z(
        cell_1959_and_in[0]) );
  XOR2_X1 cell_1959_a_HPC2_and_U14 ( .A(Fresh[245]), .B(cell_1959_and_in[0]), 
        .Z(cell_1959_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1959_a_HPC2_and_U13 ( .A(Fresh[245]), .B(cell_1959_and_in[1]), 
        .Z(cell_1959_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1959_a_HPC2_and_U12 ( .A1(cell_1959_a_HPC2_and_a_reg[1]), .A2(
        cell_1959_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1959_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1959_a_HPC2_and_U11 ( .A1(cell_1959_a_HPC2_and_a_reg[0]), .A2(
        cell_1959_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1959_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1959_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1959_a_HPC2_and_n9), 
        .ZN(cell_1959_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1959_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1959_a_HPC2_and_n9), 
        .ZN(cell_1959_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1959_a_HPC2_and_U8 ( .A(Fresh[245]), .ZN(cell_1959_a_HPC2_and_n9) );
  AND2_X1 cell_1959_a_HPC2_and_U7 ( .A1(cell_1959_and_in[1]), .A2(n446), .ZN(
        cell_1959_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1959_a_HPC2_and_U6 ( .A1(cell_1959_and_in[0]), .A2(n432), .ZN(
        cell_1959_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1959_a_HPC2_and_U5 ( .A(cell_1959_a_HPC2_and_n8), .B(
        cell_1959_a_HPC2_and_z_1__1_), .ZN(cell_1959_and_out[1]) );
  XNOR2_X1 cell_1959_a_HPC2_and_U4 ( .A(
        cell_1959_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1959_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1959_a_HPC2_and_n8) );
  XNOR2_X1 cell_1959_a_HPC2_and_U3 ( .A(cell_1959_a_HPC2_and_n7), .B(
        cell_1959_a_HPC2_and_z_0__0_), .ZN(cell_1959_and_out[0]) );
  XNOR2_X1 cell_1959_a_HPC2_and_U2 ( .A(
        cell_1959_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1959_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1959_a_HPC2_and_n7) );
  DFF_X1 cell_1959_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1959_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1959_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1959_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1959_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1959_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1959_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1959_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1959_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1959_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1960_U4 ( .A(signal_3526), .B(cell_1960_and_out[1]), .Z(
        signal_3738) );
  XOR2_X1 cell_1960_U3 ( .A(signal_2088), .B(cell_1960_and_out[0]), .Z(
        signal_2228) );
  XOR2_X1 cell_1960_U2 ( .A(signal_3526), .B(signal_3566), .Z(
        cell_1960_and_in[1]) );
  XOR2_X1 cell_1960_U1 ( .A(signal_2088), .B(signal_2128), .Z(
        cell_1960_and_in[0]) );
  XOR2_X1 cell_1960_a_HPC2_and_U14 ( .A(Fresh[246]), .B(cell_1960_and_in[0]), 
        .Z(cell_1960_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1960_a_HPC2_and_U13 ( .A(Fresh[246]), .B(cell_1960_and_in[1]), 
        .Z(cell_1960_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1960_a_HPC2_and_U12 ( .A1(cell_1960_a_HPC2_and_a_reg[1]), .A2(
        cell_1960_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1960_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1960_a_HPC2_and_U11 ( .A1(cell_1960_a_HPC2_and_a_reg[0]), .A2(
        cell_1960_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1960_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1960_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1960_a_HPC2_and_n9), 
        .ZN(cell_1960_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1960_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1960_a_HPC2_and_n9), 
        .ZN(cell_1960_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1960_a_HPC2_and_U8 ( .A(Fresh[246]), .ZN(cell_1960_a_HPC2_and_n9) );
  AND2_X1 cell_1960_a_HPC2_and_U7 ( .A1(cell_1960_and_in[1]), .A2(n446), .ZN(
        cell_1960_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1960_a_HPC2_and_U6 ( .A1(cell_1960_and_in[0]), .A2(n432), .ZN(
        cell_1960_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1960_a_HPC2_and_U5 ( .A(cell_1960_a_HPC2_and_n8), .B(
        cell_1960_a_HPC2_and_z_1__1_), .ZN(cell_1960_and_out[1]) );
  XNOR2_X1 cell_1960_a_HPC2_and_U4 ( .A(
        cell_1960_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1960_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1960_a_HPC2_and_n8) );
  XNOR2_X1 cell_1960_a_HPC2_and_U3 ( .A(cell_1960_a_HPC2_and_n7), .B(
        cell_1960_a_HPC2_and_z_0__0_), .ZN(cell_1960_and_out[0]) );
  XNOR2_X1 cell_1960_a_HPC2_and_U2 ( .A(
        cell_1960_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1960_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1960_a_HPC2_and_n7) );
  DFF_X1 cell_1960_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1960_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1960_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1960_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1960_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1960_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1960_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1960_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1960_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1960_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1961_U4 ( .A(signal_3464), .B(cell_1961_and_out[1]), .Z(
        signal_3739) );
  XOR2_X1 cell_1961_U3 ( .A(signal_2026), .B(cell_1961_and_out[0]), .Z(
        signal_2229) );
  XOR2_X1 cell_1961_U2 ( .A(signal_3464), .B(signal_3538), .Z(
        cell_1961_and_in[1]) );
  XOR2_X1 cell_1961_U1 ( .A(signal_2026), .B(signal_2100), .Z(
        cell_1961_and_in[0]) );
  XOR2_X1 cell_1961_a_HPC2_and_U14 ( .A(Fresh[247]), .B(cell_1961_and_in[0]), 
        .Z(cell_1961_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1961_a_HPC2_and_U13 ( .A(Fresh[247]), .B(cell_1961_and_in[1]), 
        .Z(cell_1961_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1961_a_HPC2_and_U12 ( .A1(cell_1961_a_HPC2_and_a_reg[1]), .A2(
        cell_1961_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1961_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1961_a_HPC2_and_U11 ( .A1(cell_1961_a_HPC2_and_a_reg[0]), .A2(
        cell_1961_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1961_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1961_a_HPC2_and_U10 ( .A1(n446), .A2(cell_1961_a_HPC2_and_n9), 
        .ZN(cell_1961_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1961_a_HPC2_and_U9 ( .A1(n432), .A2(cell_1961_a_HPC2_and_n9), 
        .ZN(cell_1961_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1961_a_HPC2_and_U8 ( .A(Fresh[247]), .ZN(cell_1961_a_HPC2_and_n9) );
  AND2_X1 cell_1961_a_HPC2_and_U7 ( .A1(cell_1961_and_in[1]), .A2(n446), .ZN(
        cell_1961_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1961_a_HPC2_and_U6 ( .A1(cell_1961_and_in[0]), .A2(n432), .ZN(
        cell_1961_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1961_a_HPC2_and_U5 ( .A(cell_1961_a_HPC2_and_n8), .B(
        cell_1961_a_HPC2_and_z_1__1_), .ZN(cell_1961_and_out[1]) );
  XNOR2_X1 cell_1961_a_HPC2_and_U4 ( .A(
        cell_1961_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1961_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1961_a_HPC2_and_n8) );
  XNOR2_X1 cell_1961_a_HPC2_and_U3 ( .A(cell_1961_a_HPC2_and_n7), .B(
        cell_1961_a_HPC2_and_z_0__0_), .ZN(cell_1961_and_out[0]) );
  XNOR2_X1 cell_1961_a_HPC2_and_U2 ( .A(
        cell_1961_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1961_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1961_a_HPC2_and_n7) );
  DFF_X1 cell_1961_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1961_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1961_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n432), .CK(clk), 
        .Q(cell_1961_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1961_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1961_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n446), .CK(clk), 
        .Q(cell_1961_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1961_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1961_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1961_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1962_U4 ( .A(signal_3528), .B(cell_1962_and_out[1]), .Z(
        signal_3740) );
  XOR2_X1 cell_1962_U3 ( .A(signal_2090), .B(cell_1962_and_out[0]), .Z(
        signal_2230) );
  XOR2_X1 cell_1962_U2 ( .A(signal_3528), .B(signal_3485), .Z(
        cell_1962_and_in[1]) );
  XOR2_X1 cell_1962_U1 ( .A(signal_2090), .B(signal_2047), .Z(
        cell_1962_and_in[0]) );
  XOR2_X1 cell_1962_a_HPC2_and_U14 ( .A(Fresh[248]), .B(cell_1962_and_in[0]), 
        .Z(cell_1962_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1962_a_HPC2_and_U13 ( .A(Fresh[248]), .B(cell_1962_and_in[1]), 
        .Z(cell_1962_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1962_a_HPC2_and_U12 ( .A1(cell_1962_a_HPC2_and_a_reg[1]), .A2(
        cell_1962_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1962_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1962_a_HPC2_and_U11 ( .A1(cell_1962_a_HPC2_and_a_reg[0]), .A2(
        cell_1962_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1962_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1962_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1962_a_HPC2_and_n9), 
        .ZN(cell_1962_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1962_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1962_a_HPC2_and_n9), 
        .ZN(cell_1962_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1962_a_HPC2_and_U8 ( .A(Fresh[248]), .ZN(cell_1962_a_HPC2_and_n9) );
  AND2_X1 cell_1962_a_HPC2_and_U7 ( .A1(cell_1962_and_in[1]), .A2(n447), .ZN(
        cell_1962_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1962_a_HPC2_and_U6 ( .A1(cell_1962_and_in[0]), .A2(n433), .ZN(
        cell_1962_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1962_a_HPC2_and_U5 ( .A(cell_1962_a_HPC2_and_n8), .B(
        cell_1962_a_HPC2_and_z_1__1_), .ZN(cell_1962_and_out[1]) );
  XNOR2_X1 cell_1962_a_HPC2_and_U4 ( .A(
        cell_1962_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1962_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1962_a_HPC2_and_n8) );
  XNOR2_X1 cell_1962_a_HPC2_and_U3 ( .A(cell_1962_a_HPC2_and_n7), .B(
        cell_1962_a_HPC2_and_z_0__0_), .ZN(cell_1962_and_out[0]) );
  XNOR2_X1 cell_1962_a_HPC2_and_U2 ( .A(
        cell_1962_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1962_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1962_a_HPC2_and_n7) );
  DFF_X1 cell_1962_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1962_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1962_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1962_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1962_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1962_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1962_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1962_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1962_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1962_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1963_U4 ( .A(signal_3510), .B(cell_1963_and_out[1]), .Z(
        signal_3741) );
  XOR2_X1 cell_1963_U3 ( .A(signal_2072), .B(cell_1963_and_out[0]), .Z(
        signal_2231) );
  XOR2_X1 cell_1963_U2 ( .A(signal_3510), .B(signal_3493), .Z(
        cell_1963_and_in[1]) );
  XOR2_X1 cell_1963_U1 ( .A(signal_2072), .B(signal_2055), .Z(
        cell_1963_and_in[0]) );
  XOR2_X1 cell_1963_a_HPC2_and_U14 ( .A(Fresh[249]), .B(cell_1963_and_in[0]), 
        .Z(cell_1963_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1963_a_HPC2_and_U13 ( .A(Fresh[249]), .B(cell_1963_and_in[1]), 
        .Z(cell_1963_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1963_a_HPC2_and_U12 ( .A1(cell_1963_a_HPC2_and_a_reg[1]), .A2(
        cell_1963_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1963_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1963_a_HPC2_and_U11 ( .A1(cell_1963_a_HPC2_and_a_reg[0]), .A2(
        cell_1963_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1963_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1963_a_HPC2_and_U10 ( .A1(n452), .A2(cell_1963_a_HPC2_and_n9), 
        .ZN(cell_1963_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1963_a_HPC2_and_U9 ( .A1(n438), .A2(cell_1963_a_HPC2_and_n9), 
        .ZN(cell_1963_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1963_a_HPC2_and_U8 ( .A(Fresh[249]), .ZN(cell_1963_a_HPC2_and_n9) );
  AND2_X1 cell_1963_a_HPC2_and_U7 ( .A1(cell_1963_and_in[1]), .A2(n452), .ZN(
        cell_1963_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1963_a_HPC2_and_U6 ( .A1(cell_1963_and_in[0]), .A2(n438), .ZN(
        cell_1963_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1963_a_HPC2_and_U5 ( .A(cell_1963_a_HPC2_and_n8), .B(
        cell_1963_a_HPC2_and_z_1__1_), .ZN(cell_1963_and_out[1]) );
  XNOR2_X1 cell_1963_a_HPC2_and_U4 ( .A(
        cell_1963_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1963_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1963_a_HPC2_and_n8) );
  XNOR2_X1 cell_1963_a_HPC2_and_U3 ( .A(cell_1963_a_HPC2_and_n7), .B(
        cell_1963_a_HPC2_and_z_0__0_), .ZN(cell_1963_and_out[0]) );
  XNOR2_X1 cell_1963_a_HPC2_and_U2 ( .A(
        cell_1963_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1963_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1963_a_HPC2_and_n7) );
  DFF_X1 cell_1963_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1963_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1963_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n438), .CK(clk), 
        .Q(cell_1963_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1963_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1963_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n452), .CK(clk), 
        .Q(cell_1963_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1963_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1963_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1963_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1964_U4 ( .A(signal_3566), .B(cell_1964_and_out[1]), .Z(
        signal_3742) );
  XOR2_X1 cell_1964_U3 ( .A(signal_2128), .B(cell_1964_and_out[0]), .Z(
        signal_2232) );
  XOR2_X1 cell_1964_U2 ( .A(signal_3566), .B(signal_3484), .Z(
        cell_1964_and_in[1]) );
  XOR2_X1 cell_1964_U1 ( .A(signal_2128), .B(signal_2046), .Z(
        cell_1964_and_in[0]) );
  XOR2_X1 cell_1964_a_HPC2_and_U14 ( .A(Fresh[250]), .B(cell_1964_and_in[0]), 
        .Z(cell_1964_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1964_a_HPC2_and_U13 ( .A(Fresh[250]), .B(cell_1964_and_in[1]), 
        .Z(cell_1964_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1964_a_HPC2_and_U12 ( .A1(cell_1964_a_HPC2_and_a_reg[1]), .A2(
        cell_1964_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1964_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1964_a_HPC2_and_U11 ( .A1(cell_1964_a_HPC2_and_a_reg[0]), .A2(
        cell_1964_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1964_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1964_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1964_a_HPC2_and_n9), 
        .ZN(cell_1964_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1964_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1964_a_HPC2_and_n9), 
        .ZN(cell_1964_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1964_a_HPC2_and_U8 ( .A(Fresh[250]), .ZN(cell_1964_a_HPC2_and_n9) );
  AND2_X1 cell_1964_a_HPC2_and_U7 ( .A1(cell_1964_and_in[1]), .A2(n447), .ZN(
        cell_1964_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1964_a_HPC2_and_U6 ( .A1(cell_1964_and_in[0]), .A2(n433), .ZN(
        cell_1964_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1964_a_HPC2_and_U5 ( .A(cell_1964_a_HPC2_and_n8), .B(
        cell_1964_a_HPC2_and_z_1__1_), .ZN(cell_1964_and_out[1]) );
  XNOR2_X1 cell_1964_a_HPC2_and_U4 ( .A(
        cell_1964_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1964_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1964_a_HPC2_and_n8) );
  XNOR2_X1 cell_1964_a_HPC2_and_U3 ( .A(cell_1964_a_HPC2_and_n7), .B(
        cell_1964_a_HPC2_and_z_0__0_), .ZN(cell_1964_and_out[0]) );
  XNOR2_X1 cell_1964_a_HPC2_and_U2 ( .A(
        cell_1964_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1964_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1964_a_HPC2_and_n7) );
  DFF_X1 cell_1964_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1964_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1964_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1964_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1964_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1964_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1964_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1964_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1964_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1964_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1965_U4 ( .A(signal_3585), .B(cell_1965_and_out[1]), .Z(
        signal_3743) );
  XOR2_X1 cell_1965_U3 ( .A(signal_2147), .B(cell_1965_and_out[0]), .Z(
        signal_2233) );
  XOR2_X1 cell_1965_U2 ( .A(signal_3585), .B(signal_3527), .Z(
        cell_1965_and_in[1]) );
  XOR2_X1 cell_1965_U1 ( .A(signal_2147), .B(signal_2089), .Z(
        cell_1965_and_in[0]) );
  XOR2_X1 cell_1965_a_HPC2_and_U14 ( .A(Fresh[251]), .B(cell_1965_and_in[0]), 
        .Z(cell_1965_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1965_a_HPC2_and_U13 ( .A(Fresh[251]), .B(cell_1965_and_in[1]), 
        .Z(cell_1965_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1965_a_HPC2_and_U12 ( .A1(cell_1965_a_HPC2_and_a_reg[1]), .A2(
        cell_1965_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1965_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1965_a_HPC2_and_U11 ( .A1(cell_1965_a_HPC2_and_a_reg[0]), .A2(
        cell_1965_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1965_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1965_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1965_a_HPC2_and_n9), 
        .ZN(cell_1965_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1965_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1965_a_HPC2_and_n9), 
        .ZN(cell_1965_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1965_a_HPC2_and_U8 ( .A(Fresh[251]), .ZN(cell_1965_a_HPC2_and_n9) );
  AND2_X1 cell_1965_a_HPC2_and_U7 ( .A1(cell_1965_and_in[1]), .A2(n447), .ZN(
        cell_1965_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1965_a_HPC2_and_U6 ( .A1(cell_1965_and_in[0]), .A2(n433), .ZN(
        cell_1965_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1965_a_HPC2_and_U5 ( .A(cell_1965_a_HPC2_and_n8), .B(
        cell_1965_a_HPC2_and_z_1__1_), .ZN(cell_1965_and_out[1]) );
  XNOR2_X1 cell_1965_a_HPC2_and_U4 ( .A(
        cell_1965_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1965_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1965_a_HPC2_and_n8) );
  XNOR2_X1 cell_1965_a_HPC2_and_U3 ( .A(cell_1965_a_HPC2_and_n7), .B(
        cell_1965_a_HPC2_and_z_0__0_), .ZN(cell_1965_and_out[0]) );
  XNOR2_X1 cell_1965_a_HPC2_and_U2 ( .A(
        cell_1965_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1965_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1965_a_HPC2_and_n7) );
  DFF_X1 cell_1965_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1965_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1965_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1965_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1965_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1965_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1965_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1965_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1965_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1965_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1966_U4 ( .A(signal_3524), .B(cell_1966_and_out[1]), .Z(
        signal_3744) );
  XOR2_X1 cell_1966_U3 ( .A(signal_2086), .B(cell_1966_and_out[0]), .Z(
        signal_2234) );
  XOR2_X1 cell_1966_U2 ( .A(signal_3524), .B(signal_3431), .Z(
        cell_1966_and_in[1]) );
  XOR2_X1 cell_1966_U1 ( .A(signal_2086), .B(signal_2017), .Z(
        cell_1966_and_in[0]) );
  XOR2_X1 cell_1966_a_HPC2_and_U14 ( .A(Fresh[252]), .B(cell_1966_and_in[0]), 
        .Z(cell_1966_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1966_a_HPC2_and_U13 ( .A(Fresh[252]), .B(cell_1966_and_in[1]), 
        .Z(cell_1966_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1966_a_HPC2_and_U12 ( .A1(cell_1966_a_HPC2_and_a_reg[1]), .A2(
        cell_1966_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1966_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1966_a_HPC2_and_U11 ( .A1(cell_1966_a_HPC2_and_a_reg[0]), .A2(
        cell_1966_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1966_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1966_a_HPC2_and_U10 ( .A1(n451), .A2(cell_1966_a_HPC2_and_n9), 
        .ZN(cell_1966_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1966_a_HPC2_and_U9 ( .A1(n437), .A2(cell_1966_a_HPC2_and_n9), 
        .ZN(cell_1966_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1966_a_HPC2_and_U8 ( .A(Fresh[252]), .ZN(cell_1966_a_HPC2_and_n9) );
  AND2_X1 cell_1966_a_HPC2_and_U7 ( .A1(cell_1966_and_in[1]), .A2(n451), .ZN(
        cell_1966_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1966_a_HPC2_and_U6 ( .A1(cell_1966_and_in[0]), .A2(n437), .ZN(
        cell_1966_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1966_a_HPC2_and_U5 ( .A(cell_1966_a_HPC2_and_n8), .B(
        cell_1966_a_HPC2_and_z_1__1_), .ZN(cell_1966_and_out[1]) );
  XNOR2_X1 cell_1966_a_HPC2_and_U4 ( .A(
        cell_1966_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1966_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1966_a_HPC2_and_n8) );
  XNOR2_X1 cell_1966_a_HPC2_and_U3 ( .A(cell_1966_a_HPC2_and_n7), .B(
        cell_1966_a_HPC2_and_z_0__0_), .ZN(cell_1966_and_out[0]) );
  XNOR2_X1 cell_1966_a_HPC2_and_U2 ( .A(
        cell_1966_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1966_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1966_a_HPC2_and_n7) );
  DFF_X1 cell_1966_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1966_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1966_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n437), .CK(clk), 
        .Q(cell_1966_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1966_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1966_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n451), .CK(clk), 
        .Q(cell_1966_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1966_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1966_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1966_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1967_U4 ( .A(signal_3460), .B(cell_1967_and_out[1]), .Z(
        signal_3745) );
  XOR2_X1 cell_1967_U3 ( .A(signal_2022), .B(cell_1967_and_out[0]), .Z(
        signal_2235) );
  XOR2_X1 cell_1967_U2 ( .A(signal_3460), .B(signal_3550), .Z(
        cell_1967_and_in[1]) );
  XOR2_X1 cell_1967_U1 ( .A(signal_2022), .B(signal_2112), .Z(
        cell_1967_and_in[0]) );
  XOR2_X1 cell_1967_a_HPC2_and_U14 ( .A(Fresh[253]), .B(cell_1967_and_in[0]), 
        .Z(cell_1967_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1967_a_HPC2_and_U13 ( .A(Fresh[253]), .B(cell_1967_and_in[1]), 
        .Z(cell_1967_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1967_a_HPC2_and_U12 ( .A1(cell_1967_a_HPC2_and_a_reg[1]), .A2(
        cell_1967_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1967_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1967_a_HPC2_and_U11 ( .A1(cell_1967_a_HPC2_and_a_reg[0]), .A2(
        cell_1967_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1967_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1967_a_HPC2_and_U10 ( .A1(n450), .A2(cell_1967_a_HPC2_and_n9), 
        .ZN(cell_1967_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1967_a_HPC2_and_U9 ( .A1(n436), .A2(cell_1967_a_HPC2_and_n9), 
        .ZN(cell_1967_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1967_a_HPC2_and_U8 ( .A(Fresh[253]), .ZN(cell_1967_a_HPC2_and_n9) );
  AND2_X1 cell_1967_a_HPC2_and_U7 ( .A1(cell_1967_and_in[1]), .A2(n450), .ZN(
        cell_1967_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1967_a_HPC2_and_U6 ( .A1(cell_1967_and_in[0]), .A2(n436), .ZN(
        cell_1967_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1967_a_HPC2_and_U5 ( .A(cell_1967_a_HPC2_and_n8), .B(
        cell_1967_a_HPC2_and_z_1__1_), .ZN(cell_1967_and_out[1]) );
  XNOR2_X1 cell_1967_a_HPC2_and_U4 ( .A(
        cell_1967_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1967_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1967_a_HPC2_and_n8) );
  XNOR2_X1 cell_1967_a_HPC2_and_U3 ( .A(cell_1967_a_HPC2_and_n7), .B(
        cell_1967_a_HPC2_and_z_0__0_), .ZN(cell_1967_and_out[0]) );
  XNOR2_X1 cell_1967_a_HPC2_and_U2 ( .A(
        cell_1967_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1967_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1967_a_HPC2_and_n7) );
  DFF_X1 cell_1967_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1967_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1967_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_1967_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1967_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1967_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_1967_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1967_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1967_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1967_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1968_U4 ( .A(signal_3484), .B(cell_1968_and_out[1]), .Z(
        signal_3746) );
  XOR2_X1 cell_1968_U3 ( .A(signal_2046), .B(cell_1968_and_out[0]), .Z(
        signal_2236) );
  XOR2_X1 cell_1968_U2 ( .A(signal_3484), .B(signal_3544), .Z(
        cell_1968_and_in[1]) );
  XOR2_X1 cell_1968_U1 ( .A(signal_2046), .B(signal_2106), .Z(
        cell_1968_and_in[0]) );
  XOR2_X1 cell_1968_a_HPC2_and_U14 ( .A(Fresh[254]), .B(cell_1968_and_in[0]), 
        .Z(cell_1968_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1968_a_HPC2_and_U13 ( .A(Fresh[254]), .B(cell_1968_and_in[1]), 
        .Z(cell_1968_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1968_a_HPC2_and_U12 ( .A1(cell_1968_a_HPC2_and_a_reg[1]), .A2(
        cell_1968_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1968_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1968_a_HPC2_and_U11 ( .A1(cell_1968_a_HPC2_and_a_reg[0]), .A2(
        cell_1968_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1968_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1968_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1968_a_HPC2_and_n9), 
        .ZN(cell_1968_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1968_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1968_a_HPC2_and_n9), 
        .ZN(cell_1968_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1968_a_HPC2_and_U8 ( .A(Fresh[254]), .ZN(cell_1968_a_HPC2_and_n9) );
  AND2_X1 cell_1968_a_HPC2_and_U7 ( .A1(cell_1968_and_in[1]), .A2(n447), .ZN(
        cell_1968_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1968_a_HPC2_and_U6 ( .A1(cell_1968_and_in[0]), .A2(n433), .ZN(
        cell_1968_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1968_a_HPC2_and_U5 ( .A(cell_1968_a_HPC2_and_n8), .B(
        cell_1968_a_HPC2_and_z_1__1_), .ZN(cell_1968_and_out[1]) );
  XNOR2_X1 cell_1968_a_HPC2_and_U4 ( .A(
        cell_1968_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1968_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1968_a_HPC2_and_n8) );
  XNOR2_X1 cell_1968_a_HPC2_and_U3 ( .A(cell_1968_a_HPC2_and_n7), .B(
        cell_1968_a_HPC2_and_z_0__0_), .ZN(cell_1968_and_out[0]) );
  XNOR2_X1 cell_1968_a_HPC2_and_U2 ( .A(
        cell_1968_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1968_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1968_a_HPC2_and_n7) );
  DFF_X1 cell_1968_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1968_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1968_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1968_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1968_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1968_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1968_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1968_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1968_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1968_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1969_U4 ( .A(signal_3587), .B(cell_1969_and_out[1]), .Z(
        signal_3747) );
  XOR2_X1 cell_1969_U3 ( .A(signal_2149), .B(cell_1969_and_out[0]), .Z(
        signal_2237) );
  XOR2_X1 cell_1969_U2 ( .A(signal_3587), .B(signal_3487), .Z(
        cell_1969_and_in[1]) );
  XOR2_X1 cell_1969_U1 ( .A(signal_2149), .B(signal_2049), .Z(
        cell_1969_and_in[0]) );
  XOR2_X1 cell_1969_a_HPC2_and_U14 ( .A(Fresh[255]), .B(cell_1969_and_in[0]), 
        .Z(cell_1969_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1969_a_HPC2_and_U13 ( .A(Fresh[255]), .B(cell_1969_and_in[1]), 
        .Z(cell_1969_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1969_a_HPC2_and_U12 ( .A1(cell_1969_a_HPC2_and_a_reg[1]), .A2(
        cell_1969_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1969_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1969_a_HPC2_and_U11 ( .A1(cell_1969_a_HPC2_and_a_reg[0]), .A2(
        cell_1969_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1969_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1969_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1969_a_HPC2_and_n9), 
        .ZN(cell_1969_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1969_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1969_a_HPC2_and_n9), 
        .ZN(cell_1969_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1969_a_HPC2_and_U8 ( .A(Fresh[255]), .ZN(cell_1969_a_HPC2_and_n9) );
  AND2_X1 cell_1969_a_HPC2_and_U7 ( .A1(cell_1969_and_in[1]), .A2(n454), .ZN(
        cell_1969_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1969_a_HPC2_and_U6 ( .A1(cell_1969_and_in[0]), .A2(n440), .ZN(
        cell_1969_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1969_a_HPC2_and_U5 ( .A(cell_1969_a_HPC2_and_n8), .B(
        cell_1969_a_HPC2_and_z_1__1_), .ZN(cell_1969_and_out[1]) );
  XNOR2_X1 cell_1969_a_HPC2_and_U4 ( .A(
        cell_1969_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1969_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1969_a_HPC2_and_n8) );
  XNOR2_X1 cell_1969_a_HPC2_and_U3 ( .A(cell_1969_a_HPC2_and_n7), .B(
        cell_1969_a_HPC2_and_z_0__0_), .ZN(cell_1969_and_out[0]) );
  XNOR2_X1 cell_1969_a_HPC2_and_U2 ( .A(
        cell_1969_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1969_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1969_a_HPC2_and_n7) );
  DFF_X1 cell_1969_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1969_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1969_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1969_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1969_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1969_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1969_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1969_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1969_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1969_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1970_U4 ( .A(signal_3422), .B(cell_1970_and_out[1]), .Z(
        signal_3748) );
  XOR2_X1 cell_1970_U3 ( .A(signal_2008), .B(cell_1970_and_out[0]), .Z(
        signal_2238) );
  XOR2_X1 cell_1970_U2 ( .A(signal_3422), .B(signal_3463), .Z(
        cell_1970_and_in[1]) );
  XOR2_X1 cell_1970_U1 ( .A(signal_2008), .B(signal_2025), .Z(
        cell_1970_and_in[0]) );
  XOR2_X1 cell_1970_a_HPC2_and_U14 ( .A(Fresh[256]), .B(cell_1970_and_in[0]), 
        .Z(cell_1970_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1970_a_HPC2_and_U13 ( .A(Fresh[256]), .B(cell_1970_and_in[1]), 
        .Z(cell_1970_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1970_a_HPC2_and_U12 ( .A1(cell_1970_a_HPC2_and_a_reg[1]), .A2(
        cell_1970_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1970_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1970_a_HPC2_and_U11 ( .A1(cell_1970_a_HPC2_and_a_reg[0]), .A2(
        cell_1970_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1970_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1970_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1970_a_HPC2_and_n9), 
        .ZN(cell_1970_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1970_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1970_a_HPC2_and_n9), 
        .ZN(cell_1970_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1970_a_HPC2_and_U8 ( .A(Fresh[256]), .ZN(cell_1970_a_HPC2_and_n9) );
  AND2_X1 cell_1970_a_HPC2_and_U7 ( .A1(cell_1970_and_in[1]), .A2(n447), .ZN(
        cell_1970_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1970_a_HPC2_and_U6 ( .A1(cell_1970_and_in[0]), .A2(n433), .ZN(
        cell_1970_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1970_a_HPC2_and_U5 ( .A(cell_1970_a_HPC2_and_n8), .B(
        cell_1970_a_HPC2_and_z_1__1_), .ZN(cell_1970_and_out[1]) );
  XNOR2_X1 cell_1970_a_HPC2_and_U4 ( .A(
        cell_1970_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1970_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1970_a_HPC2_and_n8) );
  XNOR2_X1 cell_1970_a_HPC2_and_U3 ( .A(cell_1970_a_HPC2_and_n7), .B(
        cell_1970_a_HPC2_and_z_0__0_), .ZN(cell_1970_and_out[0]) );
  XNOR2_X1 cell_1970_a_HPC2_and_U2 ( .A(
        cell_1970_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1970_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1970_a_HPC2_and_n7) );
  DFF_X1 cell_1970_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1970_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1970_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1970_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1970_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1970_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1970_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1970_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1970_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1970_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1971_U4 ( .A(signal_3505), .B(cell_1971_and_out[1]), .Z(
        signal_3749) );
  XOR2_X1 cell_1971_U3 ( .A(signal_2067), .B(cell_1971_and_out[0]), .Z(
        signal_2239) );
  XOR2_X1 cell_1971_U2 ( .A(signal_3505), .B(signal_3561), .Z(
        cell_1971_and_in[1]) );
  XOR2_X1 cell_1971_U1 ( .A(signal_2067), .B(signal_2123), .Z(
        cell_1971_and_in[0]) );
  XOR2_X1 cell_1971_a_HPC2_and_U14 ( .A(Fresh[257]), .B(cell_1971_and_in[0]), 
        .Z(cell_1971_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1971_a_HPC2_and_U13 ( .A(Fresh[257]), .B(cell_1971_and_in[1]), 
        .Z(cell_1971_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1971_a_HPC2_and_U12 ( .A1(cell_1971_a_HPC2_and_a_reg[1]), .A2(
        cell_1971_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1971_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1971_a_HPC2_and_U11 ( .A1(cell_1971_a_HPC2_and_a_reg[0]), .A2(
        cell_1971_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1971_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1971_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1971_a_HPC2_and_n9), 
        .ZN(cell_1971_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1971_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1971_a_HPC2_and_n9), 
        .ZN(cell_1971_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1971_a_HPC2_and_U8 ( .A(Fresh[257]), .ZN(cell_1971_a_HPC2_and_n9) );
  AND2_X1 cell_1971_a_HPC2_and_U7 ( .A1(cell_1971_and_in[1]), .A2(n454), .ZN(
        cell_1971_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1971_a_HPC2_and_U6 ( .A1(cell_1971_and_in[0]), .A2(n440), .ZN(
        cell_1971_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1971_a_HPC2_and_U5 ( .A(cell_1971_a_HPC2_and_n8), .B(
        cell_1971_a_HPC2_and_z_1__1_), .ZN(cell_1971_and_out[1]) );
  XNOR2_X1 cell_1971_a_HPC2_and_U4 ( .A(
        cell_1971_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1971_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1971_a_HPC2_and_n8) );
  XNOR2_X1 cell_1971_a_HPC2_and_U3 ( .A(cell_1971_a_HPC2_and_n7), .B(
        cell_1971_a_HPC2_and_z_0__0_), .ZN(cell_1971_and_out[0]) );
  XNOR2_X1 cell_1971_a_HPC2_and_U2 ( .A(
        cell_1971_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1971_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1971_a_HPC2_and_n7) );
  DFF_X1 cell_1971_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1971_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1971_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1971_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1971_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1971_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1971_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1971_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1971_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1971_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1972_U4 ( .A(signal_3527), .B(cell_1972_and_out[1]), .Z(
        signal_3750) );
  XOR2_X1 cell_1972_U3 ( .A(signal_2089), .B(cell_1972_and_out[0]), .Z(
        signal_2240) );
  XOR2_X1 cell_1972_U2 ( .A(signal_3527), .B(signal_3478), .Z(
        cell_1972_and_in[1]) );
  XOR2_X1 cell_1972_U1 ( .A(signal_2089), .B(signal_2040), .Z(
        cell_1972_and_in[0]) );
  XOR2_X1 cell_1972_a_HPC2_and_U14 ( .A(Fresh[258]), .B(cell_1972_and_in[0]), 
        .Z(cell_1972_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1972_a_HPC2_and_U13 ( .A(Fresh[258]), .B(cell_1972_and_in[1]), 
        .Z(cell_1972_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1972_a_HPC2_and_U12 ( .A1(cell_1972_a_HPC2_and_a_reg[1]), .A2(
        cell_1972_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1972_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1972_a_HPC2_and_U11 ( .A1(cell_1972_a_HPC2_and_a_reg[0]), .A2(
        cell_1972_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1972_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1972_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1972_a_HPC2_and_n9), 
        .ZN(cell_1972_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1972_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1972_a_HPC2_and_n9), 
        .ZN(cell_1972_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1972_a_HPC2_and_U8 ( .A(Fresh[258]), .ZN(cell_1972_a_HPC2_and_n9) );
  AND2_X1 cell_1972_a_HPC2_and_U7 ( .A1(cell_1972_and_in[1]), .A2(n447), .ZN(
        cell_1972_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1972_a_HPC2_and_U6 ( .A1(cell_1972_and_in[0]), .A2(n433), .ZN(
        cell_1972_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1972_a_HPC2_and_U5 ( .A(cell_1972_a_HPC2_and_n8), .B(
        cell_1972_a_HPC2_and_z_1__1_), .ZN(cell_1972_and_out[1]) );
  XNOR2_X1 cell_1972_a_HPC2_and_U4 ( .A(
        cell_1972_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1972_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1972_a_HPC2_and_n8) );
  XNOR2_X1 cell_1972_a_HPC2_and_U3 ( .A(cell_1972_a_HPC2_and_n7), .B(
        cell_1972_a_HPC2_and_z_0__0_), .ZN(cell_1972_and_out[0]) );
  XNOR2_X1 cell_1972_a_HPC2_and_U2 ( .A(
        cell_1972_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1972_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1972_a_HPC2_and_n7) );
  DFF_X1 cell_1972_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1972_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1972_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1972_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1972_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1972_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1972_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1972_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1972_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1972_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1973_U4 ( .A(signal_3530), .B(cell_1973_and_out[1]), .Z(
        signal_3751) );
  XOR2_X1 cell_1973_U3 ( .A(signal_2092), .B(cell_1973_and_out[0]), .Z(
        signal_2241) );
  XOR2_X1 cell_1973_U2 ( .A(signal_3530), .B(signal_3509), .Z(
        cell_1973_and_in[1]) );
  XOR2_X1 cell_1973_U1 ( .A(signal_2092), .B(signal_2071), .Z(
        cell_1973_and_in[0]) );
  XOR2_X1 cell_1973_a_HPC2_and_U14 ( .A(Fresh[259]), .B(cell_1973_and_in[0]), 
        .Z(cell_1973_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1973_a_HPC2_and_U13 ( .A(Fresh[259]), .B(cell_1973_and_in[1]), 
        .Z(cell_1973_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1973_a_HPC2_and_U12 ( .A1(cell_1973_a_HPC2_and_a_reg[1]), .A2(
        cell_1973_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1973_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1973_a_HPC2_and_U11 ( .A1(cell_1973_a_HPC2_and_a_reg[0]), .A2(
        cell_1973_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1973_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1973_a_HPC2_and_U10 ( .A1(n447), .A2(cell_1973_a_HPC2_and_n9), 
        .ZN(cell_1973_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1973_a_HPC2_and_U9 ( .A1(n433), .A2(cell_1973_a_HPC2_and_n9), 
        .ZN(cell_1973_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1973_a_HPC2_and_U8 ( .A(Fresh[259]), .ZN(cell_1973_a_HPC2_and_n9) );
  AND2_X1 cell_1973_a_HPC2_and_U7 ( .A1(cell_1973_and_in[1]), .A2(n447), .ZN(
        cell_1973_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1973_a_HPC2_and_U6 ( .A1(cell_1973_and_in[0]), .A2(n433), .ZN(
        cell_1973_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1973_a_HPC2_and_U5 ( .A(cell_1973_a_HPC2_and_n8), .B(
        cell_1973_a_HPC2_and_z_1__1_), .ZN(cell_1973_and_out[1]) );
  XNOR2_X1 cell_1973_a_HPC2_and_U4 ( .A(
        cell_1973_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1973_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1973_a_HPC2_and_n8) );
  XNOR2_X1 cell_1973_a_HPC2_and_U3 ( .A(cell_1973_a_HPC2_and_n7), .B(
        cell_1973_a_HPC2_and_z_0__0_), .ZN(cell_1973_and_out[0]) );
  XNOR2_X1 cell_1973_a_HPC2_and_U2 ( .A(
        cell_1973_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1973_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1973_a_HPC2_and_n7) );
  DFF_X1 cell_1973_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1973_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1973_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n433), .CK(clk), 
        .Q(cell_1973_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1973_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1973_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n447), .CK(clk), 
        .Q(cell_1973_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1973_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1973_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1973_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1974_U4 ( .A(signal_3532), .B(cell_1974_and_out[1]), .Z(
        signal_3752) );
  XOR2_X1 cell_1974_U3 ( .A(signal_2094), .B(cell_1974_and_out[0]), .Z(
        signal_2242) );
  XOR2_X1 cell_1974_U2 ( .A(signal_3532), .B(signal_3572), .Z(
        cell_1974_and_in[1]) );
  XOR2_X1 cell_1974_U1 ( .A(signal_2094), .B(signal_2134), .Z(
        cell_1974_and_in[0]) );
  XOR2_X1 cell_1974_a_HPC2_and_U14 ( .A(Fresh[260]), .B(cell_1974_and_in[0]), 
        .Z(cell_1974_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1974_a_HPC2_and_U13 ( .A(Fresh[260]), .B(cell_1974_and_in[1]), 
        .Z(cell_1974_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1974_a_HPC2_and_U12 ( .A1(cell_1974_a_HPC2_and_a_reg[1]), .A2(
        cell_1974_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1974_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1974_a_HPC2_and_U11 ( .A1(cell_1974_a_HPC2_and_a_reg[0]), .A2(
        cell_1974_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1974_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1974_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1974_a_HPC2_and_n9), 
        .ZN(cell_1974_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1974_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1974_a_HPC2_and_n9), 
        .ZN(cell_1974_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1974_a_HPC2_and_U8 ( .A(Fresh[260]), .ZN(cell_1974_a_HPC2_and_n9) );
  AND2_X1 cell_1974_a_HPC2_and_U7 ( .A1(cell_1974_and_in[1]), .A2(n454), .ZN(
        cell_1974_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1974_a_HPC2_and_U6 ( .A1(cell_1974_and_in[0]), .A2(n440), .ZN(
        cell_1974_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1974_a_HPC2_and_U5 ( .A(cell_1974_a_HPC2_and_n8), .B(
        cell_1974_a_HPC2_and_z_1__1_), .ZN(cell_1974_and_out[1]) );
  XNOR2_X1 cell_1974_a_HPC2_and_U4 ( .A(
        cell_1974_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1974_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1974_a_HPC2_and_n8) );
  XNOR2_X1 cell_1974_a_HPC2_and_U3 ( .A(cell_1974_a_HPC2_and_n7), .B(
        cell_1974_a_HPC2_and_z_0__0_), .ZN(cell_1974_and_out[0]) );
  XNOR2_X1 cell_1974_a_HPC2_and_U2 ( .A(
        cell_1974_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1974_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1974_a_HPC2_and_n7) );
  DFF_X1 cell_1974_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1974_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1974_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1974_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1974_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1974_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1974_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1974_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1974_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1974_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1975_U4 ( .A(signal_3428), .B(cell_1975_and_out[1]), .Z(
        signal_3753) );
  XOR2_X1 cell_1975_U3 ( .A(signal_2014), .B(cell_1975_and_out[0]), .Z(
        signal_2243) );
  XOR2_X1 cell_1975_U2 ( .A(signal_3428), .B(signal_3581), .Z(
        cell_1975_and_in[1]) );
  XOR2_X1 cell_1975_U1 ( .A(signal_2014), .B(signal_2143), .Z(
        cell_1975_and_in[0]) );
  XOR2_X1 cell_1975_a_HPC2_and_U14 ( .A(Fresh[261]), .B(cell_1975_and_in[0]), 
        .Z(cell_1975_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1975_a_HPC2_and_U13 ( .A(Fresh[261]), .B(cell_1975_and_in[1]), 
        .Z(cell_1975_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1975_a_HPC2_and_U12 ( .A1(cell_1975_a_HPC2_and_a_reg[1]), .A2(
        cell_1975_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1975_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1975_a_HPC2_and_U11 ( .A1(cell_1975_a_HPC2_and_a_reg[0]), .A2(
        cell_1975_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1975_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1975_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1975_a_HPC2_and_n9), 
        .ZN(cell_1975_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1975_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1975_a_HPC2_and_n9), 
        .ZN(cell_1975_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1975_a_HPC2_and_U8 ( .A(Fresh[261]), .ZN(cell_1975_a_HPC2_and_n9) );
  AND2_X1 cell_1975_a_HPC2_and_U7 ( .A1(cell_1975_and_in[1]), .A2(n454), .ZN(
        cell_1975_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1975_a_HPC2_and_U6 ( .A1(cell_1975_and_in[0]), .A2(n440), .ZN(
        cell_1975_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1975_a_HPC2_and_U5 ( .A(cell_1975_a_HPC2_and_n8), .B(
        cell_1975_a_HPC2_and_z_1__1_), .ZN(cell_1975_and_out[1]) );
  XNOR2_X1 cell_1975_a_HPC2_and_U4 ( .A(
        cell_1975_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1975_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1975_a_HPC2_and_n8) );
  XNOR2_X1 cell_1975_a_HPC2_and_U3 ( .A(cell_1975_a_HPC2_and_n7), .B(
        cell_1975_a_HPC2_and_z_0__0_), .ZN(cell_1975_and_out[0]) );
  XNOR2_X1 cell_1975_a_HPC2_and_U2 ( .A(
        cell_1975_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1975_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1975_a_HPC2_and_n7) );
  DFF_X1 cell_1975_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1975_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1975_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1975_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1975_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1975_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1975_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1975_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1975_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1975_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1976_U4 ( .A(signal_3522), .B(cell_1976_and_out[1]), .Z(
        signal_3754) );
  XOR2_X1 cell_1976_U3 ( .A(signal_2084), .B(cell_1976_and_out[0]), .Z(
        signal_2244) );
  XOR2_X1 cell_1976_U2 ( .A(signal_3522), .B(n367), .Z(cell_1976_and_in[1]) );
  XOR2_X1 cell_1976_U1 ( .A(signal_2084), .B(n366), .Z(cell_1976_and_in[0]) );
  XOR2_X1 cell_1976_a_HPC2_and_U14 ( .A(Fresh[262]), .B(cell_1976_and_in[0]), 
        .Z(cell_1976_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1976_a_HPC2_and_U13 ( .A(Fresh[262]), .B(cell_1976_and_in[1]), 
        .Z(cell_1976_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1976_a_HPC2_and_U12 ( .A1(cell_1976_a_HPC2_and_a_reg[1]), .A2(
        cell_1976_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1976_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1976_a_HPC2_and_U11 ( .A1(cell_1976_a_HPC2_and_a_reg[0]), .A2(
        cell_1976_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1976_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1976_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1976_a_HPC2_and_n9), 
        .ZN(cell_1976_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1976_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1976_a_HPC2_and_n9), 
        .ZN(cell_1976_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1976_a_HPC2_and_U8 ( .A(Fresh[262]), .ZN(cell_1976_a_HPC2_and_n9) );
  AND2_X1 cell_1976_a_HPC2_and_U7 ( .A1(cell_1976_and_in[1]), .A2(n448), .ZN(
        cell_1976_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1976_a_HPC2_and_U6 ( .A1(cell_1976_and_in[0]), .A2(n434), .ZN(
        cell_1976_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1976_a_HPC2_and_U5 ( .A(cell_1976_a_HPC2_and_n8), .B(
        cell_1976_a_HPC2_and_z_1__1_), .ZN(cell_1976_and_out[1]) );
  XNOR2_X1 cell_1976_a_HPC2_and_U4 ( .A(
        cell_1976_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1976_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1976_a_HPC2_and_n8) );
  XNOR2_X1 cell_1976_a_HPC2_and_U3 ( .A(cell_1976_a_HPC2_and_n7), .B(
        cell_1976_a_HPC2_and_z_0__0_), .ZN(cell_1976_and_out[0]) );
  XNOR2_X1 cell_1976_a_HPC2_and_U2 ( .A(
        cell_1976_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1976_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1976_a_HPC2_and_n7) );
  DFF_X1 cell_1976_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1976_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1976_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1976_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1976_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1976_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1976_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1976_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1976_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1976_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1977_U4 ( .A(signal_3421), .B(cell_1977_and_out[1]), .Z(
        signal_3755) );
  XOR2_X1 cell_1977_U3 ( .A(signal_2007), .B(cell_1977_and_out[0]), .Z(
        signal_2245) );
  XOR2_X1 cell_1977_U2 ( .A(signal_3421), .B(signal_3557), .Z(
        cell_1977_and_in[1]) );
  XOR2_X1 cell_1977_U1 ( .A(signal_2007), .B(signal_2119), .Z(
        cell_1977_and_in[0]) );
  XOR2_X1 cell_1977_a_HPC2_and_U14 ( .A(Fresh[263]), .B(cell_1977_and_in[0]), 
        .Z(cell_1977_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1977_a_HPC2_and_U13 ( .A(Fresh[263]), .B(cell_1977_and_in[1]), 
        .Z(cell_1977_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1977_a_HPC2_and_U12 ( .A1(cell_1977_a_HPC2_and_a_reg[1]), .A2(
        cell_1977_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1977_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1977_a_HPC2_and_U11 ( .A1(cell_1977_a_HPC2_and_a_reg[0]), .A2(
        cell_1977_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1977_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1977_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1977_a_HPC2_and_n9), 
        .ZN(cell_1977_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1977_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1977_a_HPC2_and_n9), 
        .ZN(cell_1977_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1977_a_HPC2_and_U8 ( .A(Fresh[263]), .ZN(cell_1977_a_HPC2_and_n9) );
  AND2_X1 cell_1977_a_HPC2_and_U7 ( .A1(cell_1977_and_in[1]), .A2(n448), .ZN(
        cell_1977_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1977_a_HPC2_and_U6 ( .A1(cell_1977_and_in[0]), .A2(n434), .ZN(
        cell_1977_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1977_a_HPC2_and_U5 ( .A(cell_1977_a_HPC2_and_n8), .B(
        cell_1977_a_HPC2_and_z_1__1_), .ZN(cell_1977_and_out[1]) );
  XNOR2_X1 cell_1977_a_HPC2_and_U4 ( .A(
        cell_1977_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1977_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1977_a_HPC2_and_n8) );
  XNOR2_X1 cell_1977_a_HPC2_and_U3 ( .A(cell_1977_a_HPC2_and_n7), .B(
        cell_1977_a_HPC2_and_z_0__0_), .ZN(cell_1977_and_out[0]) );
  XNOR2_X1 cell_1977_a_HPC2_and_U2 ( .A(
        cell_1977_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1977_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1977_a_HPC2_and_n7) );
  DFF_X1 cell_1977_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1977_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1977_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1977_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1977_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1977_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1977_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1977_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1977_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1977_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1978_U4 ( .A(signal_3525), .B(cell_1978_and_out[1]), .Z(
        signal_3756) );
  XOR2_X1 cell_1978_U3 ( .A(signal_2087), .B(cell_1978_and_out[0]), .Z(
        signal_2246) );
  XOR2_X1 cell_1978_U2 ( .A(signal_3525), .B(signal_3481), .Z(
        cell_1978_and_in[1]) );
  XOR2_X1 cell_1978_U1 ( .A(signal_2087), .B(signal_2043), .Z(
        cell_1978_and_in[0]) );
  XOR2_X1 cell_1978_a_HPC2_and_U14 ( .A(Fresh[264]), .B(cell_1978_and_in[0]), 
        .Z(cell_1978_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1978_a_HPC2_and_U13 ( .A(Fresh[264]), .B(cell_1978_and_in[1]), 
        .Z(cell_1978_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1978_a_HPC2_and_U12 ( .A1(cell_1978_a_HPC2_and_a_reg[1]), .A2(
        cell_1978_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1978_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1978_a_HPC2_and_U11 ( .A1(cell_1978_a_HPC2_and_a_reg[0]), .A2(
        cell_1978_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1978_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1978_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1978_a_HPC2_and_n9), 
        .ZN(cell_1978_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1978_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1978_a_HPC2_and_n9), 
        .ZN(cell_1978_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1978_a_HPC2_and_U8 ( .A(Fresh[264]), .ZN(cell_1978_a_HPC2_and_n9) );
  AND2_X1 cell_1978_a_HPC2_and_U7 ( .A1(cell_1978_and_in[1]), .A2(n454), .ZN(
        cell_1978_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1978_a_HPC2_and_U6 ( .A1(cell_1978_and_in[0]), .A2(n440), .ZN(
        cell_1978_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1978_a_HPC2_and_U5 ( .A(cell_1978_a_HPC2_and_n8), .B(
        cell_1978_a_HPC2_and_z_1__1_), .ZN(cell_1978_and_out[1]) );
  XNOR2_X1 cell_1978_a_HPC2_and_U4 ( .A(
        cell_1978_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1978_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1978_a_HPC2_and_n8) );
  XNOR2_X1 cell_1978_a_HPC2_and_U3 ( .A(cell_1978_a_HPC2_and_n7), .B(
        cell_1978_a_HPC2_and_z_0__0_), .ZN(cell_1978_and_out[0]) );
  XNOR2_X1 cell_1978_a_HPC2_and_U2 ( .A(
        cell_1978_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1978_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1978_a_HPC2_and_n7) );
  DFF_X1 cell_1978_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1978_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1978_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1978_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1978_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1978_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1978_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1978_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1978_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1978_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1979_U4 ( .A(signal_3490), .B(cell_1979_and_out[1]), .Z(
        signal_3757) );
  XOR2_X1 cell_1979_U3 ( .A(signal_2052), .B(cell_1979_and_out[0]), .Z(
        signal_2247) );
  XOR2_X1 cell_1979_U2 ( .A(signal_3490), .B(signal_3416), .Z(
        cell_1979_and_in[1]) );
  XOR2_X1 cell_1979_U1 ( .A(signal_2052), .B(signal_2002), .Z(
        cell_1979_and_in[0]) );
  XOR2_X1 cell_1979_a_HPC2_and_U14 ( .A(Fresh[265]), .B(cell_1979_and_in[0]), 
        .Z(cell_1979_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1979_a_HPC2_and_U13 ( .A(Fresh[265]), .B(cell_1979_and_in[1]), 
        .Z(cell_1979_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1979_a_HPC2_and_U12 ( .A1(cell_1979_a_HPC2_and_a_reg[1]), .A2(
        cell_1979_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1979_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1979_a_HPC2_and_U11 ( .A1(cell_1979_a_HPC2_and_a_reg[0]), .A2(
        cell_1979_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1979_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1979_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1979_a_HPC2_and_n9), 
        .ZN(cell_1979_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1979_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1979_a_HPC2_and_n9), 
        .ZN(cell_1979_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1979_a_HPC2_and_U8 ( .A(Fresh[265]), .ZN(cell_1979_a_HPC2_and_n9) );
  AND2_X1 cell_1979_a_HPC2_and_U7 ( .A1(cell_1979_and_in[1]), .A2(n454), .ZN(
        cell_1979_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1979_a_HPC2_and_U6 ( .A1(cell_1979_and_in[0]), .A2(n440), .ZN(
        cell_1979_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1979_a_HPC2_and_U5 ( .A(cell_1979_a_HPC2_and_n8), .B(
        cell_1979_a_HPC2_and_z_1__1_), .ZN(cell_1979_and_out[1]) );
  XNOR2_X1 cell_1979_a_HPC2_and_U4 ( .A(
        cell_1979_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1979_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1979_a_HPC2_and_n8) );
  XNOR2_X1 cell_1979_a_HPC2_and_U3 ( .A(cell_1979_a_HPC2_and_n7), .B(
        cell_1979_a_HPC2_and_z_0__0_), .ZN(cell_1979_and_out[0]) );
  XNOR2_X1 cell_1979_a_HPC2_and_U2 ( .A(
        cell_1979_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1979_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1979_a_HPC2_and_n7) );
  DFF_X1 cell_1979_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1979_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1979_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1979_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1979_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1979_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1979_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1979_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1979_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1979_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1980_U4 ( .A(signal_3486), .B(cell_1980_and_out[1]), .Z(
        signal_3758) );
  XOR2_X1 cell_1980_U3 ( .A(signal_2048), .B(cell_1980_and_out[0]), .Z(
        signal_2248) );
  XOR2_X1 cell_1980_U2 ( .A(signal_3486), .B(signal_3586), .Z(
        cell_1980_and_in[1]) );
  XOR2_X1 cell_1980_U1 ( .A(signal_2048), .B(signal_2148), .Z(
        cell_1980_and_in[0]) );
  XOR2_X1 cell_1980_a_HPC2_and_U14 ( .A(Fresh[266]), .B(cell_1980_and_in[0]), 
        .Z(cell_1980_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1980_a_HPC2_and_U13 ( .A(Fresh[266]), .B(cell_1980_and_in[1]), 
        .Z(cell_1980_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1980_a_HPC2_and_U12 ( .A1(cell_1980_a_HPC2_and_a_reg[1]), .A2(
        cell_1980_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1980_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1980_a_HPC2_and_U11 ( .A1(cell_1980_a_HPC2_and_a_reg[0]), .A2(
        cell_1980_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1980_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1980_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1980_a_HPC2_and_n9), 
        .ZN(cell_1980_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1980_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1980_a_HPC2_and_n9), 
        .ZN(cell_1980_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1980_a_HPC2_and_U8 ( .A(Fresh[266]), .ZN(cell_1980_a_HPC2_and_n9) );
  AND2_X1 cell_1980_a_HPC2_and_U7 ( .A1(cell_1980_and_in[1]), .A2(n448), .ZN(
        cell_1980_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1980_a_HPC2_and_U6 ( .A1(cell_1980_and_in[0]), .A2(n434), .ZN(
        cell_1980_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1980_a_HPC2_and_U5 ( .A(cell_1980_a_HPC2_and_n8), .B(
        cell_1980_a_HPC2_and_z_1__1_), .ZN(cell_1980_and_out[1]) );
  XNOR2_X1 cell_1980_a_HPC2_and_U4 ( .A(
        cell_1980_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1980_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1980_a_HPC2_and_n8) );
  XNOR2_X1 cell_1980_a_HPC2_and_U3 ( .A(cell_1980_a_HPC2_and_n7), .B(
        cell_1980_a_HPC2_and_z_0__0_), .ZN(cell_1980_and_out[0]) );
  XNOR2_X1 cell_1980_a_HPC2_and_U2 ( .A(
        cell_1980_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1980_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1980_a_HPC2_and_n7) );
  DFF_X1 cell_1980_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1980_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1980_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1980_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1980_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1980_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1980_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1980_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1980_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1980_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1981_U4 ( .A(signal_3508), .B(cell_1981_and_out[1]), .Z(
        signal_3759) );
  XOR2_X1 cell_1981_U3 ( .A(signal_2070), .B(cell_1981_and_out[0]), .Z(
        signal_2249) );
  XOR2_X1 cell_1981_U2 ( .A(signal_3508), .B(signal_3584), .Z(
        cell_1981_and_in[1]) );
  XOR2_X1 cell_1981_U1 ( .A(signal_2070), .B(signal_2146), .Z(
        cell_1981_and_in[0]) );
  XOR2_X1 cell_1981_a_HPC2_and_U14 ( .A(Fresh[267]), .B(cell_1981_and_in[0]), 
        .Z(cell_1981_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1981_a_HPC2_and_U13 ( .A(Fresh[267]), .B(cell_1981_and_in[1]), 
        .Z(cell_1981_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1981_a_HPC2_and_U12 ( .A1(cell_1981_a_HPC2_and_a_reg[1]), .A2(
        cell_1981_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1981_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1981_a_HPC2_and_U11 ( .A1(cell_1981_a_HPC2_and_a_reg[0]), .A2(
        cell_1981_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1981_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1981_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1981_a_HPC2_and_n9), 
        .ZN(cell_1981_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1981_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1981_a_HPC2_and_n9), 
        .ZN(cell_1981_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1981_a_HPC2_and_U8 ( .A(Fresh[267]), .ZN(cell_1981_a_HPC2_and_n9) );
  AND2_X1 cell_1981_a_HPC2_and_U7 ( .A1(cell_1981_and_in[1]), .A2(n448), .ZN(
        cell_1981_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1981_a_HPC2_and_U6 ( .A1(cell_1981_and_in[0]), .A2(n434), .ZN(
        cell_1981_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1981_a_HPC2_and_U5 ( .A(cell_1981_a_HPC2_and_n8), .B(
        cell_1981_a_HPC2_and_z_1__1_), .ZN(cell_1981_and_out[1]) );
  XNOR2_X1 cell_1981_a_HPC2_and_U4 ( .A(
        cell_1981_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1981_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1981_a_HPC2_and_n8) );
  XNOR2_X1 cell_1981_a_HPC2_and_U3 ( .A(cell_1981_a_HPC2_and_n7), .B(
        cell_1981_a_HPC2_and_z_0__0_), .ZN(cell_1981_and_out[0]) );
  XNOR2_X1 cell_1981_a_HPC2_and_U2 ( .A(
        cell_1981_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1981_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1981_a_HPC2_and_n7) );
  DFF_X1 cell_1981_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1981_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1981_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1981_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1981_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1981_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1981_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1981_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1981_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1981_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1982_U4 ( .A(signal_3549), .B(cell_1982_and_out[1]), .Z(
        signal_3760) );
  XOR2_X1 cell_1982_U3 ( .A(signal_2111), .B(cell_1982_and_out[0]), .Z(
        signal_2250) );
  XOR2_X1 cell_1982_U2 ( .A(signal_3549), .B(signal_3476), .Z(
        cell_1982_and_in[1]) );
  XOR2_X1 cell_1982_U1 ( .A(signal_2111), .B(signal_2038), .Z(
        cell_1982_and_in[0]) );
  XOR2_X1 cell_1982_a_HPC2_and_U14 ( .A(Fresh[268]), .B(cell_1982_and_in[0]), 
        .Z(cell_1982_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1982_a_HPC2_and_U13 ( .A(Fresh[268]), .B(cell_1982_and_in[1]), 
        .Z(cell_1982_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1982_a_HPC2_and_U12 ( .A1(cell_1982_a_HPC2_and_a_reg[1]), .A2(
        cell_1982_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1982_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1982_a_HPC2_and_U11 ( .A1(cell_1982_a_HPC2_and_a_reg[0]), .A2(
        cell_1982_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1982_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1982_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1982_a_HPC2_and_n9), 
        .ZN(cell_1982_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1982_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1982_a_HPC2_and_n9), 
        .ZN(cell_1982_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1982_a_HPC2_and_U8 ( .A(Fresh[268]), .ZN(cell_1982_a_HPC2_and_n9) );
  AND2_X1 cell_1982_a_HPC2_and_U7 ( .A1(cell_1982_and_in[1]), .A2(n448), .ZN(
        cell_1982_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1982_a_HPC2_and_U6 ( .A1(cell_1982_and_in[0]), .A2(n434), .ZN(
        cell_1982_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1982_a_HPC2_and_U5 ( .A(cell_1982_a_HPC2_and_n8), .B(
        cell_1982_a_HPC2_and_z_1__1_), .ZN(cell_1982_and_out[1]) );
  XNOR2_X1 cell_1982_a_HPC2_and_U4 ( .A(
        cell_1982_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1982_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1982_a_HPC2_and_n8) );
  XNOR2_X1 cell_1982_a_HPC2_and_U3 ( .A(cell_1982_a_HPC2_and_n7), .B(
        cell_1982_a_HPC2_and_z_0__0_), .ZN(cell_1982_and_out[0]) );
  XNOR2_X1 cell_1982_a_HPC2_and_U2 ( .A(
        cell_1982_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1982_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1982_a_HPC2_and_n7) );
  DFF_X1 cell_1982_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1982_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1982_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1982_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1982_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1982_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1982_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1982_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1982_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1982_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1983_U4 ( .A(n367), .B(cell_1983_and_out[1]), .Z(signal_3761)
         );
  XOR2_X1 cell_1983_U3 ( .A(n366), .B(cell_1983_and_out[0]), .Z(signal_2251)
         );
  XOR2_X1 cell_1983_U2 ( .A(n367), .B(signal_3539), .Z(cell_1983_and_in[1]) );
  XOR2_X1 cell_1983_U1 ( .A(n366), .B(signal_2101), .Z(cell_1983_and_in[0]) );
  XOR2_X1 cell_1983_a_HPC2_and_U14 ( .A(Fresh[269]), .B(cell_1983_and_in[0]), 
        .Z(cell_1983_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1983_a_HPC2_and_U13 ( .A(Fresh[269]), .B(cell_1983_and_in[1]), 
        .Z(cell_1983_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1983_a_HPC2_and_U12 ( .A1(cell_1983_a_HPC2_and_a_reg[1]), .A2(
        cell_1983_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1983_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1983_a_HPC2_and_U11 ( .A1(cell_1983_a_HPC2_and_a_reg[0]), .A2(
        cell_1983_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1983_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1983_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1983_a_HPC2_and_n9), 
        .ZN(cell_1983_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1983_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1983_a_HPC2_and_n9), 
        .ZN(cell_1983_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1983_a_HPC2_and_U8 ( .A(Fresh[269]), .ZN(cell_1983_a_HPC2_and_n9) );
  AND2_X1 cell_1983_a_HPC2_and_U7 ( .A1(cell_1983_and_in[1]), .A2(n448), .ZN(
        cell_1983_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1983_a_HPC2_and_U6 ( .A1(cell_1983_and_in[0]), .A2(n434), .ZN(
        cell_1983_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1983_a_HPC2_and_U5 ( .A(cell_1983_a_HPC2_and_n8), .B(
        cell_1983_a_HPC2_and_z_1__1_), .ZN(cell_1983_and_out[1]) );
  XNOR2_X1 cell_1983_a_HPC2_and_U4 ( .A(
        cell_1983_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1983_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1983_a_HPC2_and_n8) );
  XNOR2_X1 cell_1983_a_HPC2_and_U3 ( .A(cell_1983_a_HPC2_and_n7), .B(
        cell_1983_a_HPC2_and_z_0__0_), .ZN(cell_1983_and_out[0]) );
  XNOR2_X1 cell_1983_a_HPC2_and_U2 ( .A(
        cell_1983_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1983_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1983_a_HPC2_and_n7) );
  DFF_X1 cell_1983_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1983_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1983_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1983_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1983_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1983_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1983_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1983_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1983_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1983_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1984_U4 ( .A(signal_3503), .B(cell_1984_and_out[1]), .Z(
        signal_3762) );
  XOR2_X1 cell_1984_U3 ( .A(signal_2065), .B(cell_1984_and_out[0]), .Z(
        signal_2252) );
  XOR2_X1 cell_1984_U2 ( .A(signal_3503), .B(signal_3469), .Z(
        cell_1984_and_in[1]) );
  XOR2_X1 cell_1984_U1 ( .A(signal_2065), .B(signal_2031), .Z(
        cell_1984_and_in[0]) );
  XOR2_X1 cell_1984_a_HPC2_and_U14 ( .A(Fresh[270]), .B(cell_1984_and_in[0]), 
        .Z(cell_1984_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1984_a_HPC2_and_U13 ( .A(Fresh[270]), .B(cell_1984_and_in[1]), 
        .Z(cell_1984_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1984_a_HPC2_and_U12 ( .A1(cell_1984_a_HPC2_and_a_reg[1]), .A2(
        cell_1984_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1984_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1984_a_HPC2_and_U11 ( .A1(cell_1984_a_HPC2_and_a_reg[0]), .A2(
        cell_1984_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1984_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1984_a_HPC2_and_U10 ( .A1(n454), .A2(cell_1984_a_HPC2_and_n9), 
        .ZN(cell_1984_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1984_a_HPC2_and_U9 ( .A1(n440), .A2(cell_1984_a_HPC2_and_n9), 
        .ZN(cell_1984_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1984_a_HPC2_and_U8 ( .A(Fresh[270]), .ZN(cell_1984_a_HPC2_and_n9) );
  AND2_X1 cell_1984_a_HPC2_and_U7 ( .A1(cell_1984_and_in[1]), .A2(n454), .ZN(
        cell_1984_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1984_a_HPC2_and_U6 ( .A1(cell_1984_and_in[0]), .A2(n440), .ZN(
        cell_1984_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1984_a_HPC2_and_U5 ( .A(cell_1984_a_HPC2_and_n8), .B(
        cell_1984_a_HPC2_and_z_1__1_), .ZN(cell_1984_and_out[1]) );
  XNOR2_X1 cell_1984_a_HPC2_and_U4 ( .A(
        cell_1984_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1984_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1984_a_HPC2_and_n8) );
  XNOR2_X1 cell_1984_a_HPC2_and_U3 ( .A(cell_1984_a_HPC2_and_n7), .B(
        cell_1984_a_HPC2_and_z_0__0_), .ZN(cell_1984_and_out[0]) );
  XNOR2_X1 cell_1984_a_HPC2_and_U2 ( .A(
        cell_1984_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1984_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1984_a_HPC2_and_n7) );
  DFF_X1 cell_1984_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1984_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1984_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n440), .CK(clk), 
        .Q(cell_1984_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1984_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1984_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n454), .CK(clk), 
        .Q(cell_1984_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1984_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1984_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1984_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1985_U4 ( .A(signal_3480), .B(cell_1985_and_out[1]), .Z(
        signal_3763) );
  XOR2_X1 cell_1985_U3 ( .A(signal_2042), .B(cell_1985_and_out[0]), .Z(
        signal_2253) );
  XOR2_X1 cell_1985_U2 ( .A(signal_3480), .B(signal_3425), .Z(
        cell_1985_and_in[1]) );
  XOR2_X1 cell_1985_U1 ( .A(signal_2042), .B(signal_2011), .Z(
        cell_1985_and_in[0]) );
  XOR2_X1 cell_1985_a_HPC2_and_U14 ( .A(Fresh[271]), .B(cell_1985_and_in[0]), 
        .Z(cell_1985_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1985_a_HPC2_and_U13 ( .A(Fresh[271]), .B(cell_1985_and_in[1]), 
        .Z(cell_1985_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1985_a_HPC2_and_U12 ( .A1(cell_1985_a_HPC2_and_a_reg[1]), .A2(
        cell_1985_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1985_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1985_a_HPC2_and_U11 ( .A1(cell_1985_a_HPC2_and_a_reg[0]), .A2(
        cell_1985_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1985_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1985_a_HPC2_and_U10 ( .A1(n448), .A2(cell_1985_a_HPC2_and_n9), 
        .ZN(cell_1985_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1985_a_HPC2_and_U9 ( .A1(n434), .A2(cell_1985_a_HPC2_and_n9), 
        .ZN(cell_1985_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1985_a_HPC2_and_U8 ( .A(Fresh[271]), .ZN(cell_1985_a_HPC2_and_n9) );
  AND2_X1 cell_1985_a_HPC2_and_U7 ( .A1(cell_1985_and_in[1]), .A2(n448), .ZN(
        cell_1985_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1985_a_HPC2_and_U6 ( .A1(cell_1985_and_in[0]), .A2(n434), .ZN(
        cell_1985_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1985_a_HPC2_and_U5 ( .A(cell_1985_a_HPC2_and_n8), .B(
        cell_1985_a_HPC2_and_z_1__1_), .ZN(cell_1985_and_out[1]) );
  XNOR2_X1 cell_1985_a_HPC2_and_U4 ( .A(
        cell_1985_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1985_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1985_a_HPC2_and_n8) );
  XNOR2_X1 cell_1985_a_HPC2_and_U3 ( .A(cell_1985_a_HPC2_and_n7), .B(
        cell_1985_a_HPC2_and_z_0__0_), .ZN(cell_1985_and_out[0]) );
  XNOR2_X1 cell_1985_a_HPC2_and_U2 ( .A(
        cell_1985_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1985_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1985_a_HPC2_and_n7) );
  DFF_X1 cell_1985_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1985_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1985_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n434), .CK(clk), 
        .Q(cell_1985_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1985_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1985_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n448), .CK(clk), 
        .Q(cell_1985_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1985_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1985_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1985_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1986_U4 ( .A(signal_3541), .B(cell_1986_and_out[1]), .Z(
        signal_3764) );
  XOR2_X1 cell_1986_U3 ( .A(signal_2103), .B(cell_1986_and_out[0]), .Z(
        signal_2254) );
  XOR2_X1 cell_1986_U2 ( .A(signal_3541), .B(signal_3472), .Z(
        cell_1986_and_in[1]) );
  XOR2_X1 cell_1986_U1 ( .A(signal_2103), .B(signal_2034), .Z(
        cell_1986_and_in[0]) );
  XOR2_X1 cell_1986_a_HPC2_and_U14 ( .A(Fresh[272]), .B(cell_1986_and_in[0]), 
        .Z(cell_1986_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1986_a_HPC2_and_U13 ( .A(Fresh[272]), .B(cell_1986_and_in[1]), 
        .Z(cell_1986_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1986_a_HPC2_and_U12 ( .A1(cell_1986_a_HPC2_and_a_reg[1]), .A2(
        cell_1986_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1986_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1986_a_HPC2_and_U11 ( .A1(cell_1986_a_HPC2_and_a_reg[0]), .A2(
        cell_1986_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1986_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1986_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1986_a_HPC2_and_n9), 
        .ZN(cell_1986_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1986_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1986_a_HPC2_and_n9), 
        .ZN(cell_1986_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1986_a_HPC2_and_U8 ( .A(Fresh[272]), .ZN(cell_1986_a_HPC2_and_n9) );
  AND2_X1 cell_1986_a_HPC2_and_U7 ( .A1(cell_1986_and_in[1]), .A2(n449), .ZN(
        cell_1986_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1986_a_HPC2_and_U6 ( .A1(cell_1986_and_in[0]), .A2(n435), .ZN(
        cell_1986_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1986_a_HPC2_and_U5 ( .A(cell_1986_a_HPC2_and_n8), .B(
        cell_1986_a_HPC2_and_z_1__1_), .ZN(cell_1986_and_out[1]) );
  XNOR2_X1 cell_1986_a_HPC2_and_U4 ( .A(
        cell_1986_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1986_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1986_a_HPC2_and_n8) );
  XNOR2_X1 cell_1986_a_HPC2_and_U3 ( .A(cell_1986_a_HPC2_and_n7), .B(
        cell_1986_a_HPC2_and_z_0__0_), .ZN(cell_1986_and_out[0]) );
  XNOR2_X1 cell_1986_a_HPC2_and_U2 ( .A(
        cell_1986_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1986_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1986_a_HPC2_and_n7) );
  DFF_X1 cell_1986_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1986_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1986_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1986_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1986_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1986_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1986_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1986_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1986_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1986_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1987_U4 ( .A(signal_3484), .B(cell_1987_and_out[1]), .Z(
        signal_3765) );
  XOR2_X1 cell_1987_U3 ( .A(signal_2046), .B(cell_1987_and_out[0]), .Z(
        signal_2255) );
  XOR2_X1 cell_1987_U2 ( .A(signal_3484), .B(signal_3549), .Z(
        cell_1987_and_in[1]) );
  XOR2_X1 cell_1987_U1 ( .A(signal_2046), .B(signal_2111), .Z(
        cell_1987_and_in[0]) );
  XOR2_X1 cell_1987_a_HPC2_and_U14 ( .A(Fresh[273]), .B(cell_1987_and_in[0]), 
        .Z(cell_1987_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1987_a_HPC2_and_U13 ( .A(Fresh[273]), .B(cell_1987_and_in[1]), 
        .Z(cell_1987_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1987_a_HPC2_and_U12 ( .A1(cell_1987_a_HPC2_and_a_reg[1]), .A2(
        cell_1987_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1987_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1987_a_HPC2_and_U11 ( .A1(cell_1987_a_HPC2_and_a_reg[0]), .A2(
        cell_1987_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1987_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1987_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1987_a_HPC2_and_n9), 
        .ZN(cell_1987_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1987_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1987_a_HPC2_and_n9), 
        .ZN(cell_1987_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1987_a_HPC2_and_U8 ( .A(Fresh[273]), .ZN(cell_1987_a_HPC2_and_n9) );
  AND2_X1 cell_1987_a_HPC2_and_U7 ( .A1(cell_1987_and_in[1]), .A2(n449), .ZN(
        cell_1987_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1987_a_HPC2_and_U6 ( .A1(cell_1987_and_in[0]), .A2(n435), .ZN(
        cell_1987_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1987_a_HPC2_and_U5 ( .A(cell_1987_a_HPC2_and_n8), .B(
        cell_1987_a_HPC2_and_z_1__1_), .ZN(cell_1987_and_out[1]) );
  XNOR2_X1 cell_1987_a_HPC2_and_U4 ( .A(
        cell_1987_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1987_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1987_a_HPC2_and_n8) );
  XNOR2_X1 cell_1987_a_HPC2_and_U3 ( .A(cell_1987_a_HPC2_and_n7), .B(
        cell_1987_a_HPC2_and_z_0__0_), .ZN(cell_1987_and_out[0]) );
  XNOR2_X1 cell_1987_a_HPC2_and_U2 ( .A(
        cell_1987_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1987_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1987_a_HPC2_and_n7) );
  DFF_X1 cell_1987_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1987_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1987_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1987_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1987_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1987_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1987_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1987_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1987_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1987_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1988_U4 ( .A(signal_3531), .B(cell_1988_and_out[1]), .Z(
        signal_3766) );
  XOR2_X1 cell_1988_U3 ( .A(signal_2093), .B(cell_1988_and_out[0]), .Z(
        signal_2256) );
  XOR2_X1 cell_1988_U2 ( .A(signal_3531), .B(signal_3258), .Z(
        cell_1988_and_in[1]) );
  XOR2_X1 cell_1988_U1 ( .A(signal_2093), .B(signal_1984), .Z(
        cell_1988_and_in[0]) );
  XOR2_X1 cell_1988_a_HPC2_and_U14 ( .A(Fresh[274]), .B(cell_1988_and_in[0]), 
        .Z(cell_1988_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1988_a_HPC2_and_U13 ( .A(Fresh[274]), .B(cell_1988_and_in[1]), 
        .Z(cell_1988_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1988_a_HPC2_and_U12 ( .A1(cell_1988_a_HPC2_and_a_reg[1]), .A2(
        cell_1988_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1988_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1988_a_HPC2_and_U11 ( .A1(cell_1988_a_HPC2_and_a_reg[0]), .A2(
        cell_1988_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1988_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1988_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1988_a_HPC2_and_n9), 
        .ZN(cell_1988_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1988_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1988_a_HPC2_and_n9), 
        .ZN(cell_1988_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1988_a_HPC2_and_U8 ( .A(Fresh[274]), .ZN(cell_1988_a_HPC2_and_n9) );
  AND2_X1 cell_1988_a_HPC2_and_U7 ( .A1(cell_1988_and_in[1]), .A2(n449), .ZN(
        cell_1988_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1988_a_HPC2_and_U6 ( .A1(cell_1988_and_in[0]), .A2(n435), .ZN(
        cell_1988_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1988_a_HPC2_and_U5 ( .A(cell_1988_a_HPC2_and_n8), .B(
        cell_1988_a_HPC2_and_z_1__1_), .ZN(cell_1988_and_out[1]) );
  XNOR2_X1 cell_1988_a_HPC2_and_U4 ( .A(
        cell_1988_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1988_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1988_a_HPC2_and_n8) );
  XNOR2_X1 cell_1988_a_HPC2_and_U3 ( .A(cell_1988_a_HPC2_and_n7), .B(
        cell_1988_a_HPC2_and_z_0__0_), .ZN(cell_1988_and_out[0]) );
  XNOR2_X1 cell_1988_a_HPC2_and_U2 ( .A(
        cell_1988_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1988_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1988_a_HPC2_and_n7) );
  DFF_X1 cell_1988_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1988_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1988_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1988_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1988_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1988_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1988_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1988_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1988_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1988_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1989_U4 ( .A(signal_3464), .B(cell_1989_and_out[1]), .Z(
        signal_3767) );
  XOR2_X1 cell_1989_U3 ( .A(signal_2026), .B(cell_1989_and_out[0]), .Z(
        signal_2257) );
  XOR2_X1 cell_1989_U2 ( .A(signal_3464), .B(signal_3583), .Z(
        cell_1989_and_in[1]) );
  XOR2_X1 cell_1989_U1 ( .A(signal_2026), .B(signal_2145), .Z(
        cell_1989_and_in[0]) );
  XOR2_X1 cell_1989_a_HPC2_and_U14 ( .A(Fresh[275]), .B(cell_1989_and_in[0]), 
        .Z(cell_1989_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1989_a_HPC2_and_U13 ( .A(Fresh[275]), .B(cell_1989_and_in[1]), 
        .Z(cell_1989_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1989_a_HPC2_and_U12 ( .A1(cell_1989_a_HPC2_and_a_reg[1]), .A2(
        cell_1989_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1989_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1989_a_HPC2_and_U11 ( .A1(cell_1989_a_HPC2_and_a_reg[0]), .A2(
        cell_1989_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1989_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1989_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1989_a_HPC2_and_n9), 
        .ZN(cell_1989_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1989_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1989_a_HPC2_and_n9), 
        .ZN(cell_1989_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1989_a_HPC2_and_U8 ( .A(Fresh[275]), .ZN(cell_1989_a_HPC2_and_n9) );
  AND2_X1 cell_1989_a_HPC2_and_U7 ( .A1(cell_1989_and_in[1]), .A2(n449), .ZN(
        cell_1989_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1989_a_HPC2_and_U6 ( .A1(cell_1989_and_in[0]), .A2(n435), .ZN(
        cell_1989_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1989_a_HPC2_and_U5 ( .A(cell_1989_a_HPC2_and_n8), .B(
        cell_1989_a_HPC2_and_z_1__1_), .ZN(cell_1989_and_out[1]) );
  XNOR2_X1 cell_1989_a_HPC2_and_U4 ( .A(
        cell_1989_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1989_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1989_a_HPC2_and_n8) );
  XNOR2_X1 cell_1989_a_HPC2_and_U3 ( .A(cell_1989_a_HPC2_and_n7), .B(
        cell_1989_a_HPC2_and_z_0__0_), .ZN(cell_1989_and_out[0]) );
  XNOR2_X1 cell_1989_a_HPC2_and_U2 ( .A(
        cell_1989_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1989_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1989_a_HPC2_and_n7) );
  DFF_X1 cell_1989_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1989_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1989_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1989_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1989_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1989_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1989_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1989_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1989_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1989_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1990_U4 ( .A(signal_3552), .B(cell_1990_and_out[1]), .Z(
        signal_3768) );
  XOR2_X1 cell_1990_U3 ( .A(signal_2114), .B(cell_1990_and_out[0]), .Z(
        signal_2258) );
  XOR2_X1 cell_1990_U2 ( .A(signal_3552), .B(signal_3562), .Z(
        cell_1990_and_in[1]) );
  XOR2_X1 cell_1990_U1 ( .A(signal_2114), .B(signal_2124), .Z(
        cell_1990_and_in[0]) );
  XOR2_X1 cell_1990_a_HPC2_and_U14 ( .A(Fresh[276]), .B(cell_1990_and_in[0]), 
        .Z(cell_1990_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1990_a_HPC2_and_U13 ( .A(Fresh[276]), .B(cell_1990_and_in[1]), 
        .Z(cell_1990_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1990_a_HPC2_and_U12 ( .A1(cell_1990_a_HPC2_and_a_reg[1]), .A2(
        cell_1990_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1990_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1990_a_HPC2_and_U11 ( .A1(cell_1990_a_HPC2_and_a_reg[0]), .A2(
        cell_1990_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1990_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1990_a_HPC2_and_U10 ( .A1(n450), .A2(cell_1990_a_HPC2_and_n9), 
        .ZN(cell_1990_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1990_a_HPC2_and_U9 ( .A1(n436), .A2(cell_1990_a_HPC2_and_n9), 
        .ZN(cell_1990_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1990_a_HPC2_and_U8 ( .A(Fresh[276]), .ZN(cell_1990_a_HPC2_and_n9) );
  AND2_X1 cell_1990_a_HPC2_and_U7 ( .A1(cell_1990_and_in[1]), .A2(n450), .ZN(
        cell_1990_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1990_a_HPC2_and_U6 ( .A1(cell_1990_and_in[0]), .A2(n436), .ZN(
        cell_1990_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1990_a_HPC2_and_U5 ( .A(cell_1990_a_HPC2_and_n8), .B(
        cell_1990_a_HPC2_and_z_1__1_), .ZN(cell_1990_and_out[1]) );
  XNOR2_X1 cell_1990_a_HPC2_and_U4 ( .A(
        cell_1990_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1990_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1990_a_HPC2_and_n8) );
  XNOR2_X1 cell_1990_a_HPC2_and_U3 ( .A(cell_1990_a_HPC2_and_n7), .B(
        cell_1990_a_HPC2_and_z_0__0_), .ZN(cell_1990_and_out[0]) );
  XNOR2_X1 cell_1990_a_HPC2_and_U2 ( .A(
        cell_1990_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1990_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1990_a_HPC2_and_n7) );
  DFF_X1 cell_1990_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1990_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1990_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_1990_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1990_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1990_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_1990_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1990_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1990_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1990_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1991_U4 ( .A(signal_3515), .B(cell_1991_and_out[1]), .Z(
        signal_3769) );
  XOR2_X1 cell_1991_U3 ( .A(signal_2077), .B(cell_1991_and_out[0]), .Z(
        signal_2259) );
  XOR2_X1 cell_1991_U2 ( .A(signal_3515), .B(signal_3496), .Z(
        cell_1991_and_in[1]) );
  XOR2_X1 cell_1991_U1 ( .A(signal_2077), .B(signal_2058), .Z(
        cell_1991_and_in[0]) );
  XOR2_X1 cell_1991_a_HPC2_and_U14 ( .A(Fresh[277]), .B(cell_1991_and_in[0]), 
        .Z(cell_1991_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1991_a_HPC2_and_U13 ( .A(Fresh[277]), .B(cell_1991_and_in[1]), 
        .Z(cell_1991_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1991_a_HPC2_and_U12 ( .A1(cell_1991_a_HPC2_and_a_reg[1]), .A2(
        cell_1991_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1991_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1991_a_HPC2_and_U11 ( .A1(cell_1991_a_HPC2_and_a_reg[0]), .A2(
        cell_1991_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1991_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1991_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1991_a_HPC2_and_n9), 
        .ZN(cell_1991_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1991_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1991_a_HPC2_and_n9), 
        .ZN(cell_1991_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1991_a_HPC2_and_U8 ( .A(Fresh[277]), .ZN(cell_1991_a_HPC2_and_n9) );
  AND2_X1 cell_1991_a_HPC2_and_U7 ( .A1(cell_1991_and_in[1]), .A2(n442), .ZN(
        cell_1991_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1991_a_HPC2_and_U6 ( .A1(cell_1991_and_in[0]), .A2(n428), .ZN(
        cell_1991_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1991_a_HPC2_and_U5 ( .A(cell_1991_a_HPC2_and_n8), .B(
        cell_1991_a_HPC2_and_z_1__1_), .ZN(cell_1991_and_out[1]) );
  XNOR2_X1 cell_1991_a_HPC2_and_U4 ( .A(
        cell_1991_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1991_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1991_a_HPC2_and_n8) );
  XNOR2_X1 cell_1991_a_HPC2_and_U3 ( .A(cell_1991_a_HPC2_and_n7), .B(
        cell_1991_a_HPC2_and_z_0__0_), .ZN(cell_1991_and_out[0]) );
  XNOR2_X1 cell_1991_a_HPC2_and_U2 ( .A(
        cell_1991_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1991_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1991_a_HPC2_and_n7) );
  DFF_X1 cell_1991_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1991_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1991_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1991_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1991_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1991_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1991_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1991_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1991_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1991_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1992_U4 ( .A(signal_3524), .B(cell_1992_and_out[1]), .Z(
        signal_3770) );
  XOR2_X1 cell_1992_U3 ( .A(signal_2086), .B(cell_1992_and_out[0]), .Z(
        signal_2260) );
  XOR2_X1 cell_1992_U2 ( .A(signal_3524), .B(n365), .Z(cell_1992_and_in[1]) );
  XOR2_X1 cell_1992_U1 ( .A(signal_2086), .B(n363), .Z(cell_1992_and_in[0]) );
  XOR2_X1 cell_1992_a_HPC2_and_U14 ( .A(Fresh[278]), .B(cell_1992_and_in[0]), 
        .Z(cell_1992_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1992_a_HPC2_and_U13 ( .A(Fresh[278]), .B(cell_1992_and_in[1]), 
        .Z(cell_1992_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1992_a_HPC2_and_U12 ( .A1(cell_1992_a_HPC2_and_a_reg[1]), .A2(
        cell_1992_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1992_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1992_a_HPC2_and_U11 ( .A1(cell_1992_a_HPC2_and_a_reg[0]), .A2(
        cell_1992_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1992_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1992_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1992_a_HPC2_and_n9), 
        .ZN(cell_1992_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1992_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1992_a_HPC2_and_n9), 
        .ZN(cell_1992_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1992_a_HPC2_and_U8 ( .A(Fresh[278]), .ZN(cell_1992_a_HPC2_and_n9) );
  AND2_X1 cell_1992_a_HPC2_and_U7 ( .A1(cell_1992_and_in[1]), .A2(n449), .ZN(
        cell_1992_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1992_a_HPC2_and_U6 ( .A1(cell_1992_and_in[0]), .A2(n435), .ZN(
        cell_1992_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1992_a_HPC2_and_U5 ( .A(cell_1992_a_HPC2_and_n8), .B(
        cell_1992_a_HPC2_and_z_1__1_), .ZN(cell_1992_and_out[1]) );
  XNOR2_X1 cell_1992_a_HPC2_and_U4 ( .A(
        cell_1992_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1992_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1992_a_HPC2_and_n8) );
  XNOR2_X1 cell_1992_a_HPC2_and_U3 ( .A(cell_1992_a_HPC2_and_n7), .B(
        cell_1992_a_HPC2_and_z_0__0_), .ZN(cell_1992_and_out[0]) );
  XNOR2_X1 cell_1992_a_HPC2_and_U2 ( .A(
        cell_1992_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1992_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1992_a_HPC2_and_n7) );
  DFF_X1 cell_1992_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1992_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1992_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1992_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1992_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1992_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1992_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1992_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1992_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1992_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1993_U4 ( .A(signal_3480), .B(cell_1993_and_out[1]), .Z(
        signal_3771) );
  XOR2_X1 cell_1993_U3 ( .A(signal_2042), .B(cell_1993_and_out[0]), .Z(
        signal_2261) );
  XOR2_X1 cell_1993_U2 ( .A(signal_3480), .B(signal_3499), .Z(
        cell_1993_and_in[1]) );
  XOR2_X1 cell_1993_U1 ( .A(signal_2042), .B(signal_2061), .Z(
        cell_1993_and_in[0]) );
  XOR2_X1 cell_1993_a_HPC2_and_U14 ( .A(Fresh[279]), .B(cell_1993_and_in[0]), 
        .Z(cell_1993_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1993_a_HPC2_and_U13 ( .A(Fresh[279]), .B(cell_1993_and_in[1]), 
        .Z(cell_1993_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1993_a_HPC2_and_U12 ( .A1(cell_1993_a_HPC2_and_a_reg[1]), .A2(
        cell_1993_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1993_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1993_a_HPC2_and_U11 ( .A1(cell_1993_a_HPC2_and_a_reg[0]), .A2(
        cell_1993_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1993_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1993_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1993_a_HPC2_and_n9), 
        .ZN(cell_1993_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1993_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1993_a_HPC2_and_n9), 
        .ZN(cell_1993_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1993_a_HPC2_and_U8 ( .A(Fresh[279]), .ZN(cell_1993_a_HPC2_and_n9) );
  AND2_X1 cell_1993_a_HPC2_and_U7 ( .A1(cell_1993_and_in[1]), .A2(n449), .ZN(
        cell_1993_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1993_a_HPC2_and_U6 ( .A1(cell_1993_and_in[0]), .A2(n435), .ZN(
        cell_1993_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1993_a_HPC2_and_U5 ( .A(cell_1993_a_HPC2_and_n8), .B(
        cell_1993_a_HPC2_and_z_1__1_), .ZN(cell_1993_and_out[1]) );
  XNOR2_X1 cell_1993_a_HPC2_and_U4 ( .A(
        cell_1993_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1993_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1993_a_HPC2_and_n8) );
  XNOR2_X1 cell_1993_a_HPC2_and_U3 ( .A(cell_1993_a_HPC2_and_n7), .B(
        cell_1993_a_HPC2_and_z_0__0_), .ZN(cell_1993_and_out[0]) );
  XNOR2_X1 cell_1993_a_HPC2_and_U2 ( .A(
        cell_1993_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1993_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1993_a_HPC2_and_n7) );
  DFF_X1 cell_1993_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1993_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1993_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1993_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1993_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1993_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1993_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1993_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1993_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1993_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1994_U4 ( .A(signal_3494), .B(cell_1994_and_out[1]), .Z(
        signal_3772) );
  XOR2_X1 cell_1994_U3 ( .A(signal_2056), .B(cell_1994_and_out[0]), .Z(
        signal_2262) );
  XOR2_X1 cell_1994_U2 ( .A(signal_3494), .B(signal_3556), .Z(
        cell_1994_and_in[1]) );
  XOR2_X1 cell_1994_U1 ( .A(signal_2056), .B(signal_2118), .Z(
        cell_1994_and_in[0]) );
  XOR2_X1 cell_1994_a_HPC2_and_U14 ( .A(Fresh[280]), .B(cell_1994_and_in[0]), 
        .Z(cell_1994_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1994_a_HPC2_and_U13 ( .A(Fresh[280]), .B(cell_1994_and_in[1]), 
        .Z(cell_1994_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1994_a_HPC2_and_U12 ( .A1(cell_1994_a_HPC2_and_a_reg[1]), .A2(
        cell_1994_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1994_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1994_a_HPC2_and_U11 ( .A1(cell_1994_a_HPC2_and_a_reg[0]), .A2(
        cell_1994_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1994_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1994_a_HPC2_and_U10 ( .A1(signal_3235), .A2(
        cell_1994_a_HPC2_and_n9), .ZN(cell_1994_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1994_a_HPC2_and_U9 ( .A1(signal_1514), .A2(
        cell_1994_a_HPC2_and_n9), .ZN(cell_1994_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1994_a_HPC2_and_U8 ( .A(Fresh[280]), .ZN(cell_1994_a_HPC2_and_n9) );
  AND2_X1 cell_1994_a_HPC2_and_U7 ( .A1(cell_1994_and_in[1]), .A2(signal_3235), 
        .ZN(cell_1994_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1994_a_HPC2_and_U6 ( .A1(cell_1994_and_in[0]), .A2(signal_1514), 
        .ZN(cell_1994_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1994_a_HPC2_and_U5 ( .A(cell_1994_a_HPC2_and_n8), .B(
        cell_1994_a_HPC2_and_z_1__1_), .ZN(cell_1994_and_out[1]) );
  XNOR2_X1 cell_1994_a_HPC2_and_U4 ( .A(
        cell_1994_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1994_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1994_a_HPC2_and_n8) );
  XNOR2_X1 cell_1994_a_HPC2_and_U3 ( .A(cell_1994_a_HPC2_and_n7), .B(
        cell_1994_a_HPC2_and_z_0__0_), .ZN(cell_1994_and_out[0]) );
  XNOR2_X1 cell_1994_a_HPC2_and_U2 ( .A(
        cell_1994_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1994_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1994_a_HPC2_and_n7) );
  DFF_X1 cell_1994_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1994_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1994_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1514), 
        .CK(clk), .Q(cell_1994_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1994_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1994_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3235), 
        .CK(clk), .Q(cell_1994_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1994_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1994_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1994_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1995_U4 ( .A(signal_3510), .B(cell_1995_and_out[1]), .Z(
        signal_3773) );
  XOR2_X1 cell_1995_U3 ( .A(signal_2072), .B(cell_1995_and_out[0]), .Z(
        signal_2263) );
  XOR2_X1 cell_1995_U2 ( .A(signal_3510), .B(signal_3506), .Z(
        cell_1995_and_in[1]) );
  XOR2_X1 cell_1995_U1 ( .A(signal_2072), .B(signal_2068), .Z(
        cell_1995_and_in[0]) );
  XOR2_X1 cell_1995_a_HPC2_and_U14 ( .A(Fresh[281]), .B(cell_1995_and_in[0]), 
        .Z(cell_1995_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1995_a_HPC2_and_U13 ( .A(Fresh[281]), .B(cell_1995_and_in[1]), 
        .Z(cell_1995_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1995_a_HPC2_and_U12 ( .A1(cell_1995_a_HPC2_and_a_reg[1]), .A2(
        cell_1995_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1995_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1995_a_HPC2_and_U11 ( .A1(cell_1995_a_HPC2_and_a_reg[0]), .A2(
        cell_1995_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1995_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1995_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1995_a_HPC2_and_n9), 
        .ZN(cell_1995_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1995_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1995_a_HPC2_and_n9), 
        .ZN(cell_1995_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1995_a_HPC2_and_U8 ( .A(Fresh[281]), .ZN(cell_1995_a_HPC2_and_n9) );
  AND2_X1 cell_1995_a_HPC2_and_U7 ( .A1(cell_1995_and_in[1]), .A2(n449), .ZN(
        cell_1995_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1995_a_HPC2_and_U6 ( .A1(cell_1995_and_in[0]), .A2(n435), .ZN(
        cell_1995_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1995_a_HPC2_and_U5 ( .A(cell_1995_a_HPC2_and_n8), .B(
        cell_1995_a_HPC2_and_z_1__1_), .ZN(cell_1995_and_out[1]) );
  XNOR2_X1 cell_1995_a_HPC2_and_U4 ( .A(
        cell_1995_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1995_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1995_a_HPC2_and_n8) );
  XNOR2_X1 cell_1995_a_HPC2_and_U3 ( .A(cell_1995_a_HPC2_and_n7), .B(
        cell_1995_a_HPC2_and_z_0__0_), .ZN(cell_1995_and_out[0]) );
  XNOR2_X1 cell_1995_a_HPC2_and_U2 ( .A(
        cell_1995_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1995_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1995_a_HPC2_and_n7) );
  DFF_X1 cell_1995_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1995_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1995_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1995_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1995_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1995_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1995_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1995_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1995_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1995_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1996_U4 ( .A(n389), .B(cell_1996_and_out[1]), .Z(signal_3774)
         );
  XOR2_X1 cell_1996_U3 ( .A(n388), .B(cell_1996_and_out[0]), .Z(signal_2264)
         );
  XOR2_X1 cell_1996_U2 ( .A(n389), .B(signal_3512), .Z(cell_1996_and_in[1]) );
  XOR2_X1 cell_1996_U1 ( .A(n388), .B(signal_2074), .Z(cell_1996_and_in[0]) );
  XOR2_X1 cell_1996_a_HPC2_and_U14 ( .A(Fresh[282]), .B(cell_1996_and_in[0]), 
        .Z(cell_1996_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1996_a_HPC2_and_U13 ( .A(Fresh[282]), .B(cell_1996_and_in[1]), 
        .Z(cell_1996_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1996_a_HPC2_and_U12 ( .A1(cell_1996_a_HPC2_and_a_reg[1]), .A2(
        cell_1996_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1996_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1996_a_HPC2_and_U11 ( .A1(cell_1996_a_HPC2_and_a_reg[0]), .A2(
        cell_1996_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1996_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1996_a_HPC2_and_U10 ( .A1(n449), .A2(cell_1996_a_HPC2_and_n9), 
        .ZN(cell_1996_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1996_a_HPC2_and_U9 ( .A1(n435), .A2(cell_1996_a_HPC2_and_n9), 
        .ZN(cell_1996_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1996_a_HPC2_and_U8 ( .A(Fresh[282]), .ZN(cell_1996_a_HPC2_and_n9) );
  AND2_X1 cell_1996_a_HPC2_and_U7 ( .A1(cell_1996_and_in[1]), .A2(n449), .ZN(
        cell_1996_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1996_a_HPC2_and_U6 ( .A1(cell_1996_and_in[0]), .A2(n435), .ZN(
        cell_1996_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1996_a_HPC2_and_U5 ( .A(cell_1996_a_HPC2_and_n8), .B(
        cell_1996_a_HPC2_and_z_1__1_), .ZN(cell_1996_and_out[1]) );
  XNOR2_X1 cell_1996_a_HPC2_and_U4 ( .A(
        cell_1996_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1996_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1996_a_HPC2_and_n8) );
  XNOR2_X1 cell_1996_a_HPC2_and_U3 ( .A(cell_1996_a_HPC2_and_n7), .B(
        cell_1996_a_HPC2_and_z_0__0_), .ZN(cell_1996_and_out[0]) );
  XNOR2_X1 cell_1996_a_HPC2_and_U2 ( .A(
        cell_1996_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1996_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1996_a_HPC2_and_n7) );
  DFF_X1 cell_1996_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1996_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1996_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n435), .CK(clk), 
        .Q(cell_1996_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1996_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1996_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n449), .CK(clk), 
        .Q(cell_1996_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1996_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1996_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1996_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1997_U4 ( .A(signal_3529), .B(cell_1997_and_out[1]), .Z(
        signal_3775) );
  XOR2_X1 cell_1997_U3 ( .A(signal_2091), .B(cell_1997_and_out[0]), .Z(
        signal_2265) );
  XOR2_X1 cell_1997_U2 ( .A(signal_3529), .B(signal_3553), .Z(
        cell_1997_and_in[1]) );
  XOR2_X1 cell_1997_U1 ( .A(signal_2091), .B(signal_2115), .Z(
        cell_1997_and_in[0]) );
  XOR2_X1 cell_1997_a_HPC2_and_U14 ( .A(Fresh[283]), .B(cell_1997_and_in[0]), 
        .Z(cell_1997_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1997_a_HPC2_and_U13 ( .A(Fresh[283]), .B(cell_1997_and_in[1]), 
        .Z(cell_1997_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1997_a_HPC2_and_U12 ( .A1(cell_1997_a_HPC2_and_a_reg[1]), .A2(
        cell_1997_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1997_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1997_a_HPC2_and_U11 ( .A1(cell_1997_a_HPC2_and_a_reg[0]), .A2(
        cell_1997_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1997_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1997_a_HPC2_and_U10 ( .A1(n443), .A2(cell_1997_a_HPC2_and_n9), 
        .ZN(cell_1997_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1997_a_HPC2_and_U9 ( .A1(n429), .A2(cell_1997_a_HPC2_and_n9), 
        .ZN(cell_1997_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1997_a_HPC2_and_U8 ( .A(Fresh[283]), .ZN(cell_1997_a_HPC2_and_n9) );
  AND2_X1 cell_1997_a_HPC2_and_U7 ( .A1(cell_1997_and_in[1]), .A2(n443), .ZN(
        cell_1997_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1997_a_HPC2_and_U6 ( .A1(cell_1997_and_in[0]), .A2(n429), .ZN(
        cell_1997_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1997_a_HPC2_and_U5 ( .A(cell_1997_a_HPC2_and_n8), .B(
        cell_1997_a_HPC2_and_z_1__1_), .ZN(cell_1997_and_out[1]) );
  XNOR2_X1 cell_1997_a_HPC2_and_U4 ( .A(
        cell_1997_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1997_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1997_a_HPC2_and_n8) );
  XNOR2_X1 cell_1997_a_HPC2_and_U3 ( .A(cell_1997_a_HPC2_and_n7), .B(
        cell_1997_a_HPC2_and_z_0__0_), .ZN(cell_1997_and_out[0]) );
  XNOR2_X1 cell_1997_a_HPC2_and_U2 ( .A(
        cell_1997_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1997_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1997_a_HPC2_and_n7) );
  DFF_X1 cell_1997_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1997_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1997_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n429), .CK(clk), 
        .Q(cell_1997_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1997_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1997_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n443), .CK(clk), 
        .Q(cell_1997_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1997_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1997_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1997_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1998_U4 ( .A(signal_3467), .B(cell_1998_and_out[1]), .Z(
        signal_3776) );
  XOR2_X1 cell_1998_U3 ( .A(signal_2029), .B(cell_1998_and_out[0]), .Z(
        signal_2266) );
  XOR2_X1 cell_1998_U2 ( .A(signal_3467), .B(signal_3459), .Z(
        cell_1998_and_in[1]) );
  XOR2_X1 cell_1998_U1 ( .A(signal_2029), .B(signal_2021), .Z(
        cell_1998_and_in[0]) );
  XOR2_X1 cell_1998_a_HPC2_and_U14 ( .A(Fresh[284]), .B(cell_1998_and_in[0]), 
        .Z(cell_1998_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1998_a_HPC2_and_U13 ( .A(Fresh[284]), .B(cell_1998_and_in[1]), 
        .Z(cell_1998_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1998_a_HPC2_and_U12 ( .A1(cell_1998_a_HPC2_and_a_reg[1]), .A2(
        cell_1998_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1998_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1998_a_HPC2_and_U11 ( .A1(cell_1998_a_HPC2_and_a_reg[0]), .A2(
        cell_1998_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1998_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1998_a_HPC2_and_U10 ( .A1(n442), .A2(cell_1998_a_HPC2_and_n9), 
        .ZN(cell_1998_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1998_a_HPC2_and_U9 ( .A1(n428), .A2(cell_1998_a_HPC2_and_n9), 
        .ZN(cell_1998_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1998_a_HPC2_and_U8 ( .A(Fresh[284]), .ZN(cell_1998_a_HPC2_and_n9) );
  AND2_X1 cell_1998_a_HPC2_and_U7 ( .A1(cell_1998_and_in[1]), .A2(n442), .ZN(
        cell_1998_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1998_a_HPC2_and_U6 ( .A1(cell_1998_and_in[0]), .A2(n428), .ZN(
        cell_1998_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1998_a_HPC2_and_U5 ( .A(cell_1998_a_HPC2_and_n8), .B(
        cell_1998_a_HPC2_and_z_1__1_), .ZN(cell_1998_and_out[1]) );
  XNOR2_X1 cell_1998_a_HPC2_and_U4 ( .A(
        cell_1998_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1998_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1998_a_HPC2_and_n8) );
  XNOR2_X1 cell_1998_a_HPC2_and_U3 ( .A(cell_1998_a_HPC2_and_n7), .B(
        cell_1998_a_HPC2_and_z_0__0_), .ZN(cell_1998_and_out[0]) );
  XNOR2_X1 cell_1998_a_HPC2_and_U2 ( .A(
        cell_1998_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1998_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1998_a_HPC2_and_n7) );
  DFF_X1 cell_1998_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1998_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1998_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n428), .CK(clk), 
        .Q(cell_1998_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1998_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1998_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n442), .CK(clk), 
        .Q(cell_1998_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1998_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1998_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1998_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_1999_U4 ( .A(signal_3575), .B(cell_1999_and_out[1]), .Z(
        signal_3777) );
  XOR2_X1 cell_1999_U3 ( .A(signal_2137), .B(cell_1999_and_out[0]), .Z(
        signal_2267) );
  XOR2_X1 cell_1999_U2 ( .A(signal_3575), .B(signal_3503), .Z(
        cell_1999_and_in[1]) );
  XOR2_X1 cell_1999_U1 ( .A(signal_2137), .B(signal_2065), .Z(
        cell_1999_and_in[0]) );
  XOR2_X1 cell_1999_a_HPC2_and_U14 ( .A(Fresh[285]), .B(cell_1999_and_in[0]), 
        .Z(cell_1999_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_1999_a_HPC2_and_U13 ( .A(Fresh[285]), .B(cell_1999_and_in[1]), 
        .Z(cell_1999_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_1999_a_HPC2_and_U12 ( .A1(cell_1999_a_HPC2_and_a_reg[1]), .A2(
        cell_1999_a_HPC2_and_s_out_1__0_), .ZN(
        cell_1999_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_1999_a_HPC2_and_U11 ( .A1(cell_1999_a_HPC2_and_a_reg[0]), .A2(
        cell_1999_a_HPC2_and_s_out_0__1_), .ZN(
        cell_1999_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_1999_a_HPC2_and_U10 ( .A1(n450), .A2(cell_1999_a_HPC2_and_n9), 
        .ZN(cell_1999_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_1999_a_HPC2_and_U9 ( .A1(n436), .A2(cell_1999_a_HPC2_and_n9), 
        .ZN(cell_1999_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_1999_a_HPC2_and_U8 ( .A(Fresh[285]), .ZN(cell_1999_a_HPC2_and_n9) );
  AND2_X1 cell_1999_a_HPC2_and_U7 ( .A1(cell_1999_and_in[1]), .A2(n450), .ZN(
        cell_1999_a_HPC2_and_mul[1]) );
  AND2_X1 cell_1999_a_HPC2_and_U6 ( .A1(cell_1999_and_in[0]), .A2(n436), .ZN(
        cell_1999_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_1999_a_HPC2_and_U5 ( .A(cell_1999_a_HPC2_and_n8), .B(
        cell_1999_a_HPC2_and_z_1__1_), .ZN(cell_1999_and_out[1]) );
  XNOR2_X1 cell_1999_a_HPC2_and_U4 ( .A(
        cell_1999_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_1999_a_HPC2_and_p_1_out_1__0_), .ZN(cell_1999_a_HPC2_and_n8) );
  XNOR2_X1 cell_1999_a_HPC2_and_U3 ( .A(cell_1999_a_HPC2_and_n7), .B(
        cell_1999_a_HPC2_and_z_0__0_), .ZN(cell_1999_and_out[0]) );
  XNOR2_X1 cell_1999_a_HPC2_and_U2 ( .A(
        cell_1999_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_1999_a_HPC2_and_p_1_out_0__1_), .ZN(cell_1999_a_HPC2_and_n7) );
  DFF_X1 cell_1999_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_1999_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_1999_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_1999_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_1999_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_1999_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_1999_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_1999_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_1999_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_1999_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2000_U4 ( .A(signal_3516), .B(cell_2000_and_out[1]), .Z(
        signal_3778) );
  XOR2_X1 cell_2000_U3 ( .A(signal_2078), .B(cell_2000_and_out[0]), .Z(
        signal_2268) );
  XOR2_X1 cell_2000_U2 ( .A(signal_3516), .B(signal_3484), .Z(
        cell_2000_and_in[1]) );
  XOR2_X1 cell_2000_U1 ( .A(signal_2078), .B(signal_2046), .Z(
        cell_2000_and_in[0]) );
  XOR2_X1 cell_2000_a_HPC2_and_U14 ( .A(Fresh[286]), .B(cell_2000_and_in[0]), 
        .Z(cell_2000_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2000_a_HPC2_and_U13 ( .A(Fresh[286]), .B(cell_2000_and_in[1]), 
        .Z(cell_2000_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2000_a_HPC2_and_U12 ( .A1(cell_2000_a_HPC2_and_a_reg[1]), .A2(
        cell_2000_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2000_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2000_a_HPC2_and_U11 ( .A1(cell_2000_a_HPC2_and_a_reg[0]), .A2(
        cell_2000_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2000_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2000_a_HPC2_and_U10 ( .A1(n450), .A2(cell_2000_a_HPC2_and_n9), 
        .ZN(cell_2000_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2000_a_HPC2_and_U9 ( .A1(n436), .A2(cell_2000_a_HPC2_and_n9), 
        .ZN(cell_2000_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2000_a_HPC2_and_U8 ( .A(Fresh[286]), .ZN(cell_2000_a_HPC2_and_n9) );
  AND2_X1 cell_2000_a_HPC2_and_U7 ( .A1(cell_2000_and_in[1]), .A2(n450), .ZN(
        cell_2000_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2000_a_HPC2_and_U6 ( .A1(cell_2000_and_in[0]), .A2(n436), .ZN(
        cell_2000_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2000_a_HPC2_and_U5 ( .A(cell_2000_a_HPC2_and_n8), .B(
        cell_2000_a_HPC2_and_z_1__1_), .ZN(cell_2000_and_out[1]) );
  XNOR2_X1 cell_2000_a_HPC2_and_U4 ( .A(
        cell_2000_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2000_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2000_a_HPC2_and_n8) );
  XNOR2_X1 cell_2000_a_HPC2_and_U3 ( .A(cell_2000_a_HPC2_and_n7), .B(
        cell_2000_a_HPC2_and_z_0__0_), .ZN(cell_2000_and_out[0]) );
  XNOR2_X1 cell_2000_a_HPC2_and_U2 ( .A(
        cell_2000_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2000_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2000_a_HPC2_and_n7) );
  DFF_X1 cell_2000_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2000_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2000_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_2000_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2000_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2000_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_2000_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2000_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2000_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2000_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2001_U4 ( .A(signal_3480), .B(cell_2001_and_out[1]), .Z(
        signal_3779) );
  XOR2_X1 cell_2001_U3 ( .A(signal_2042), .B(cell_2001_and_out[0]), .Z(
        signal_2269) );
  XOR2_X1 cell_2001_U2 ( .A(signal_3480), .B(signal_3462), .Z(
        cell_2001_and_in[1]) );
  XOR2_X1 cell_2001_U1 ( .A(signal_2042), .B(signal_2024), .Z(
        cell_2001_and_in[0]) );
  XOR2_X1 cell_2001_a_HPC2_and_U14 ( .A(Fresh[287]), .B(cell_2001_and_in[0]), 
        .Z(cell_2001_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2001_a_HPC2_and_U13 ( .A(Fresh[287]), .B(cell_2001_and_in[1]), 
        .Z(cell_2001_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2001_a_HPC2_and_U12 ( .A1(cell_2001_a_HPC2_and_a_reg[1]), .A2(
        cell_2001_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2001_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2001_a_HPC2_and_U11 ( .A1(cell_2001_a_HPC2_and_a_reg[0]), .A2(
        cell_2001_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2001_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2001_a_HPC2_and_U10 ( .A1(n450), .A2(cell_2001_a_HPC2_and_n9), 
        .ZN(cell_2001_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2001_a_HPC2_and_U9 ( .A1(n436), .A2(cell_2001_a_HPC2_and_n9), 
        .ZN(cell_2001_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2001_a_HPC2_and_U8 ( .A(Fresh[287]), .ZN(cell_2001_a_HPC2_and_n9) );
  AND2_X1 cell_2001_a_HPC2_and_U7 ( .A1(cell_2001_and_in[1]), .A2(n450), .ZN(
        cell_2001_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2001_a_HPC2_and_U6 ( .A1(cell_2001_and_in[0]), .A2(n436), .ZN(
        cell_2001_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2001_a_HPC2_and_U5 ( .A(cell_2001_a_HPC2_and_n8), .B(
        cell_2001_a_HPC2_and_z_1__1_), .ZN(cell_2001_and_out[1]) );
  XNOR2_X1 cell_2001_a_HPC2_and_U4 ( .A(
        cell_2001_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2001_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2001_a_HPC2_and_n8) );
  XNOR2_X1 cell_2001_a_HPC2_and_U3 ( .A(cell_2001_a_HPC2_and_n7), .B(
        cell_2001_a_HPC2_and_z_0__0_), .ZN(cell_2001_and_out[0]) );
  XNOR2_X1 cell_2001_a_HPC2_and_U2 ( .A(
        cell_2001_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2001_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2001_a_HPC2_and_n7) );
  DFF_X1 cell_2001_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2001_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2001_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_2001_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2001_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2001_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_2001_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2001_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2001_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2001_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2002_U4 ( .A(signal_3488), .B(cell_2002_and_out[1]), .Z(
        signal_3780) );
  XOR2_X1 cell_2002_U3 ( .A(signal_2050), .B(cell_2002_and_out[0]), .Z(
        signal_2270) );
  XOR2_X1 cell_2002_U2 ( .A(signal_3488), .B(signal_3516), .Z(
        cell_2002_and_in[1]) );
  XOR2_X1 cell_2002_U1 ( .A(signal_2050), .B(signal_2078), .Z(
        cell_2002_and_in[0]) );
  XOR2_X1 cell_2002_a_HPC2_and_U14 ( .A(Fresh[288]), .B(cell_2002_and_in[0]), 
        .Z(cell_2002_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2002_a_HPC2_and_U13 ( .A(Fresh[288]), .B(cell_2002_and_in[1]), 
        .Z(cell_2002_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2002_a_HPC2_and_U12 ( .A1(cell_2002_a_HPC2_and_a_reg[1]), .A2(
        cell_2002_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2002_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2002_a_HPC2_and_U11 ( .A1(cell_2002_a_HPC2_and_a_reg[0]), .A2(
        cell_2002_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2002_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2002_a_HPC2_and_U10 ( .A1(n450), .A2(cell_2002_a_HPC2_and_n9), 
        .ZN(cell_2002_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2002_a_HPC2_and_U9 ( .A1(n436), .A2(cell_2002_a_HPC2_and_n9), 
        .ZN(cell_2002_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2002_a_HPC2_and_U8 ( .A(Fresh[288]), .ZN(cell_2002_a_HPC2_and_n9) );
  AND2_X1 cell_2002_a_HPC2_and_U7 ( .A1(cell_2002_and_in[1]), .A2(n450), .ZN(
        cell_2002_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2002_a_HPC2_and_U6 ( .A1(cell_2002_and_in[0]), .A2(n436), .ZN(
        cell_2002_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2002_a_HPC2_and_U5 ( .A(cell_2002_a_HPC2_and_n8), .B(
        cell_2002_a_HPC2_and_z_1__1_), .ZN(cell_2002_and_out[1]) );
  XNOR2_X1 cell_2002_a_HPC2_and_U4 ( .A(
        cell_2002_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2002_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2002_a_HPC2_and_n8) );
  XNOR2_X1 cell_2002_a_HPC2_and_U3 ( .A(cell_2002_a_HPC2_and_n7), .B(
        cell_2002_a_HPC2_and_z_0__0_), .ZN(cell_2002_and_out[0]) );
  XNOR2_X1 cell_2002_a_HPC2_and_U2 ( .A(
        cell_2002_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2002_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2002_a_HPC2_and_n7) );
  DFF_X1 cell_2002_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2002_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2002_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_2002_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2002_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2002_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_2002_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2002_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2002_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2002_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2003_U4 ( .A(signal_3461), .B(cell_2003_and_out[1]), .Z(
        signal_3781) );
  XOR2_X1 cell_2003_U3 ( .A(signal_2023), .B(cell_2003_and_out[0]), .Z(
        signal_2271) );
  XOR2_X1 cell_2003_U2 ( .A(signal_3461), .B(signal_3415), .Z(
        cell_2003_and_in[1]) );
  XOR2_X1 cell_2003_U1 ( .A(signal_2023), .B(signal_2001), .Z(
        cell_2003_and_in[0]) );
  XOR2_X1 cell_2003_a_HPC2_and_U14 ( .A(Fresh[289]), .B(cell_2003_and_in[0]), 
        .Z(cell_2003_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2003_a_HPC2_and_U13 ( .A(Fresh[289]), .B(cell_2003_and_in[1]), 
        .Z(cell_2003_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2003_a_HPC2_and_U12 ( .A1(cell_2003_a_HPC2_and_a_reg[1]), .A2(
        cell_2003_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2003_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2003_a_HPC2_and_U11 ( .A1(cell_2003_a_HPC2_and_a_reg[0]), .A2(
        cell_2003_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2003_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2003_a_HPC2_and_U10 ( .A1(n450), .A2(cell_2003_a_HPC2_and_n9), 
        .ZN(cell_2003_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2003_a_HPC2_and_U9 ( .A1(n436), .A2(cell_2003_a_HPC2_and_n9), 
        .ZN(cell_2003_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2003_a_HPC2_and_U8 ( .A(Fresh[289]), .ZN(cell_2003_a_HPC2_and_n9) );
  AND2_X1 cell_2003_a_HPC2_and_U7 ( .A1(cell_2003_and_in[1]), .A2(n450), .ZN(
        cell_2003_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2003_a_HPC2_and_U6 ( .A1(cell_2003_and_in[0]), .A2(n436), .ZN(
        cell_2003_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2003_a_HPC2_and_U5 ( .A(cell_2003_a_HPC2_and_n8), .B(
        cell_2003_a_HPC2_and_z_1__1_), .ZN(cell_2003_and_out[1]) );
  XNOR2_X1 cell_2003_a_HPC2_and_U4 ( .A(
        cell_2003_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2003_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2003_a_HPC2_and_n8) );
  XNOR2_X1 cell_2003_a_HPC2_and_U3 ( .A(cell_2003_a_HPC2_and_n7), .B(
        cell_2003_a_HPC2_and_z_0__0_), .ZN(cell_2003_and_out[0]) );
  XNOR2_X1 cell_2003_a_HPC2_and_U2 ( .A(
        cell_2003_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2003_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2003_a_HPC2_and_n7) );
  DFF_X1 cell_2003_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2003_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2003_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_2003_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2003_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2003_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_2003_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2003_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2003_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2003_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2004_U4 ( .A(signal_3465), .B(cell_2004_and_out[1]), .Z(
        signal_3782) );
  XOR2_X1 cell_2004_U3 ( .A(signal_2027), .B(cell_2004_and_out[0]), .Z(
        signal_2272) );
  XOR2_X1 cell_2004_U2 ( .A(signal_3465), .B(signal_3554), .Z(
        cell_2004_and_in[1]) );
  XOR2_X1 cell_2004_U1 ( .A(signal_2027), .B(signal_2116), .Z(
        cell_2004_and_in[0]) );
  XOR2_X1 cell_2004_a_HPC2_and_U14 ( .A(Fresh[290]), .B(cell_2004_and_in[0]), 
        .Z(cell_2004_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2004_a_HPC2_and_U13 ( .A(Fresh[290]), .B(cell_2004_and_in[1]), 
        .Z(cell_2004_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2004_a_HPC2_and_U12 ( .A1(cell_2004_a_HPC2_and_a_reg[1]), .A2(
        cell_2004_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2004_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2004_a_HPC2_and_U11 ( .A1(cell_2004_a_HPC2_and_a_reg[0]), .A2(
        cell_2004_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2004_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2004_a_HPC2_and_U10 ( .A1(n444), .A2(cell_2004_a_HPC2_and_n9), 
        .ZN(cell_2004_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2004_a_HPC2_and_U9 ( .A1(n430), .A2(cell_2004_a_HPC2_and_n9), 
        .ZN(cell_2004_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2004_a_HPC2_and_U8 ( .A(Fresh[290]), .ZN(cell_2004_a_HPC2_and_n9) );
  AND2_X1 cell_2004_a_HPC2_and_U7 ( .A1(cell_2004_and_in[1]), .A2(n444), .ZN(
        cell_2004_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2004_a_HPC2_and_U6 ( .A1(cell_2004_and_in[0]), .A2(n430), .ZN(
        cell_2004_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2004_a_HPC2_and_U5 ( .A(cell_2004_a_HPC2_and_n8), .B(
        cell_2004_a_HPC2_and_z_1__1_), .ZN(cell_2004_and_out[1]) );
  XNOR2_X1 cell_2004_a_HPC2_and_U4 ( .A(
        cell_2004_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2004_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2004_a_HPC2_and_n8) );
  XNOR2_X1 cell_2004_a_HPC2_and_U3 ( .A(cell_2004_a_HPC2_and_n7), .B(
        cell_2004_a_HPC2_and_z_0__0_), .ZN(cell_2004_and_out[0]) );
  XNOR2_X1 cell_2004_a_HPC2_and_U2 ( .A(
        cell_2004_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2004_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2004_a_HPC2_and_n7) );
  DFF_X1 cell_2004_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2004_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2004_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n430), .CK(clk), 
        .Q(cell_2004_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2004_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2004_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n444), .CK(clk), 
        .Q(cell_2004_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2004_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2004_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2004_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2005_U4 ( .A(signal_3505), .B(cell_2005_and_out[1]), .Z(
        signal_3783) );
  XOR2_X1 cell_2005_U3 ( .A(signal_2067), .B(cell_2005_and_out[0]), .Z(
        signal_2273) );
  XOR2_X1 cell_2005_U2 ( .A(signal_3505), .B(signal_3473), .Z(
        cell_2005_and_in[1]) );
  XOR2_X1 cell_2005_U1 ( .A(signal_2067), .B(signal_2035), .Z(
        cell_2005_and_in[0]) );
  XOR2_X1 cell_2005_a_HPC2_and_U14 ( .A(Fresh[291]), .B(cell_2005_and_in[0]), 
        .Z(cell_2005_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2005_a_HPC2_and_U13 ( .A(Fresh[291]), .B(cell_2005_and_in[1]), 
        .Z(cell_2005_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2005_a_HPC2_and_U12 ( .A1(cell_2005_a_HPC2_and_a_reg[1]), .A2(
        cell_2005_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2005_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2005_a_HPC2_and_U11 ( .A1(cell_2005_a_HPC2_and_a_reg[0]), .A2(
        cell_2005_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2005_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2005_a_HPC2_and_U10 ( .A1(n455), .A2(cell_2005_a_HPC2_and_n9), 
        .ZN(cell_2005_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2005_a_HPC2_and_U9 ( .A1(n441), .A2(cell_2005_a_HPC2_and_n9), 
        .ZN(cell_2005_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2005_a_HPC2_and_U8 ( .A(Fresh[291]), .ZN(cell_2005_a_HPC2_and_n9) );
  AND2_X1 cell_2005_a_HPC2_and_U7 ( .A1(cell_2005_and_in[1]), .A2(n455), .ZN(
        cell_2005_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2005_a_HPC2_and_U6 ( .A1(cell_2005_and_in[0]), .A2(n441), .ZN(
        cell_2005_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2005_a_HPC2_and_U5 ( .A(cell_2005_a_HPC2_and_n8), .B(
        cell_2005_a_HPC2_and_z_1__1_), .ZN(cell_2005_and_out[1]) );
  XNOR2_X1 cell_2005_a_HPC2_and_U4 ( .A(
        cell_2005_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2005_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2005_a_HPC2_and_n8) );
  XNOR2_X1 cell_2005_a_HPC2_and_U3 ( .A(cell_2005_a_HPC2_and_n7), .B(
        cell_2005_a_HPC2_and_z_0__0_), .ZN(cell_2005_and_out[0]) );
  XNOR2_X1 cell_2005_a_HPC2_and_U2 ( .A(
        cell_2005_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2005_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2005_a_HPC2_and_n7) );
  DFF_X1 cell_2005_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2005_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2005_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_2005_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2005_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2005_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_2005_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2005_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2005_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2005_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2006_U4 ( .A(signal_3524), .B(cell_2006_and_out[1]), .Z(
        signal_3784) );
  XOR2_X1 cell_2006_U3 ( .A(signal_2086), .B(cell_2006_and_out[0]), .Z(
        signal_2274) );
  XOR2_X1 cell_2006_U2 ( .A(signal_3524), .B(signal_3492), .Z(
        cell_2006_and_in[1]) );
  XOR2_X1 cell_2006_U1 ( .A(signal_2086), .B(signal_2054), .Z(
        cell_2006_and_in[0]) );
  XOR2_X1 cell_2006_a_HPC2_and_U14 ( .A(Fresh[292]), .B(cell_2006_and_in[0]), 
        .Z(cell_2006_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2006_a_HPC2_and_U13 ( .A(Fresh[292]), .B(cell_2006_and_in[1]), 
        .Z(cell_2006_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2006_a_HPC2_and_U12 ( .A1(cell_2006_a_HPC2_and_a_reg[1]), .A2(
        cell_2006_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2006_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2006_a_HPC2_and_U11 ( .A1(cell_2006_a_HPC2_and_a_reg[0]), .A2(
        cell_2006_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2006_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2006_a_HPC2_and_U10 ( .A1(n455), .A2(cell_2006_a_HPC2_and_n9), 
        .ZN(cell_2006_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2006_a_HPC2_and_U9 ( .A1(n441), .A2(cell_2006_a_HPC2_and_n9), 
        .ZN(cell_2006_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2006_a_HPC2_and_U8 ( .A(Fresh[292]), .ZN(cell_2006_a_HPC2_and_n9) );
  AND2_X1 cell_2006_a_HPC2_and_U7 ( .A1(cell_2006_and_in[1]), .A2(n455), .ZN(
        cell_2006_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2006_a_HPC2_and_U6 ( .A1(cell_2006_and_in[0]), .A2(n441), .ZN(
        cell_2006_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2006_a_HPC2_and_U5 ( .A(cell_2006_a_HPC2_and_n8), .B(
        cell_2006_a_HPC2_and_z_1__1_), .ZN(cell_2006_and_out[1]) );
  XNOR2_X1 cell_2006_a_HPC2_and_U4 ( .A(
        cell_2006_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2006_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2006_a_HPC2_and_n8) );
  XNOR2_X1 cell_2006_a_HPC2_and_U3 ( .A(cell_2006_a_HPC2_and_n7), .B(
        cell_2006_a_HPC2_and_z_0__0_), .ZN(cell_2006_and_out[0]) );
  XNOR2_X1 cell_2006_a_HPC2_and_U2 ( .A(
        cell_2006_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2006_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2006_a_HPC2_and_n7) );
  DFF_X1 cell_2006_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2006_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2006_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n441), .CK(clk), 
        .Q(cell_2006_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2006_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2006_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n455), .CK(clk), 
        .Q(cell_2006_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2006_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2006_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2006_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2007_U4 ( .A(signal_3578), .B(cell_2007_and_out[1]), .Z(
        signal_3785) );
  XOR2_X1 cell_2007_U3 ( .A(signal_2140), .B(cell_2007_and_out[0]), .Z(
        signal_2275) );
  XOR2_X1 cell_2007_U2 ( .A(signal_3578), .B(signal_3527), .Z(
        cell_2007_and_in[1]) );
  XOR2_X1 cell_2007_U1 ( .A(signal_2140), .B(signal_2089), .Z(
        cell_2007_and_in[0]) );
  XOR2_X1 cell_2007_a_HPC2_and_U14 ( .A(Fresh[293]), .B(cell_2007_and_in[0]), 
        .Z(cell_2007_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2007_a_HPC2_and_U13 ( .A(Fresh[293]), .B(cell_2007_and_in[1]), 
        .Z(cell_2007_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2007_a_HPC2_and_U12 ( .A1(cell_2007_a_HPC2_and_a_reg[1]), .A2(
        cell_2007_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2007_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2007_a_HPC2_and_U11 ( .A1(cell_2007_a_HPC2_and_a_reg[0]), .A2(
        cell_2007_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2007_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2007_a_HPC2_and_U10 ( .A1(n450), .A2(cell_2007_a_HPC2_and_n9), 
        .ZN(cell_2007_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2007_a_HPC2_and_U9 ( .A1(n436), .A2(cell_2007_a_HPC2_and_n9), 
        .ZN(cell_2007_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2007_a_HPC2_and_U8 ( .A(Fresh[293]), .ZN(cell_2007_a_HPC2_and_n9) );
  AND2_X1 cell_2007_a_HPC2_and_U7 ( .A1(cell_2007_and_in[1]), .A2(n450), .ZN(
        cell_2007_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2007_a_HPC2_and_U6 ( .A1(cell_2007_and_in[0]), .A2(n436), .ZN(
        cell_2007_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2007_a_HPC2_and_U5 ( .A(cell_2007_a_HPC2_and_n8), .B(
        cell_2007_a_HPC2_and_z_1__1_), .ZN(cell_2007_and_out[1]) );
  XNOR2_X1 cell_2007_a_HPC2_and_U4 ( .A(
        cell_2007_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2007_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2007_a_HPC2_and_n8) );
  XNOR2_X1 cell_2007_a_HPC2_and_U3 ( .A(cell_2007_a_HPC2_and_n7), .B(
        cell_2007_a_HPC2_and_z_0__0_), .ZN(cell_2007_and_out[0]) );
  XNOR2_X1 cell_2007_a_HPC2_and_U2 ( .A(
        cell_2007_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2007_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2007_a_HPC2_and_n7) );
  DFF_X1 cell_2007_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2007_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2007_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n436), .CK(clk), 
        .Q(cell_2007_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2007_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2007_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n450), .CK(clk), 
        .Q(cell_2007_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2007_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2007_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2007_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2008_U4 ( .A(signal_3742), .B(cell_2008_and_out[1]), .Z(
        signal_3922) );
  XOR2_X1 cell_2008_U3 ( .A(signal_2232), .B(cell_2008_and_out[0]), .Z(
        signal_2276) );
  XOR2_X1 cell_2008_U2 ( .A(signal_3742), .B(signal_3722), .Z(
        cell_2008_and_in[1]) );
  XOR2_X1 cell_2008_U1 ( .A(signal_2232), .B(signal_2212), .Z(
        cell_2008_and_in[0]) );
  XOR2_X1 cell_2008_a_HPC2_and_U14 ( .A(Fresh[294]), .B(cell_2008_and_in[0]), 
        .Z(cell_2008_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2008_a_HPC2_and_U13 ( .A(Fresh[294]), .B(cell_2008_and_in[1]), 
        .Z(cell_2008_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2008_a_HPC2_and_U12 ( .A1(cell_2008_a_HPC2_and_a_reg[1]), .A2(
        cell_2008_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2008_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2008_a_HPC2_and_U11 ( .A1(cell_2008_a_HPC2_and_a_reg[0]), .A2(
        cell_2008_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2008_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2008_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2008_a_HPC2_and_n9), 
        .ZN(cell_2008_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2008_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2008_a_HPC2_and_n9), 
        .ZN(cell_2008_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2008_a_HPC2_and_U8 ( .A(Fresh[294]), .ZN(cell_2008_a_HPC2_and_n9) );
  AND2_X1 cell_2008_a_HPC2_and_U7 ( .A1(cell_2008_and_in[1]), .A2(n466), .ZN(
        cell_2008_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2008_a_HPC2_and_U6 ( .A1(cell_2008_and_in[0]), .A2(n462), .ZN(
        cell_2008_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2008_a_HPC2_and_U5 ( .A(cell_2008_a_HPC2_and_n8), .B(
        cell_2008_a_HPC2_and_z_1__1_), .ZN(cell_2008_and_out[1]) );
  XNOR2_X1 cell_2008_a_HPC2_and_U4 ( .A(
        cell_2008_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2008_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2008_a_HPC2_and_n8) );
  XNOR2_X1 cell_2008_a_HPC2_and_U3 ( .A(cell_2008_a_HPC2_and_n7), .B(
        cell_2008_a_HPC2_and_z_0__0_), .ZN(cell_2008_and_out[0]) );
  XNOR2_X1 cell_2008_a_HPC2_and_U2 ( .A(
        cell_2008_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2008_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2008_a_HPC2_and_n7) );
  DFF_X1 cell_2008_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2008_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2008_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2008_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2008_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2008_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2008_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2008_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2008_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2008_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2009_U4 ( .A(signal_3783), .B(cell_2009_and_out[1]), .Z(
        signal_3923) );
  XOR2_X1 cell_2009_U3 ( .A(signal_2273), .B(cell_2009_and_out[0]), .Z(
        signal_2277) );
  XOR2_X1 cell_2009_U2 ( .A(signal_3783), .B(signal_3754), .Z(
        cell_2009_and_in[1]) );
  XOR2_X1 cell_2009_U1 ( .A(signal_2273), .B(signal_2244), .Z(
        cell_2009_and_in[0]) );
  XOR2_X1 cell_2009_a_HPC2_and_U14 ( .A(Fresh[295]), .B(cell_2009_and_in[0]), 
        .Z(cell_2009_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2009_a_HPC2_and_U13 ( .A(Fresh[295]), .B(cell_2009_and_in[1]), 
        .Z(cell_2009_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2009_a_HPC2_and_U12 ( .A1(cell_2009_a_HPC2_and_a_reg[1]), .A2(
        cell_2009_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2009_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2009_a_HPC2_and_U11 ( .A1(cell_2009_a_HPC2_and_a_reg[0]), .A2(
        cell_2009_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2009_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2009_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2009_a_HPC2_and_n9), 
        .ZN(cell_2009_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2009_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2009_a_HPC2_and_n9), 
        .ZN(cell_2009_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2009_a_HPC2_and_U8 ( .A(Fresh[295]), .ZN(cell_2009_a_HPC2_and_n9) );
  AND2_X1 cell_2009_a_HPC2_and_U7 ( .A1(cell_2009_and_in[1]), .A2(n466), .ZN(
        cell_2009_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2009_a_HPC2_and_U6 ( .A1(cell_2009_and_in[0]), .A2(n462), .ZN(
        cell_2009_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2009_a_HPC2_and_U5 ( .A(cell_2009_a_HPC2_and_n8), .B(
        cell_2009_a_HPC2_and_z_1__1_), .ZN(cell_2009_and_out[1]) );
  XNOR2_X1 cell_2009_a_HPC2_and_U4 ( .A(
        cell_2009_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2009_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2009_a_HPC2_and_n8) );
  XNOR2_X1 cell_2009_a_HPC2_and_U3 ( .A(cell_2009_a_HPC2_and_n7), .B(
        cell_2009_a_HPC2_and_z_0__0_), .ZN(cell_2009_and_out[0]) );
  XNOR2_X1 cell_2009_a_HPC2_and_U2 ( .A(
        cell_2009_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2009_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2009_a_HPC2_and_n7) );
  DFF_X1 cell_2009_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2009_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2009_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2009_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2009_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2009_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2009_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2009_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2009_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2009_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2010_U4 ( .A(signal_3723), .B(cell_2010_and_out[1]), .Z(
        signal_3924) );
  XOR2_X1 cell_2010_U3 ( .A(signal_2213), .B(cell_2010_and_out[0]), .Z(
        signal_2278) );
  XOR2_X1 cell_2010_U2 ( .A(signal_3723), .B(signal_3667), .Z(
        cell_2010_and_in[1]) );
  XOR2_X1 cell_2010_U1 ( .A(signal_2213), .B(signal_2157), .Z(
        cell_2010_and_in[0]) );
  XOR2_X1 cell_2010_a_HPC2_and_U14 ( .A(Fresh[296]), .B(cell_2010_and_in[0]), 
        .Z(cell_2010_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2010_a_HPC2_and_U13 ( .A(Fresh[296]), .B(cell_2010_and_in[1]), 
        .Z(cell_2010_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2010_a_HPC2_and_U12 ( .A1(cell_2010_a_HPC2_and_a_reg[1]), .A2(
        cell_2010_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2010_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2010_a_HPC2_and_U11 ( .A1(cell_2010_a_HPC2_and_a_reg[0]), .A2(
        cell_2010_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2010_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2010_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2010_a_HPC2_and_n9), 
        .ZN(cell_2010_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2010_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2010_a_HPC2_and_n9), 
        .ZN(cell_2010_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2010_a_HPC2_and_U8 ( .A(Fresh[296]), .ZN(cell_2010_a_HPC2_and_n9) );
  AND2_X1 cell_2010_a_HPC2_and_U7 ( .A1(cell_2010_and_in[1]), .A2(n466), .ZN(
        cell_2010_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2010_a_HPC2_and_U6 ( .A1(cell_2010_and_in[0]), .A2(n462), .ZN(
        cell_2010_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2010_a_HPC2_and_U5 ( .A(cell_2010_a_HPC2_and_n8), .B(
        cell_2010_a_HPC2_and_z_1__1_), .ZN(cell_2010_and_out[1]) );
  XNOR2_X1 cell_2010_a_HPC2_and_U4 ( .A(
        cell_2010_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2010_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2010_a_HPC2_and_n8) );
  XNOR2_X1 cell_2010_a_HPC2_and_U3 ( .A(cell_2010_a_HPC2_and_n7), .B(
        cell_2010_a_HPC2_and_z_0__0_), .ZN(cell_2010_and_out[0]) );
  XNOR2_X1 cell_2010_a_HPC2_and_U2 ( .A(
        cell_2010_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2010_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2010_a_HPC2_and_n7) );
  DFF_X1 cell_2010_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2010_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2010_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2010_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2010_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2010_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2010_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2010_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2010_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2010_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2011_U4 ( .A(signal_3743), .B(cell_2011_and_out[1]), .Z(
        signal_3925) );
  XOR2_X1 cell_2011_U3 ( .A(signal_2233), .B(cell_2011_and_out[0]), .Z(
        signal_2279) );
  XOR2_X1 cell_2011_U2 ( .A(signal_3743), .B(signal_3692), .Z(
        cell_2011_and_in[1]) );
  XOR2_X1 cell_2011_U1 ( .A(signal_2233), .B(signal_2182), .Z(
        cell_2011_and_in[0]) );
  XOR2_X1 cell_2011_a_HPC2_and_U14 ( .A(Fresh[297]), .B(cell_2011_and_in[0]), 
        .Z(cell_2011_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2011_a_HPC2_and_U13 ( .A(Fresh[297]), .B(cell_2011_and_in[1]), 
        .Z(cell_2011_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2011_a_HPC2_and_U12 ( .A1(cell_2011_a_HPC2_and_a_reg[1]), .A2(
        cell_2011_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2011_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2011_a_HPC2_and_U11 ( .A1(cell_2011_a_HPC2_and_a_reg[0]), .A2(
        cell_2011_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2011_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2011_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2011_a_HPC2_and_n9), 
        .ZN(cell_2011_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2011_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2011_a_HPC2_and_n9), 
        .ZN(cell_2011_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2011_a_HPC2_and_U8 ( .A(Fresh[297]), .ZN(cell_2011_a_HPC2_and_n9) );
  AND2_X1 cell_2011_a_HPC2_and_U7 ( .A1(cell_2011_and_in[1]), .A2(n466), .ZN(
        cell_2011_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2011_a_HPC2_and_U6 ( .A1(cell_2011_and_in[0]), .A2(n462), .ZN(
        cell_2011_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2011_a_HPC2_and_U5 ( .A(cell_2011_a_HPC2_and_n8), .B(
        cell_2011_a_HPC2_and_z_1__1_), .ZN(cell_2011_and_out[1]) );
  XNOR2_X1 cell_2011_a_HPC2_and_U4 ( .A(
        cell_2011_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2011_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2011_a_HPC2_and_n8) );
  XNOR2_X1 cell_2011_a_HPC2_and_U3 ( .A(cell_2011_a_HPC2_and_n7), .B(
        cell_2011_a_HPC2_and_z_0__0_), .ZN(cell_2011_and_out[0]) );
  XNOR2_X1 cell_2011_a_HPC2_and_U2 ( .A(
        cell_2011_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2011_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2011_a_HPC2_and_n7) );
  DFF_X1 cell_2011_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2011_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2011_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2011_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2011_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2011_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2011_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2011_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2011_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2011_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2012_U4 ( .A(signal_3712), .B(cell_2012_and_out[1]), .Z(
        signal_3926) );
  XOR2_X1 cell_2012_U3 ( .A(signal_2202), .B(cell_2012_and_out[0]), .Z(
        signal_2280) );
  XOR2_X1 cell_2012_U2 ( .A(signal_3712), .B(signal_3774), .Z(
        cell_2012_and_in[1]) );
  XOR2_X1 cell_2012_U1 ( .A(signal_2202), .B(signal_2264), .Z(
        cell_2012_and_in[0]) );
  XOR2_X1 cell_2012_a_HPC2_and_U14 ( .A(Fresh[298]), .B(cell_2012_and_in[0]), 
        .Z(cell_2012_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2012_a_HPC2_and_U13 ( .A(Fresh[298]), .B(cell_2012_and_in[1]), 
        .Z(cell_2012_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2012_a_HPC2_and_U12 ( .A1(cell_2012_a_HPC2_and_a_reg[1]), .A2(
        cell_2012_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2012_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2012_a_HPC2_and_U11 ( .A1(cell_2012_a_HPC2_and_a_reg[0]), .A2(
        cell_2012_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2012_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2012_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2012_a_HPC2_and_n9), 
        .ZN(cell_2012_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2012_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2012_a_HPC2_and_n9), 
        .ZN(cell_2012_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2012_a_HPC2_and_U8 ( .A(Fresh[298]), .ZN(cell_2012_a_HPC2_and_n9) );
  AND2_X1 cell_2012_a_HPC2_and_U7 ( .A1(cell_2012_and_in[1]), .A2(n466), .ZN(
        cell_2012_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2012_a_HPC2_and_U6 ( .A1(cell_2012_and_in[0]), .A2(n462), .ZN(
        cell_2012_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2012_a_HPC2_and_U5 ( .A(cell_2012_a_HPC2_and_n8), .B(
        cell_2012_a_HPC2_and_z_1__1_), .ZN(cell_2012_and_out[1]) );
  XNOR2_X1 cell_2012_a_HPC2_and_U4 ( .A(
        cell_2012_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2012_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2012_a_HPC2_and_n8) );
  XNOR2_X1 cell_2012_a_HPC2_and_U3 ( .A(cell_2012_a_HPC2_and_n7), .B(
        cell_2012_a_HPC2_and_z_0__0_), .ZN(cell_2012_and_out[0]) );
  XNOR2_X1 cell_2012_a_HPC2_and_U2 ( .A(
        cell_2012_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2012_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2012_a_HPC2_and_n7) );
  DFF_X1 cell_2012_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2012_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2012_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2012_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2012_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2012_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2012_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2012_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2012_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2012_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2013_U4 ( .A(signal_3780), .B(cell_2013_and_out[1]), .Z(
        signal_3927) );
  XOR2_X1 cell_2013_U3 ( .A(signal_2270), .B(cell_2013_and_out[0]), .Z(
        signal_2281) );
  XOR2_X1 cell_2013_U2 ( .A(signal_3780), .B(signal_3747), .Z(
        cell_2013_and_in[1]) );
  XOR2_X1 cell_2013_U1 ( .A(signal_2270), .B(signal_2237), .Z(
        cell_2013_and_in[0]) );
  XOR2_X1 cell_2013_a_HPC2_and_U14 ( .A(Fresh[299]), .B(cell_2013_and_in[0]), 
        .Z(cell_2013_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2013_a_HPC2_and_U13 ( .A(Fresh[299]), .B(cell_2013_and_in[1]), 
        .Z(cell_2013_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2013_a_HPC2_and_U12 ( .A1(cell_2013_a_HPC2_and_a_reg[1]), .A2(
        cell_2013_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2013_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2013_a_HPC2_and_U11 ( .A1(cell_2013_a_HPC2_and_a_reg[0]), .A2(
        cell_2013_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2013_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2013_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2013_a_HPC2_and_n9), 
        .ZN(cell_2013_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2013_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2013_a_HPC2_and_n9), 
        .ZN(cell_2013_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2013_a_HPC2_and_U8 ( .A(Fresh[299]), .ZN(cell_2013_a_HPC2_and_n9) );
  AND2_X1 cell_2013_a_HPC2_and_U7 ( .A1(cell_2013_and_in[1]), .A2(n466), .ZN(
        cell_2013_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2013_a_HPC2_and_U6 ( .A1(cell_2013_and_in[0]), .A2(n462), .ZN(
        cell_2013_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2013_a_HPC2_and_U5 ( .A(cell_2013_a_HPC2_and_n8), .B(
        cell_2013_a_HPC2_and_z_1__1_), .ZN(cell_2013_and_out[1]) );
  XNOR2_X1 cell_2013_a_HPC2_and_U4 ( .A(
        cell_2013_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2013_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2013_a_HPC2_and_n8) );
  XNOR2_X1 cell_2013_a_HPC2_and_U3 ( .A(cell_2013_a_HPC2_and_n7), .B(
        cell_2013_a_HPC2_and_z_0__0_), .ZN(cell_2013_and_out[0]) );
  XNOR2_X1 cell_2013_a_HPC2_and_U2 ( .A(
        cell_2013_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2013_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2013_a_HPC2_and_n7) );
  DFF_X1 cell_2013_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2013_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2013_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2013_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2013_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2013_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2013_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2013_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2013_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2013_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2014_U4 ( .A(signal_3750), .B(cell_2014_and_out[1]), .Z(
        signal_3928) );
  XOR2_X1 cell_2014_U3 ( .A(signal_2240), .B(cell_2014_and_out[0]), .Z(
        signal_2282) );
  XOR2_X1 cell_2014_U2 ( .A(signal_3750), .B(signal_3765), .Z(
        cell_2014_and_in[1]) );
  XOR2_X1 cell_2014_U1 ( .A(signal_2240), .B(signal_2255), .Z(
        cell_2014_and_in[0]) );
  XOR2_X1 cell_2014_a_HPC2_and_U14 ( .A(Fresh[300]), .B(cell_2014_and_in[0]), 
        .Z(cell_2014_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2014_a_HPC2_and_U13 ( .A(Fresh[300]), .B(cell_2014_and_in[1]), 
        .Z(cell_2014_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2014_a_HPC2_and_U12 ( .A1(cell_2014_a_HPC2_and_a_reg[1]), .A2(
        cell_2014_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2014_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2014_a_HPC2_and_U11 ( .A1(cell_2014_a_HPC2_and_a_reg[0]), .A2(
        cell_2014_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2014_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2014_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2014_a_HPC2_and_n9), 
        .ZN(cell_2014_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2014_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2014_a_HPC2_and_n9), 
        .ZN(cell_2014_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2014_a_HPC2_and_U8 ( .A(Fresh[300]), .ZN(cell_2014_a_HPC2_and_n9) );
  AND2_X1 cell_2014_a_HPC2_and_U7 ( .A1(cell_2014_and_in[1]), .A2(n466), .ZN(
        cell_2014_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2014_a_HPC2_and_U6 ( .A1(cell_2014_and_in[0]), .A2(n462), .ZN(
        cell_2014_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2014_a_HPC2_and_U5 ( .A(cell_2014_a_HPC2_and_n8), .B(
        cell_2014_a_HPC2_and_z_1__1_), .ZN(cell_2014_and_out[1]) );
  XNOR2_X1 cell_2014_a_HPC2_and_U4 ( .A(
        cell_2014_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2014_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2014_a_HPC2_and_n8) );
  XNOR2_X1 cell_2014_a_HPC2_and_U3 ( .A(cell_2014_a_HPC2_and_n7), .B(
        cell_2014_a_HPC2_and_z_0__0_), .ZN(cell_2014_and_out[0]) );
  XNOR2_X1 cell_2014_a_HPC2_and_U2 ( .A(
        cell_2014_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2014_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2014_a_HPC2_and_n7) );
  DFF_X1 cell_2014_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2014_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2014_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2014_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2014_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2014_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2014_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2014_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2014_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2014_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2015_U4 ( .A(signal_3769), .B(cell_2015_and_out[1]), .Z(
        signal_3929) );
  XOR2_X1 cell_2015_U3 ( .A(signal_2259), .B(cell_2015_and_out[0]), .Z(
        signal_2283) );
  XOR2_X1 cell_2015_U2 ( .A(signal_3769), .B(signal_3724), .Z(
        cell_2015_and_in[1]) );
  XOR2_X1 cell_2015_U1 ( .A(signal_2259), .B(signal_2214), .Z(
        cell_2015_and_in[0]) );
  XOR2_X1 cell_2015_a_HPC2_and_U14 ( .A(Fresh[301]), .B(cell_2015_and_in[0]), 
        .Z(cell_2015_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2015_a_HPC2_and_U13 ( .A(Fresh[301]), .B(cell_2015_and_in[1]), 
        .Z(cell_2015_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2015_a_HPC2_and_U12 ( .A1(cell_2015_a_HPC2_and_a_reg[1]), .A2(
        cell_2015_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2015_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2015_a_HPC2_and_U11 ( .A1(cell_2015_a_HPC2_and_a_reg[0]), .A2(
        cell_2015_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2015_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2015_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2015_a_HPC2_and_n9), 
        .ZN(cell_2015_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2015_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2015_a_HPC2_and_n9), 
        .ZN(cell_2015_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2015_a_HPC2_and_U8 ( .A(Fresh[301]), .ZN(cell_2015_a_HPC2_and_n9) );
  AND2_X1 cell_2015_a_HPC2_and_U7 ( .A1(cell_2015_and_in[1]), .A2(n466), .ZN(
        cell_2015_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2015_a_HPC2_and_U6 ( .A1(cell_2015_and_in[0]), .A2(n462), .ZN(
        cell_2015_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2015_a_HPC2_and_U5 ( .A(cell_2015_a_HPC2_and_n8), .B(
        cell_2015_a_HPC2_and_z_1__1_), .ZN(cell_2015_and_out[1]) );
  XNOR2_X1 cell_2015_a_HPC2_and_U4 ( .A(
        cell_2015_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2015_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2015_a_HPC2_and_n8) );
  XNOR2_X1 cell_2015_a_HPC2_and_U3 ( .A(cell_2015_a_HPC2_and_n7), .B(
        cell_2015_a_HPC2_and_z_0__0_), .ZN(cell_2015_and_out[0]) );
  XNOR2_X1 cell_2015_a_HPC2_and_U2 ( .A(
        cell_2015_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2015_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2015_a_HPC2_and_n7) );
  DFF_X1 cell_2015_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2015_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2015_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2015_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2015_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2015_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2015_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2015_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2015_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2015_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2016_U4 ( .A(signal_3678), .B(cell_2016_and_out[1]), .Z(
        signal_3930) );
  XOR2_X1 cell_2016_U3 ( .A(signal_2168), .B(cell_2016_and_out[0]), .Z(
        signal_2284) );
  XOR2_X1 cell_2016_U2 ( .A(signal_3678), .B(signal_3741), .Z(
        cell_2016_and_in[1]) );
  XOR2_X1 cell_2016_U1 ( .A(signal_2168), .B(signal_2231), .Z(
        cell_2016_and_in[0]) );
  XOR2_X1 cell_2016_a_HPC2_and_U14 ( .A(Fresh[302]), .B(cell_2016_and_in[0]), 
        .Z(cell_2016_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2016_a_HPC2_and_U13 ( .A(Fresh[302]), .B(cell_2016_and_in[1]), 
        .Z(cell_2016_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2016_a_HPC2_and_U12 ( .A1(cell_2016_a_HPC2_and_a_reg[1]), .A2(
        cell_2016_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2016_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2016_a_HPC2_and_U11 ( .A1(cell_2016_a_HPC2_and_a_reg[0]), .A2(
        cell_2016_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2016_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2016_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2016_a_HPC2_and_n9), 
        .ZN(cell_2016_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2016_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2016_a_HPC2_and_n9), 
        .ZN(cell_2016_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2016_a_HPC2_and_U8 ( .A(Fresh[302]), .ZN(cell_2016_a_HPC2_and_n9) );
  AND2_X1 cell_2016_a_HPC2_and_U7 ( .A1(cell_2016_and_in[1]), .A2(n466), .ZN(
        cell_2016_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2016_a_HPC2_and_U6 ( .A1(cell_2016_and_in[0]), .A2(n462), .ZN(
        cell_2016_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2016_a_HPC2_and_U5 ( .A(cell_2016_a_HPC2_and_n8), .B(
        cell_2016_a_HPC2_and_z_1__1_), .ZN(cell_2016_and_out[1]) );
  XNOR2_X1 cell_2016_a_HPC2_and_U4 ( .A(
        cell_2016_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2016_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2016_a_HPC2_and_n8) );
  XNOR2_X1 cell_2016_a_HPC2_and_U3 ( .A(cell_2016_a_HPC2_and_n7), .B(
        cell_2016_a_HPC2_and_z_0__0_), .ZN(cell_2016_and_out[0]) );
  XNOR2_X1 cell_2016_a_HPC2_and_U2 ( .A(
        cell_2016_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2016_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2016_a_HPC2_and_n7) );
  DFF_X1 cell_2016_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2016_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2016_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2016_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2016_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2016_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2016_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2016_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2016_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2016_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2017_U4 ( .A(signal_3731), .B(cell_2017_and_out[1]), .Z(
        signal_3931) );
  XOR2_X1 cell_2017_U3 ( .A(signal_2221), .B(cell_2017_and_out[0]), .Z(
        signal_2285) );
  XOR2_X1 cell_2017_U2 ( .A(signal_3731), .B(signal_3718), .Z(
        cell_2017_and_in[1]) );
  XOR2_X1 cell_2017_U1 ( .A(signal_2221), .B(signal_2208), .Z(
        cell_2017_and_in[0]) );
  XOR2_X1 cell_2017_a_HPC2_and_U14 ( .A(Fresh[303]), .B(cell_2017_and_in[0]), 
        .Z(cell_2017_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2017_a_HPC2_and_U13 ( .A(Fresh[303]), .B(cell_2017_and_in[1]), 
        .Z(cell_2017_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2017_a_HPC2_and_U12 ( .A1(cell_2017_a_HPC2_and_a_reg[1]), .A2(
        cell_2017_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2017_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2017_a_HPC2_and_U11 ( .A1(cell_2017_a_HPC2_and_a_reg[0]), .A2(
        cell_2017_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2017_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2017_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2017_a_HPC2_and_n9), 
        .ZN(cell_2017_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2017_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2017_a_HPC2_and_n9), 
        .ZN(cell_2017_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2017_a_HPC2_and_U8 ( .A(Fresh[303]), .ZN(cell_2017_a_HPC2_and_n9) );
  AND2_X1 cell_2017_a_HPC2_and_U7 ( .A1(cell_2017_and_in[1]), .A2(n466), .ZN(
        cell_2017_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2017_a_HPC2_and_U6 ( .A1(cell_2017_and_in[0]), .A2(n462), .ZN(
        cell_2017_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2017_a_HPC2_and_U5 ( .A(cell_2017_a_HPC2_and_n8), .B(
        cell_2017_a_HPC2_and_z_1__1_), .ZN(cell_2017_and_out[1]) );
  XNOR2_X1 cell_2017_a_HPC2_and_U4 ( .A(
        cell_2017_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2017_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2017_a_HPC2_and_n8) );
  XNOR2_X1 cell_2017_a_HPC2_and_U3 ( .A(cell_2017_a_HPC2_and_n7), .B(
        cell_2017_a_HPC2_and_z_0__0_), .ZN(cell_2017_and_out[0]) );
  XNOR2_X1 cell_2017_a_HPC2_and_U2 ( .A(
        cell_2017_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2017_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2017_a_HPC2_and_n7) );
  DFF_X1 cell_2017_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2017_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2017_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2017_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2017_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2017_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2017_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2017_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2017_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2017_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2018_U4 ( .A(signal_3707), .B(cell_2018_and_out[1]), .Z(
        signal_3932) );
  XOR2_X1 cell_2018_U3 ( .A(signal_2197), .B(cell_2018_and_out[0]), .Z(
        signal_2286) );
  XOR2_X1 cell_2018_U2 ( .A(signal_3707), .B(signal_3715), .Z(
        cell_2018_and_in[1]) );
  XOR2_X1 cell_2018_U1 ( .A(signal_2197), .B(signal_2205), .Z(
        cell_2018_and_in[0]) );
  XOR2_X1 cell_2018_a_HPC2_and_U14 ( .A(Fresh[304]), .B(cell_2018_and_in[0]), 
        .Z(cell_2018_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2018_a_HPC2_and_U13 ( .A(Fresh[304]), .B(cell_2018_and_in[1]), 
        .Z(cell_2018_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2018_a_HPC2_and_U12 ( .A1(cell_2018_a_HPC2_and_a_reg[1]), .A2(
        cell_2018_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2018_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2018_a_HPC2_and_U11 ( .A1(cell_2018_a_HPC2_and_a_reg[0]), .A2(
        cell_2018_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2018_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2018_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2018_a_HPC2_and_n9), 
        .ZN(cell_2018_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2018_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2018_a_HPC2_and_n9), 
        .ZN(cell_2018_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2018_a_HPC2_and_U8 ( .A(Fresh[304]), .ZN(cell_2018_a_HPC2_and_n9) );
  AND2_X1 cell_2018_a_HPC2_and_U7 ( .A1(cell_2018_and_in[1]), .A2(n466), .ZN(
        cell_2018_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2018_a_HPC2_and_U6 ( .A1(cell_2018_and_in[0]), .A2(n462), .ZN(
        cell_2018_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2018_a_HPC2_and_U5 ( .A(cell_2018_a_HPC2_and_n8), .B(
        cell_2018_a_HPC2_and_z_1__1_), .ZN(cell_2018_and_out[1]) );
  XNOR2_X1 cell_2018_a_HPC2_and_U4 ( .A(
        cell_2018_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2018_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2018_a_HPC2_and_n8) );
  XNOR2_X1 cell_2018_a_HPC2_and_U3 ( .A(cell_2018_a_HPC2_and_n7), .B(
        cell_2018_a_HPC2_and_z_0__0_), .ZN(cell_2018_and_out[0]) );
  XNOR2_X1 cell_2018_a_HPC2_and_U2 ( .A(
        cell_2018_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2018_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2018_a_HPC2_and_n7) );
  DFF_X1 cell_2018_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2018_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2018_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2018_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2018_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2018_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2018_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2018_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2018_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2018_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2019_U4 ( .A(signal_3764), .B(cell_2019_and_out[1]), .Z(
        signal_3933) );
  XOR2_X1 cell_2019_U3 ( .A(signal_2254), .B(cell_2019_and_out[0]), .Z(
        signal_2287) );
  XOR2_X1 cell_2019_U2 ( .A(signal_3764), .B(signal_3730), .Z(
        cell_2019_and_in[1]) );
  XOR2_X1 cell_2019_U1 ( .A(signal_2254), .B(signal_2220), .Z(
        cell_2019_and_in[0]) );
  XOR2_X1 cell_2019_a_HPC2_and_U14 ( .A(Fresh[305]), .B(cell_2019_and_in[0]), 
        .Z(cell_2019_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2019_a_HPC2_and_U13 ( .A(Fresh[305]), .B(cell_2019_and_in[1]), 
        .Z(cell_2019_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2019_a_HPC2_and_U12 ( .A1(cell_2019_a_HPC2_and_a_reg[1]), .A2(
        cell_2019_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2019_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2019_a_HPC2_and_U11 ( .A1(cell_2019_a_HPC2_and_a_reg[0]), .A2(
        cell_2019_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2019_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2019_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2019_a_HPC2_and_n9), 
        .ZN(cell_2019_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2019_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2019_a_HPC2_and_n9), 
        .ZN(cell_2019_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2019_a_HPC2_and_U8 ( .A(Fresh[305]), .ZN(cell_2019_a_HPC2_and_n9) );
  AND2_X1 cell_2019_a_HPC2_and_U7 ( .A1(cell_2019_and_in[1]), .A2(n466), .ZN(
        cell_2019_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2019_a_HPC2_and_U6 ( .A1(cell_2019_and_in[0]), .A2(n462), .ZN(
        cell_2019_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2019_a_HPC2_and_U5 ( .A(cell_2019_a_HPC2_and_n8), .B(
        cell_2019_a_HPC2_and_z_1__1_), .ZN(cell_2019_and_out[1]) );
  XNOR2_X1 cell_2019_a_HPC2_and_U4 ( .A(
        cell_2019_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2019_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2019_a_HPC2_and_n8) );
  XNOR2_X1 cell_2019_a_HPC2_and_U3 ( .A(cell_2019_a_HPC2_and_n7), .B(
        cell_2019_a_HPC2_and_z_0__0_), .ZN(cell_2019_and_out[0]) );
  XNOR2_X1 cell_2019_a_HPC2_and_U2 ( .A(
        cell_2019_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2019_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2019_a_HPC2_and_n7) );
  DFF_X1 cell_2019_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2019_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2019_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2019_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2019_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2019_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2019_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2019_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2019_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2019_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2020_U4 ( .A(signal_3760), .B(cell_2020_and_out[1]), .Z(
        signal_3934) );
  XOR2_X1 cell_2020_U3 ( .A(signal_2250), .B(cell_2020_and_out[0]), .Z(
        signal_2288) );
  XOR2_X1 cell_2020_U2 ( .A(signal_3760), .B(signal_3668), .Z(
        cell_2020_and_in[1]) );
  XOR2_X1 cell_2020_U1 ( .A(signal_2250), .B(signal_2158), .Z(
        cell_2020_and_in[0]) );
  XOR2_X1 cell_2020_a_HPC2_and_U14 ( .A(Fresh[306]), .B(cell_2020_and_in[0]), 
        .Z(cell_2020_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2020_a_HPC2_and_U13 ( .A(Fresh[306]), .B(cell_2020_and_in[1]), 
        .Z(cell_2020_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2020_a_HPC2_and_U12 ( .A1(cell_2020_a_HPC2_and_a_reg[1]), .A2(
        cell_2020_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2020_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2020_a_HPC2_and_U11 ( .A1(cell_2020_a_HPC2_and_a_reg[0]), .A2(
        cell_2020_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2020_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2020_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2020_a_HPC2_and_n9), 
        .ZN(cell_2020_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2020_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2020_a_HPC2_and_n9), 
        .ZN(cell_2020_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2020_a_HPC2_and_U8 ( .A(Fresh[306]), .ZN(cell_2020_a_HPC2_and_n9) );
  AND2_X1 cell_2020_a_HPC2_and_U7 ( .A1(cell_2020_and_in[1]), .A2(n467), .ZN(
        cell_2020_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2020_a_HPC2_and_U6 ( .A1(cell_2020_and_in[0]), .A2(n463), .ZN(
        cell_2020_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2020_a_HPC2_and_U5 ( .A(cell_2020_a_HPC2_and_n8), .B(
        cell_2020_a_HPC2_and_z_1__1_), .ZN(cell_2020_and_out[1]) );
  XNOR2_X1 cell_2020_a_HPC2_and_U4 ( .A(
        cell_2020_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2020_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2020_a_HPC2_and_n8) );
  XNOR2_X1 cell_2020_a_HPC2_and_U3 ( .A(cell_2020_a_HPC2_and_n7), .B(
        cell_2020_a_HPC2_and_z_0__0_), .ZN(cell_2020_and_out[0]) );
  XNOR2_X1 cell_2020_a_HPC2_and_U2 ( .A(
        cell_2020_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2020_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2020_a_HPC2_and_n7) );
  DFF_X1 cell_2020_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2020_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2020_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2020_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2020_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2020_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2020_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2020_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2020_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2020_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2021_U4 ( .A(signal_3697), .B(cell_2021_and_out[1]), .Z(
        signal_3935) );
  XOR2_X1 cell_2021_U3 ( .A(signal_2187), .B(cell_2021_and_out[0]), .Z(
        signal_2289) );
  XOR2_X1 cell_2021_U2 ( .A(signal_3697), .B(signal_3737), .Z(
        cell_2021_and_in[1]) );
  XOR2_X1 cell_2021_U1 ( .A(signal_2187), .B(signal_2227), .Z(
        cell_2021_and_in[0]) );
  XOR2_X1 cell_2021_a_HPC2_and_U14 ( .A(Fresh[307]), .B(cell_2021_and_in[0]), 
        .Z(cell_2021_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2021_a_HPC2_and_U13 ( .A(Fresh[307]), .B(cell_2021_and_in[1]), 
        .Z(cell_2021_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2021_a_HPC2_and_U12 ( .A1(cell_2021_a_HPC2_and_a_reg[1]), .A2(
        cell_2021_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2021_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2021_a_HPC2_and_U11 ( .A1(cell_2021_a_HPC2_and_a_reg[0]), .A2(
        cell_2021_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2021_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2021_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2021_a_HPC2_and_n9), 
        .ZN(cell_2021_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2021_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2021_a_HPC2_and_n9), 
        .ZN(cell_2021_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2021_a_HPC2_and_U8 ( .A(Fresh[307]), .ZN(cell_2021_a_HPC2_and_n9) );
  AND2_X1 cell_2021_a_HPC2_and_U7 ( .A1(cell_2021_and_in[1]), .A2(n467), .ZN(
        cell_2021_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2021_a_HPC2_and_U6 ( .A1(cell_2021_and_in[0]), .A2(n463), .ZN(
        cell_2021_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2021_a_HPC2_and_U5 ( .A(cell_2021_a_HPC2_and_n8), .B(
        cell_2021_a_HPC2_and_z_1__1_), .ZN(cell_2021_and_out[1]) );
  XNOR2_X1 cell_2021_a_HPC2_and_U4 ( .A(
        cell_2021_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2021_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2021_a_HPC2_and_n8) );
  XNOR2_X1 cell_2021_a_HPC2_and_U3 ( .A(cell_2021_a_HPC2_and_n7), .B(
        cell_2021_a_HPC2_and_z_0__0_), .ZN(cell_2021_and_out[0]) );
  XNOR2_X1 cell_2021_a_HPC2_and_U2 ( .A(
        cell_2021_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2021_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2021_a_HPC2_and_n7) );
  DFF_X1 cell_2021_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2021_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2021_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2021_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2021_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2021_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2021_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2021_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2021_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2021_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2022_U4 ( .A(signal_3726), .B(cell_2022_and_out[1]), .Z(
        signal_3936) );
  XOR2_X1 cell_2022_U3 ( .A(signal_2216), .B(cell_2022_and_out[0]), .Z(
        signal_2290) );
  XOR2_X1 cell_2022_U2 ( .A(signal_3726), .B(signal_3535), .Z(
        cell_2022_and_in[1]) );
  XOR2_X1 cell_2022_U1 ( .A(signal_2216), .B(signal_2097), .Z(
        cell_2022_and_in[0]) );
  XOR2_X1 cell_2022_a_HPC2_and_U14 ( .A(Fresh[308]), .B(cell_2022_and_in[0]), 
        .Z(cell_2022_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2022_a_HPC2_and_U13 ( .A(Fresh[308]), .B(cell_2022_and_in[1]), 
        .Z(cell_2022_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2022_a_HPC2_and_U12 ( .A1(cell_2022_a_HPC2_and_a_reg[1]), .A2(
        cell_2022_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2022_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2022_a_HPC2_and_U11 ( .A1(cell_2022_a_HPC2_and_a_reg[0]), .A2(
        cell_2022_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2022_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2022_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2022_a_HPC2_and_n9), 
        .ZN(cell_2022_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2022_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2022_a_HPC2_and_n9), 
        .ZN(cell_2022_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2022_a_HPC2_and_U8 ( .A(Fresh[308]), .ZN(cell_2022_a_HPC2_and_n9) );
  AND2_X1 cell_2022_a_HPC2_and_U7 ( .A1(cell_2022_and_in[1]), .A2(n467), .ZN(
        cell_2022_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2022_a_HPC2_and_U6 ( .A1(cell_2022_and_in[0]), .A2(n463), .ZN(
        cell_2022_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2022_a_HPC2_and_U5 ( .A(cell_2022_a_HPC2_and_n8), .B(
        cell_2022_a_HPC2_and_z_1__1_), .ZN(cell_2022_and_out[1]) );
  XNOR2_X1 cell_2022_a_HPC2_and_U4 ( .A(
        cell_2022_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2022_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2022_a_HPC2_and_n8) );
  XNOR2_X1 cell_2022_a_HPC2_and_U3 ( .A(cell_2022_a_HPC2_and_n7), .B(
        cell_2022_a_HPC2_and_z_0__0_), .ZN(cell_2022_and_out[0]) );
  XNOR2_X1 cell_2022_a_HPC2_and_U2 ( .A(
        cell_2022_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2022_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2022_a_HPC2_and_n7) );
  DFF_X1 cell_2022_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2022_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2022_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2022_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2022_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2022_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2022_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2022_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2022_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2022_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2023_U4 ( .A(signal_3759), .B(cell_2023_and_out[1]), .Z(
        signal_3937) );
  XOR2_X1 cell_2023_U3 ( .A(signal_2249), .B(cell_2023_and_out[0]), .Z(
        signal_2291) );
  XOR2_X1 cell_2023_U2 ( .A(signal_3759), .B(signal_3674), .Z(
        cell_2023_and_in[1]) );
  XOR2_X1 cell_2023_U1 ( .A(signal_2249), .B(signal_2164), .Z(
        cell_2023_and_in[0]) );
  XOR2_X1 cell_2023_a_HPC2_and_U14 ( .A(Fresh[309]), .B(cell_2023_and_in[0]), 
        .Z(cell_2023_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2023_a_HPC2_and_U13 ( .A(Fresh[309]), .B(cell_2023_and_in[1]), 
        .Z(cell_2023_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2023_a_HPC2_and_U12 ( .A1(cell_2023_a_HPC2_and_a_reg[1]), .A2(
        cell_2023_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2023_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2023_a_HPC2_and_U11 ( .A1(cell_2023_a_HPC2_and_a_reg[0]), .A2(
        cell_2023_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2023_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2023_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2023_a_HPC2_and_n9), 
        .ZN(cell_2023_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2023_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2023_a_HPC2_and_n9), 
        .ZN(cell_2023_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2023_a_HPC2_and_U8 ( .A(Fresh[309]), .ZN(cell_2023_a_HPC2_and_n9) );
  AND2_X1 cell_2023_a_HPC2_and_U7 ( .A1(cell_2023_and_in[1]), .A2(n467), .ZN(
        cell_2023_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2023_a_HPC2_and_U6 ( .A1(cell_2023_and_in[0]), .A2(n463), .ZN(
        cell_2023_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2023_a_HPC2_and_U5 ( .A(cell_2023_a_HPC2_and_n8), .B(
        cell_2023_a_HPC2_and_z_1__1_), .ZN(cell_2023_and_out[1]) );
  XNOR2_X1 cell_2023_a_HPC2_and_U4 ( .A(
        cell_2023_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2023_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2023_a_HPC2_and_n8) );
  XNOR2_X1 cell_2023_a_HPC2_and_U3 ( .A(cell_2023_a_HPC2_and_n7), .B(
        cell_2023_a_HPC2_and_z_0__0_), .ZN(cell_2023_and_out[0]) );
  XNOR2_X1 cell_2023_a_HPC2_and_U2 ( .A(
        cell_2023_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2023_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2023_a_HPC2_and_n7) );
  DFF_X1 cell_2023_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2023_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2023_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2023_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2023_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2023_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2023_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2023_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2023_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2023_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2024_U4 ( .A(signal_3501), .B(cell_2024_and_out[1]), .Z(
        signal_3938) );
  XOR2_X1 cell_2024_U3 ( .A(signal_2063), .B(cell_2024_and_out[0]), .Z(
        signal_2292) );
  XOR2_X1 cell_2024_U2 ( .A(signal_3501), .B(signal_3729), .Z(
        cell_2024_and_in[1]) );
  XOR2_X1 cell_2024_U1 ( .A(signal_2063), .B(signal_2219), .Z(
        cell_2024_and_in[0]) );
  XOR2_X1 cell_2024_a_HPC2_and_U14 ( .A(Fresh[310]), .B(cell_2024_and_in[0]), 
        .Z(cell_2024_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2024_a_HPC2_and_U13 ( .A(Fresh[310]), .B(cell_2024_and_in[1]), 
        .Z(cell_2024_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2024_a_HPC2_and_U12 ( .A1(cell_2024_a_HPC2_and_a_reg[1]), .A2(
        cell_2024_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2024_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2024_a_HPC2_and_U11 ( .A1(cell_2024_a_HPC2_and_a_reg[0]), .A2(
        cell_2024_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2024_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2024_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2024_a_HPC2_and_n9), 
        .ZN(cell_2024_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2024_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2024_a_HPC2_and_n9), 
        .ZN(cell_2024_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2024_a_HPC2_and_U8 ( .A(Fresh[310]), .ZN(cell_2024_a_HPC2_and_n9) );
  AND2_X1 cell_2024_a_HPC2_and_U7 ( .A1(cell_2024_and_in[1]), .A2(n467), .ZN(
        cell_2024_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2024_a_HPC2_and_U6 ( .A1(cell_2024_and_in[0]), .A2(n463), .ZN(
        cell_2024_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2024_a_HPC2_and_U5 ( .A(cell_2024_a_HPC2_and_n8), .B(
        cell_2024_a_HPC2_and_z_1__1_), .ZN(cell_2024_and_out[1]) );
  XNOR2_X1 cell_2024_a_HPC2_and_U4 ( .A(
        cell_2024_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2024_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2024_a_HPC2_and_n8) );
  XNOR2_X1 cell_2024_a_HPC2_and_U3 ( .A(cell_2024_a_HPC2_and_n7), .B(
        cell_2024_a_HPC2_and_z_0__0_), .ZN(cell_2024_and_out[0]) );
  XNOR2_X1 cell_2024_a_HPC2_and_U2 ( .A(
        cell_2024_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2024_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2024_a_HPC2_and_n7) );
  DFF_X1 cell_2024_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2024_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2024_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2024_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2024_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2024_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2024_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2024_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2024_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2024_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2025_U4 ( .A(signal_3770), .B(cell_2025_and_out[1]), .Z(
        signal_3939) );
  XOR2_X1 cell_2025_U3 ( .A(signal_2260), .B(cell_2025_and_out[0]), .Z(
        signal_2293) );
  XOR2_X1 cell_2025_U2 ( .A(signal_3770), .B(signal_3785), .Z(
        cell_2025_and_in[1]) );
  XOR2_X1 cell_2025_U1 ( .A(signal_2260), .B(signal_2275), .Z(
        cell_2025_and_in[0]) );
  XOR2_X1 cell_2025_a_HPC2_and_U14 ( .A(Fresh[311]), .B(cell_2025_and_in[0]), 
        .Z(cell_2025_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2025_a_HPC2_and_U13 ( .A(Fresh[311]), .B(cell_2025_and_in[1]), 
        .Z(cell_2025_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2025_a_HPC2_and_U12 ( .A1(cell_2025_a_HPC2_and_a_reg[1]), .A2(
        cell_2025_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2025_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2025_a_HPC2_and_U11 ( .A1(cell_2025_a_HPC2_and_a_reg[0]), .A2(
        cell_2025_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2025_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2025_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2025_a_HPC2_and_n9), 
        .ZN(cell_2025_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2025_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2025_a_HPC2_and_n9), 
        .ZN(cell_2025_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2025_a_HPC2_and_U8 ( .A(Fresh[311]), .ZN(cell_2025_a_HPC2_and_n9) );
  AND2_X1 cell_2025_a_HPC2_and_U7 ( .A1(cell_2025_and_in[1]), .A2(n467), .ZN(
        cell_2025_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2025_a_HPC2_and_U6 ( .A1(cell_2025_and_in[0]), .A2(n463), .ZN(
        cell_2025_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2025_a_HPC2_and_U5 ( .A(cell_2025_a_HPC2_and_n8), .B(
        cell_2025_a_HPC2_and_z_1__1_), .ZN(cell_2025_and_out[1]) );
  XNOR2_X1 cell_2025_a_HPC2_and_U4 ( .A(
        cell_2025_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2025_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2025_a_HPC2_and_n8) );
  XNOR2_X1 cell_2025_a_HPC2_and_U3 ( .A(cell_2025_a_HPC2_and_n7), .B(
        cell_2025_a_HPC2_and_z_0__0_), .ZN(cell_2025_and_out[0]) );
  XNOR2_X1 cell_2025_a_HPC2_and_U2 ( .A(
        cell_2025_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2025_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2025_a_HPC2_and_n7) );
  DFF_X1 cell_2025_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2025_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2025_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2025_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2025_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2025_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2025_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2025_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2025_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2025_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2026_U4 ( .A(signal_3677), .B(cell_2026_and_out[1]), .Z(
        signal_3940) );
  XOR2_X1 cell_2026_U3 ( .A(signal_2167), .B(cell_2026_and_out[0]), .Z(
        signal_2294) );
  XOR2_X1 cell_2026_U2 ( .A(signal_3677), .B(signal_3691), .Z(
        cell_2026_and_in[1]) );
  XOR2_X1 cell_2026_U1 ( .A(signal_2167), .B(signal_2181), .Z(
        cell_2026_and_in[0]) );
  XOR2_X1 cell_2026_a_HPC2_and_U14 ( .A(Fresh[312]), .B(cell_2026_and_in[0]), 
        .Z(cell_2026_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2026_a_HPC2_and_U13 ( .A(Fresh[312]), .B(cell_2026_and_in[1]), 
        .Z(cell_2026_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2026_a_HPC2_and_U12 ( .A1(cell_2026_a_HPC2_and_a_reg[1]), .A2(
        cell_2026_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2026_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2026_a_HPC2_and_U11 ( .A1(cell_2026_a_HPC2_and_a_reg[0]), .A2(
        cell_2026_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2026_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2026_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2026_a_HPC2_and_n9), 
        .ZN(cell_2026_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2026_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2026_a_HPC2_and_n9), 
        .ZN(cell_2026_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2026_a_HPC2_and_U8 ( .A(Fresh[312]), .ZN(cell_2026_a_HPC2_and_n9) );
  AND2_X1 cell_2026_a_HPC2_and_U7 ( .A1(cell_2026_and_in[1]), .A2(n467), .ZN(
        cell_2026_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2026_a_HPC2_and_U6 ( .A1(cell_2026_and_in[0]), .A2(n463), .ZN(
        cell_2026_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2026_a_HPC2_and_U5 ( .A(cell_2026_a_HPC2_and_n8), .B(
        cell_2026_a_HPC2_and_z_1__1_), .ZN(cell_2026_and_out[1]) );
  XNOR2_X1 cell_2026_a_HPC2_and_U4 ( .A(
        cell_2026_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2026_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2026_a_HPC2_and_n8) );
  XNOR2_X1 cell_2026_a_HPC2_and_U3 ( .A(cell_2026_a_HPC2_and_n7), .B(
        cell_2026_a_HPC2_and_z_0__0_), .ZN(cell_2026_and_out[0]) );
  XNOR2_X1 cell_2026_a_HPC2_and_U2 ( .A(
        cell_2026_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2026_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2026_a_HPC2_and_n7) );
  DFF_X1 cell_2026_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2026_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2026_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2026_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2026_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2026_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2026_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2026_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2026_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2026_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2027_U4 ( .A(signal_3708), .B(cell_2027_and_out[1]), .Z(
        signal_3941) );
  XOR2_X1 cell_2027_U3 ( .A(signal_2198), .B(cell_2027_and_out[0]), .Z(
        signal_2295) );
  XOR2_X1 cell_2027_U2 ( .A(signal_3708), .B(signal_3471), .Z(
        cell_2027_and_in[1]) );
  XOR2_X1 cell_2027_U1 ( .A(signal_2198), .B(signal_2033), .Z(
        cell_2027_and_in[0]) );
  XOR2_X1 cell_2027_a_HPC2_and_U14 ( .A(Fresh[313]), .B(cell_2027_and_in[0]), 
        .Z(cell_2027_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2027_a_HPC2_and_U13 ( .A(Fresh[313]), .B(cell_2027_and_in[1]), 
        .Z(cell_2027_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2027_a_HPC2_and_U12 ( .A1(cell_2027_a_HPC2_and_a_reg[1]), .A2(
        cell_2027_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2027_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2027_a_HPC2_and_U11 ( .A1(cell_2027_a_HPC2_and_a_reg[0]), .A2(
        cell_2027_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2027_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2027_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2027_a_HPC2_and_n9), 
        .ZN(cell_2027_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2027_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2027_a_HPC2_and_n9), 
        .ZN(cell_2027_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2027_a_HPC2_and_U8 ( .A(Fresh[313]), .ZN(cell_2027_a_HPC2_and_n9) );
  AND2_X1 cell_2027_a_HPC2_and_U7 ( .A1(cell_2027_and_in[1]), .A2(n467), .ZN(
        cell_2027_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2027_a_HPC2_and_U6 ( .A1(cell_2027_and_in[0]), .A2(n463), .ZN(
        cell_2027_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2027_a_HPC2_and_U5 ( .A(cell_2027_a_HPC2_and_n8), .B(
        cell_2027_a_HPC2_and_z_1__1_), .ZN(cell_2027_and_out[1]) );
  XNOR2_X1 cell_2027_a_HPC2_and_U4 ( .A(
        cell_2027_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2027_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2027_a_HPC2_and_n8) );
  XNOR2_X1 cell_2027_a_HPC2_and_U3 ( .A(cell_2027_a_HPC2_and_n7), .B(
        cell_2027_a_HPC2_and_z_0__0_), .ZN(cell_2027_and_out[0]) );
  XNOR2_X1 cell_2027_a_HPC2_and_U2 ( .A(
        cell_2027_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2027_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2027_a_HPC2_and_n7) );
  DFF_X1 cell_2027_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2027_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2027_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2027_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2027_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2027_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2027_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2027_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2027_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2027_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2028_U4 ( .A(signal_3753), .B(cell_2028_and_out[1]), .Z(
        signal_3942) );
  XOR2_X1 cell_2028_U3 ( .A(signal_2243), .B(cell_2028_and_out[0]), .Z(
        signal_2296) );
  XOR2_X1 cell_2028_U2 ( .A(signal_3753), .B(signal_3725), .Z(
        cell_2028_and_in[1]) );
  XOR2_X1 cell_2028_U1 ( .A(signal_2243), .B(signal_2215), .Z(
        cell_2028_and_in[0]) );
  XOR2_X1 cell_2028_a_HPC2_and_U14 ( .A(Fresh[314]), .B(cell_2028_and_in[0]), 
        .Z(cell_2028_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2028_a_HPC2_and_U13 ( .A(Fresh[314]), .B(cell_2028_and_in[1]), 
        .Z(cell_2028_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2028_a_HPC2_and_U12 ( .A1(cell_2028_a_HPC2_and_a_reg[1]), .A2(
        cell_2028_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2028_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2028_a_HPC2_and_U11 ( .A1(cell_2028_a_HPC2_and_a_reg[0]), .A2(
        cell_2028_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2028_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2028_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2028_a_HPC2_and_n9), 
        .ZN(cell_2028_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2028_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2028_a_HPC2_and_n9), 
        .ZN(cell_2028_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2028_a_HPC2_and_U8 ( .A(Fresh[314]), .ZN(cell_2028_a_HPC2_and_n9) );
  AND2_X1 cell_2028_a_HPC2_and_U7 ( .A1(cell_2028_and_in[1]), .A2(n467), .ZN(
        cell_2028_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2028_a_HPC2_and_U6 ( .A1(cell_2028_and_in[0]), .A2(n463), .ZN(
        cell_2028_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2028_a_HPC2_and_U5 ( .A(cell_2028_a_HPC2_and_n8), .B(
        cell_2028_a_HPC2_and_z_1__1_), .ZN(cell_2028_and_out[1]) );
  XNOR2_X1 cell_2028_a_HPC2_and_U4 ( .A(
        cell_2028_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2028_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2028_a_HPC2_and_n8) );
  XNOR2_X1 cell_2028_a_HPC2_and_U3 ( .A(cell_2028_a_HPC2_and_n7), .B(
        cell_2028_a_HPC2_and_z_0__0_), .ZN(cell_2028_and_out[0]) );
  XNOR2_X1 cell_2028_a_HPC2_and_U2 ( .A(
        cell_2028_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2028_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2028_a_HPC2_and_n7) );
  DFF_X1 cell_2028_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2028_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2028_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2028_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2028_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2028_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2028_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2028_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2028_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2028_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2029_U4 ( .A(signal_3781), .B(cell_2029_and_out[1]), .Z(
        signal_3943) );
  XOR2_X1 cell_2029_U3 ( .A(signal_2271), .B(cell_2029_and_out[0]), .Z(
        signal_2297) );
  XOR2_X1 cell_2029_U2 ( .A(signal_3781), .B(signal_3669), .Z(
        cell_2029_and_in[1]) );
  XOR2_X1 cell_2029_U1 ( .A(signal_2271), .B(signal_2159), .Z(
        cell_2029_and_in[0]) );
  XOR2_X1 cell_2029_a_HPC2_and_U14 ( .A(Fresh[315]), .B(cell_2029_and_in[0]), 
        .Z(cell_2029_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2029_a_HPC2_and_U13 ( .A(Fresh[315]), .B(cell_2029_and_in[1]), 
        .Z(cell_2029_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2029_a_HPC2_and_U12 ( .A1(cell_2029_a_HPC2_and_a_reg[1]), .A2(
        cell_2029_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2029_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2029_a_HPC2_and_U11 ( .A1(cell_2029_a_HPC2_and_a_reg[0]), .A2(
        cell_2029_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2029_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2029_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2029_a_HPC2_and_n9), 
        .ZN(cell_2029_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2029_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2029_a_HPC2_and_n9), 
        .ZN(cell_2029_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2029_a_HPC2_and_U8 ( .A(Fresh[315]), .ZN(cell_2029_a_HPC2_and_n9) );
  AND2_X1 cell_2029_a_HPC2_and_U7 ( .A1(cell_2029_and_in[1]), .A2(n467), .ZN(
        cell_2029_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2029_a_HPC2_and_U6 ( .A1(cell_2029_and_in[0]), .A2(n463), .ZN(
        cell_2029_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2029_a_HPC2_and_U5 ( .A(cell_2029_a_HPC2_and_n8), .B(
        cell_2029_a_HPC2_and_z_1__1_), .ZN(cell_2029_and_out[1]) );
  XNOR2_X1 cell_2029_a_HPC2_and_U4 ( .A(
        cell_2029_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2029_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2029_a_HPC2_and_n8) );
  XNOR2_X1 cell_2029_a_HPC2_and_U3 ( .A(cell_2029_a_HPC2_and_n7), .B(
        cell_2029_a_HPC2_and_z_0__0_), .ZN(cell_2029_and_out[0]) );
  XNOR2_X1 cell_2029_a_HPC2_and_U2 ( .A(
        cell_2029_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2029_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2029_a_HPC2_and_n7) );
  DFF_X1 cell_2029_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2029_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2029_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2029_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2029_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2029_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2029_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2029_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2029_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2029_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2030_U4 ( .A(signal_3755), .B(cell_2030_and_out[1]), .Z(
        signal_3944) );
  XOR2_X1 cell_2030_U3 ( .A(signal_2245), .B(cell_2030_and_out[0]), .Z(
        signal_2298) );
  XOR2_X1 cell_2030_U2 ( .A(signal_3755), .B(signal_3710), .Z(
        cell_2030_and_in[1]) );
  XOR2_X1 cell_2030_U1 ( .A(signal_2245), .B(signal_2200), .Z(
        cell_2030_and_in[0]) );
  XOR2_X1 cell_2030_a_HPC2_and_U14 ( .A(Fresh[316]), .B(cell_2030_and_in[0]), 
        .Z(cell_2030_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2030_a_HPC2_and_U13 ( .A(Fresh[316]), .B(cell_2030_and_in[1]), 
        .Z(cell_2030_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2030_a_HPC2_and_U12 ( .A1(cell_2030_a_HPC2_and_a_reg[1]), .A2(
        cell_2030_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2030_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2030_a_HPC2_and_U11 ( .A1(cell_2030_a_HPC2_and_a_reg[0]), .A2(
        cell_2030_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2030_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2030_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2030_a_HPC2_and_n9), 
        .ZN(cell_2030_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2030_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2030_a_HPC2_and_n9), 
        .ZN(cell_2030_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2030_a_HPC2_and_U8 ( .A(Fresh[316]), .ZN(cell_2030_a_HPC2_and_n9) );
  AND2_X1 cell_2030_a_HPC2_and_U7 ( .A1(cell_2030_and_in[1]), .A2(n467), .ZN(
        cell_2030_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2030_a_HPC2_and_U6 ( .A1(cell_2030_and_in[0]), .A2(n463), .ZN(
        cell_2030_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2030_a_HPC2_and_U5 ( .A(cell_2030_a_HPC2_and_n8), .B(
        cell_2030_a_HPC2_and_z_1__1_), .ZN(cell_2030_and_out[1]) );
  XNOR2_X1 cell_2030_a_HPC2_and_U4 ( .A(
        cell_2030_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2030_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2030_a_HPC2_and_n8) );
  XNOR2_X1 cell_2030_a_HPC2_and_U3 ( .A(cell_2030_a_HPC2_and_n7), .B(
        cell_2030_a_HPC2_and_z_0__0_), .ZN(cell_2030_and_out[0]) );
  XNOR2_X1 cell_2030_a_HPC2_and_U2 ( .A(
        cell_2030_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2030_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2030_a_HPC2_and_n7) );
  DFF_X1 cell_2030_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2030_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2030_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2030_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2030_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2030_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2030_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2030_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2030_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2030_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2031_U4 ( .A(signal_3681), .B(cell_2031_and_out[1]), .Z(
        signal_3945) );
  XOR2_X1 cell_2031_U3 ( .A(signal_2171), .B(cell_2031_and_out[0]), .Z(
        signal_2299) );
  XOR2_X1 cell_2031_U2 ( .A(signal_3681), .B(signal_3784), .Z(
        cell_2031_and_in[1]) );
  XOR2_X1 cell_2031_U1 ( .A(signal_2171), .B(signal_2274), .Z(
        cell_2031_and_in[0]) );
  XOR2_X1 cell_2031_a_HPC2_and_U14 ( .A(Fresh[317]), .B(cell_2031_and_in[0]), 
        .Z(cell_2031_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2031_a_HPC2_and_U13 ( .A(Fresh[317]), .B(cell_2031_and_in[1]), 
        .Z(cell_2031_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2031_a_HPC2_and_U12 ( .A1(cell_2031_a_HPC2_and_a_reg[1]), .A2(
        cell_2031_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2031_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2031_a_HPC2_and_U11 ( .A1(cell_2031_a_HPC2_and_a_reg[0]), .A2(
        cell_2031_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2031_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2031_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2031_a_HPC2_and_n9), 
        .ZN(cell_2031_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2031_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2031_a_HPC2_and_n9), 
        .ZN(cell_2031_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2031_a_HPC2_and_U8 ( .A(Fresh[317]), .ZN(cell_2031_a_HPC2_and_n9) );
  AND2_X1 cell_2031_a_HPC2_and_U7 ( .A1(cell_2031_and_in[1]), .A2(n467), .ZN(
        cell_2031_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2031_a_HPC2_and_U6 ( .A1(cell_2031_and_in[0]), .A2(n463), .ZN(
        cell_2031_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2031_a_HPC2_and_U5 ( .A(cell_2031_a_HPC2_and_n8), .B(
        cell_2031_a_HPC2_and_z_1__1_), .ZN(cell_2031_and_out[1]) );
  XNOR2_X1 cell_2031_a_HPC2_and_U4 ( .A(
        cell_2031_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2031_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2031_a_HPC2_and_n8) );
  XNOR2_X1 cell_2031_a_HPC2_and_U3 ( .A(cell_2031_a_HPC2_and_n7), .B(
        cell_2031_a_HPC2_and_z_0__0_), .ZN(cell_2031_and_out[0]) );
  XNOR2_X1 cell_2031_a_HPC2_and_U2 ( .A(
        cell_2031_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2031_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2031_a_HPC2_and_n7) );
  DFF_X1 cell_2031_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2031_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2031_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2031_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2031_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2031_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2031_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2031_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2031_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2031_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2032_U4 ( .A(signal_3699), .B(cell_2032_and_out[1]), .Z(
        signal_3946) );
  XOR2_X1 cell_2032_U3 ( .A(signal_2189), .B(cell_2032_and_out[0]), .Z(
        signal_2300) );
  XOR2_X1 cell_2032_U2 ( .A(signal_3699), .B(signal_3703), .Z(
        cell_2032_and_in[1]) );
  XOR2_X1 cell_2032_U1 ( .A(signal_2189), .B(signal_2193), .Z(
        cell_2032_and_in[0]) );
  XOR2_X1 cell_2032_a_HPC2_and_U14 ( .A(Fresh[318]), .B(cell_2032_and_in[0]), 
        .Z(cell_2032_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2032_a_HPC2_and_U13 ( .A(Fresh[318]), .B(cell_2032_and_in[1]), 
        .Z(cell_2032_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2032_a_HPC2_and_U12 ( .A1(cell_2032_a_HPC2_and_a_reg[1]), .A2(
        cell_2032_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2032_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2032_a_HPC2_and_U11 ( .A1(cell_2032_a_HPC2_and_a_reg[0]), .A2(
        cell_2032_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2032_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2032_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2032_a_HPC2_and_n9), 
        .ZN(cell_2032_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2032_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2032_a_HPC2_and_n9), 
        .ZN(cell_2032_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2032_a_HPC2_and_U8 ( .A(Fresh[318]), .ZN(cell_2032_a_HPC2_and_n9) );
  AND2_X1 cell_2032_a_HPC2_and_U7 ( .A1(cell_2032_and_in[1]), .A2(n469), .ZN(
        cell_2032_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2032_a_HPC2_and_U6 ( .A1(cell_2032_and_in[0]), .A2(n465), .ZN(
        cell_2032_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2032_a_HPC2_and_U5 ( .A(cell_2032_a_HPC2_and_n8), .B(
        cell_2032_a_HPC2_and_z_1__1_), .ZN(cell_2032_and_out[1]) );
  XNOR2_X1 cell_2032_a_HPC2_and_U4 ( .A(
        cell_2032_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2032_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2032_a_HPC2_and_n8) );
  XNOR2_X1 cell_2032_a_HPC2_and_U3 ( .A(cell_2032_a_HPC2_and_n7), .B(
        cell_2032_a_HPC2_and_z_0__0_), .ZN(cell_2032_and_out[0]) );
  XNOR2_X1 cell_2032_a_HPC2_and_U2 ( .A(
        cell_2032_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2032_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2032_a_HPC2_and_n7) );
  DFF_X1 cell_2032_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2032_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2032_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2032_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2032_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2032_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2032_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2032_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2032_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2032_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2033_U4 ( .A(signal_3717), .B(cell_2033_and_out[1]), .Z(
        signal_3947) );
  XOR2_X1 cell_2033_U3 ( .A(signal_2207), .B(cell_2033_and_out[0]), .Z(
        signal_2301) );
  XOR2_X1 cell_2033_U2 ( .A(signal_3717), .B(signal_3772), .Z(
        cell_2033_and_in[1]) );
  XOR2_X1 cell_2033_U1 ( .A(signal_2207), .B(signal_2262), .Z(
        cell_2033_and_in[0]) );
  XOR2_X1 cell_2033_a_HPC2_and_U14 ( .A(Fresh[319]), .B(cell_2033_and_in[0]), 
        .Z(cell_2033_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2033_a_HPC2_and_U13 ( .A(Fresh[319]), .B(cell_2033_and_in[1]), 
        .Z(cell_2033_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2033_a_HPC2_and_U12 ( .A1(cell_2033_a_HPC2_and_a_reg[1]), .A2(
        cell_2033_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2033_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2033_a_HPC2_and_U11 ( .A1(cell_2033_a_HPC2_and_a_reg[0]), .A2(
        cell_2033_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2033_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2033_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2033_a_HPC2_and_n9), 
        .ZN(cell_2033_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2033_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2033_a_HPC2_and_n9), 
        .ZN(cell_2033_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2033_a_HPC2_and_U8 ( .A(Fresh[319]), .ZN(cell_2033_a_HPC2_and_n9) );
  AND2_X1 cell_2033_a_HPC2_and_U7 ( .A1(cell_2033_and_in[1]), .A2(n466), .ZN(
        cell_2033_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2033_a_HPC2_and_U6 ( .A1(cell_2033_and_in[0]), .A2(n462), .ZN(
        cell_2033_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2033_a_HPC2_and_U5 ( .A(cell_2033_a_HPC2_and_n8), .B(
        cell_2033_a_HPC2_and_z_1__1_), .ZN(cell_2033_and_out[1]) );
  XNOR2_X1 cell_2033_a_HPC2_and_U4 ( .A(
        cell_2033_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2033_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2033_a_HPC2_and_n8) );
  XNOR2_X1 cell_2033_a_HPC2_and_U3 ( .A(cell_2033_a_HPC2_and_n7), .B(
        cell_2033_a_HPC2_and_z_0__0_), .ZN(cell_2033_and_out[0]) );
  XNOR2_X1 cell_2033_a_HPC2_and_U2 ( .A(
        cell_2033_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2033_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2033_a_HPC2_and_n7) );
  DFF_X1 cell_2033_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2033_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2033_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2033_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2033_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2033_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2033_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2033_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2033_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2033_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2034_U4 ( .A(signal_3778), .B(cell_2034_and_out[1]), .Z(
        signal_3948) );
  XOR2_X1 cell_2034_U3 ( .A(signal_2268), .B(cell_2034_and_out[0]), .Z(
        signal_2302) );
  XOR2_X1 cell_2034_U2 ( .A(signal_3778), .B(signal_3727), .Z(
        cell_2034_and_in[1]) );
  XOR2_X1 cell_2034_U1 ( .A(signal_2268), .B(signal_2217), .Z(
        cell_2034_and_in[0]) );
  XOR2_X1 cell_2034_a_HPC2_and_U14 ( .A(Fresh[320]), .B(cell_2034_and_in[0]), 
        .Z(cell_2034_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2034_a_HPC2_and_U13 ( .A(Fresh[320]), .B(cell_2034_and_in[1]), 
        .Z(cell_2034_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2034_a_HPC2_and_U12 ( .A1(cell_2034_a_HPC2_and_a_reg[1]), .A2(
        cell_2034_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2034_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2034_a_HPC2_and_U11 ( .A1(cell_2034_a_HPC2_and_a_reg[0]), .A2(
        cell_2034_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2034_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2034_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2034_a_HPC2_and_n9), 
        .ZN(cell_2034_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2034_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2034_a_HPC2_and_n9), 
        .ZN(cell_2034_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2034_a_HPC2_and_U8 ( .A(Fresh[320]), .ZN(cell_2034_a_HPC2_and_n9) );
  AND2_X1 cell_2034_a_HPC2_and_U7 ( .A1(cell_2034_and_in[1]), .A2(n467), .ZN(
        cell_2034_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2034_a_HPC2_and_U6 ( .A1(cell_2034_and_in[0]), .A2(n463), .ZN(
        cell_2034_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2034_a_HPC2_and_U5 ( .A(cell_2034_a_HPC2_and_n8), .B(
        cell_2034_a_HPC2_and_z_1__1_), .ZN(cell_2034_and_out[1]) );
  XNOR2_X1 cell_2034_a_HPC2_and_U4 ( .A(
        cell_2034_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2034_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2034_a_HPC2_and_n8) );
  XNOR2_X1 cell_2034_a_HPC2_and_U3 ( .A(cell_2034_a_HPC2_and_n7), .B(
        cell_2034_a_HPC2_and_z_0__0_), .ZN(cell_2034_and_out[0]) );
  XNOR2_X1 cell_2034_a_HPC2_and_U2 ( .A(
        cell_2034_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2034_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2034_a_HPC2_and_n7) );
  DFF_X1 cell_2034_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2034_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2034_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2034_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2034_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2034_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2034_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2034_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2034_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2034_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2035_U4 ( .A(signal_3766), .B(cell_2035_and_out[1]), .Z(
        signal_3949) );
  XOR2_X1 cell_2035_U3 ( .A(signal_2256), .B(cell_2035_and_out[0]), .Z(
        signal_2303) );
  XOR2_X1 cell_2035_U2 ( .A(signal_3766), .B(signal_3705), .Z(
        cell_2035_and_in[1]) );
  XOR2_X1 cell_2035_U1 ( .A(signal_2256), .B(signal_2195), .Z(
        cell_2035_and_in[0]) );
  XOR2_X1 cell_2035_a_HPC2_and_U14 ( .A(Fresh[321]), .B(cell_2035_and_in[0]), 
        .Z(cell_2035_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2035_a_HPC2_and_U13 ( .A(Fresh[321]), .B(cell_2035_and_in[1]), 
        .Z(cell_2035_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2035_a_HPC2_and_U12 ( .A1(cell_2035_a_HPC2_and_a_reg[1]), .A2(
        cell_2035_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2035_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2035_a_HPC2_and_U11 ( .A1(cell_2035_a_HPC2_and_a_reg[0]), .A2(
        cell_2035_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2035_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2035_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2035_a_HPC2_and_n9), 
        .ZN(cell_2035_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2035_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2035_a_HPC2_and_n9), 
        .ZN(cell_2035_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2035_a_HPC2_and_U8 ( .A(Fresh[321]), .ZN(cell_2035_a_HPC2_and_n9) );
  AND2_X1 cell_2035_a_HPC2_and_U7 ( .A1(cell_2035_and_in[1]), .A2(n468), .ZN(
        cell_2035_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2035_a_HPC2_and_U6 ( .A1(cell_2035_and_in[0]), .A2(n464), .ZN(
        cell_2035_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2035_a_HPC2_and_U5 ( .A(cell_2035_a_HPC2_and_n8), .B(
        cell_2035_a_HPC2_and_z_1__1_), .ZN(cell_2035_and_out[1]) );
  XNOR2_X1 cell_2035_a_HPC2_and_U4 ( .A(
        cell_2035_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2035_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2035_a_HPC2_and_n8) );
  XNOR2_X1 cell_2035_a_HPC2_and_U3 ( .A(cell_2035_a_HPC2_and_n7), .B(
        cell_2035_a_HPC2_and_z_0__0_), .ZN(cell_2035_and_out[0]) );
  XNOR2_X1 cell_2035_a_HPC2_and_U2 ( .A(
        cell_2035_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2035_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2035_a_HPC2_and_n7) );
  DFF_X1 cell_2035_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2035_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2035_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2035_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2035_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2035_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2035_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2035_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2035_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2035_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2036_U4 ( .A(signal_3775), .B(cell_2036_and_out[1]), .Z(
        signal_3950) );
  XOR2_X1 cell_2036_U3 ( .A(signal_2265), .B(cell_2036_and_out[0]), .Z(
        signal_2304) );
  XOR2_X1 cell_2036_U2 ( .A(signal_3775), .B(signal_3771), .Z(
        cell_2036_and_in[1]) );
  XOR2_X1 cell_2036_U1 ( .A(signal_2265), .B(signal_2261), .Z(
        cell_2036_and_in[0]) );
  XOR2_X1 cell_2036_a_HPC2_and_U14 ( .A(Fresh[322]), .B(cell_2036_and_in[0]), 
        .Z(cell_2036_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2036_a_HPC2_and_U13 ( .A(Fresh[322]), .B(cell_2036_and_in[1]), 
        .Z(cell_2036_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2036_a_HPC2_and_U12 ( .A1(cell_2036_a_HPC2_and_a_reg[1]), .A2(
        cell_2036_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2036_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2036_a_HPC2_and_U11 ( .A1(cell_2036_a_HPC2_and_a_reg[0]), .A2(
        cell_2036_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2036_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2036_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2036_a_HPC2_and_n9), 
        .ZN(cell_2036_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2036_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2036_a_HPC2_and_n9), 
        .ZN(cell_2036_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2036_a_HPC2_and_U8 ( .A(Fresh[322]), .ZN(cell_2036_a_HPC2_and_n9) );
  AND2_X1 cell_2036_a_HPC2_and_U7 ( .A1(cell_2036_and_in[1]), .A2(n469), .ZN(
        cell_2036_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2036_a_HPC2_and_U6 ( .A1(cell_2036_and_in[0]), .A2(n465), .ZN(
        cell_2036_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2036_a_HPC2_and_U5 ( .A(cell_2036_a_HPC2_and_n8), .B(
        cell_2036_a_HPC2_and_z_1__1_), .ZN(cell_2036_and_out[1]) );
  XNOR2_X1 cell_2036_a_HPC2_and_U4 ( .A(
        cell_2036_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2036_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2036_a_HPC2_and_n8) );
  XNOR2_X1 cell_2036_a_HPC2_and_U3 ( .A(cell_2036_a_HPC2_and_n7), .B(
        cell_2036_a_HPC2_and_z_0__0_), .ZN(cell_2036_and_out[0]) );
  XNOR2_X1 cell_2036_a_HPC2_and_U2 ( .A(
        cell_2036_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2036_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2036_a_HPC2_and_n7) );
  DFF_X1 cell_2036_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2036_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2036_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2036_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2036_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2036_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2036_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2036_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2036_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2036_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2037_U4 ( .A(signal_3768), .B(cell_2037_and_out[1]), .Z(
        signal_3951) );
  XOR2_X1 cell_2037_U3 ( .A(signal_2258), .B(cell_2037_and_out[0]), .Z(
        signal_2305) );
  XOR2_X1 cell_2037_U2 ( .A(signal_3768), .B(signal_3706), .Z(
        cell_2037_and_in[1]) );
  XOR2_X1 cell_2037_U1 ( .A(signal_2258), .B(signal_2196), .Z(
        cell_2037_and_in[0]) );
  XOR2_X1 cell_2037_a_HPC2_and_U14 ( .A(Fresh[323]), .B(cell_2037_and_in[0]), 
        .Z(cell_2037_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2037_a_HPC2_and_U13 ( .A(Fresh[323]), .B(cell_2037_and_in[1]), 
        .Z(cell_2037_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2037_a_HPC2_and_U12 ( .A1(cell_2037_a_HPC2_and_a_reg[1]), .A2(
        cell_2037_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2037_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2037_a_HPC2_and_U11 ( .A1(cell_2037_a_HPC2_and_a_reg[0]), .A2(
        cell_2037_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2037_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2037_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2037_a_HPC2_and_n9), 
        .ZN(cell_2037_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2037_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2037_a_HPC2_and_n9), 
        .ZN(cell_2037_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2037_a_HPC2_and_U8 ( .A(Fresh[323]), .ZN(cell_2037_a_HPC2_and_n9) );
  AND2_X1 cell_2037_a_HPC2_and_U7 ( .A1(cell_2037_and_in[1]), .A2(n466), .ZN(
        cell_2037_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2037_a_HPC2_and_U6 ( .A1(cell_2037_and_in[0]), .A2(n462), .ZN(
        cell_2037_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2037_a_HPC2_and_U5 ( .A(cell_2037_a_HPC2_and_n8), .B(
        cell_2037_a_HPC2_and_z_1__1_), .ZN(cell_2037_and_out[1]) );
  XNOR2_X1 cell_2037_a_HPC2_and_U4 ( .A(
        cell_2037_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2037_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2037_a_HPC2_and_n8) );
  XNOR2_X1 cell_2037_a_HPC2_and_U3 ( .A(cell_2037_a_HPC2_and_n7), .B(
        cell_2037_a_HPC2_and_z_0__0_), .ZN(cell_2037_and_out[0]) );
  XNOR2_X1 cell_2037_a_HPC2_and_U2 ( .A(
        cell_2037_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2037_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2037_a_HPC2_and_n7) );
  DFF_X1 cell_2037_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2037_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2037_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2037_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2037_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2037_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2037_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2037_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2037_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2037_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2038_U4 ( .A(signal_3663), .B(cell_2038_and_out[1]), .Z(
        signal_3952) );
  XOR2_X1 cell_2038_U3 ( .A(signal_2153), .B(cell_2038_and_out[0]), .Z(
        signal_2306) );
  XOR2_X1 cell_2038_U2 ( .A(signal_3663), .B(signal_3779), .Z(
        cell_2038_and_in[1]) );
  XOR2_X1 cell_2038_U1 ( .A(signal_2153), .B(signal_2269), .Z(
        cell_2038_and_in[0]) );
  XOR2_X1 cell_2038_a_HPC2_and_U14 ( .A(Fresh[324]), .B(cell_2038_and_in[0]), 
        .Z(cell_2038_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2038_a_HPC2_and_U13 ( .A(Fresh[324]), .B(cell_2038_and_in[1]), 
        .Z(cell_2038_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2038_a_HPC2_and_U12 ( .A1(cell_2038_a_HPC2_and_a_reg[1]), .A2(
        cell_2038_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2038_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2038_a_HPC2_and_U11 ( .A1(cell_2038_a_HPC2_and_a_reg[0]), .A2(
        cell_2038_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2038_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2038_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2038_a_HPC2_and_n9), 
        .ZN(cell_2038_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2038_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2038_a_HPC2_and_n9), 
        .ZN(cell_2038_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2038_a_HPC2_and_U8 ( .A(Fresh[324]), .ZN(cell_2038_a_HPC2_and_n9) );
  AND2_X1 cell_2038_a_HPC2_and_U7 ( .A1(cell_2038_and_in[1]), .A2(n467), .ZN(
        cell_2038_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2038_a_HPC2_and_U6 ( .A1(cell_2038_and_in[0]), .A2(n463), .ZN(
        cell_2038_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2038_a_HPC2_and_U5 ( .A(cell_2038_a_HPC2_and_n8), .B(
        cell_2038_a_HPC2_and_z_1__1_), .ZN(cell_2038_and_out[1]) );
  XNOR2_X1 cell_2038_a_HPC2_and_U4 ( .A(
        cell_2038_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2038_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2038_a_HPC2_and_n8) );
  XNOR2_X1 cell_2038_a_HPC2_and_U3 ( .A(cell_2038_a_HPC2_and_n7), .B(
        cell_2038_a_HPC2_and_z_0__0_), .ZN(cell_2038_and_out[0]) );
  XNOR2_X1 cell_2038_a_HPC2_and_U2 ( .A(
        cell_2038_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2038_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2038_a_HPC2_and_n7) );
  DFF_X1 cell_2038_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2038_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2038_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2038_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2038_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2038_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2038_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2038_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2038_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2038_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2039_U4 ( .A(signal_3682), .B(cell_2039_and_out[1]), .Z(
        signal_3953) );
  XOR2_X1 cell_2039_U3 ( .A(signal_2172), .B(cell_2039_and_out[0]), .Z(
        signal_2307) );
  XOR2_X1 cell_2039_U2 ( .A(signal_3682), .B(signal_3665), .Z(
        cell_2039_and_in[1]) );
  XOR2_X1 cell_2039_U1 ( .A(signal_2172), .B(signal_2155), .Z(
        cell_2039_and_in[0]) );
  XOR2_X1 cell_2039_a_HPC2_and_U14 ( .A(Fresh[325]), .B(cell_2039_and_in[0]), 
        .Z(cell_2039_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2039_a_HPC2_and_U13 ( .A(Fresh[325]), .B(cell_2039_and_in[1]), 
        .Z(cell_2039_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2039_a_HPC2_and_U12 ( .A1(cell_2039_a_HPC2_and_a_reg[1]), .A2(
        cell_2039_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2039_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2039_a_HPC2_and_U11 ( .A1(cell_2039_a_HPC2_and_a_reg[0]), .A2(
        cell_2039_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2039_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2039_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2039_a_HPC2_and_n9), 
        .ZN(cell_2039_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2039_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2039_a_HPC2_and_n9), 
        .ZN(cell_2039_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2039_a_HPC2_and_U8 ( .A(Fresh[325]), .ZN(cell_2039_a_HPC2_and_n9) );
  AND2_X1 cell_2039_a_HPC2_and_U7 ( .A1(cell_2039_and_in[1]), .A2(n468), .ZN(
        cell_2039_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2039_a_HPC2_and_U6 ( .A1(cell_2039_and_in[0]), .A2(n464), .ZN(
        cell_2039_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2039_a_HPC2_and_U5 ( .A(cell_2039_a_HPC2_and_n8), .B(
        cell_2039_a_HPC2_and_z_1__1_), .ZN(cell_2039_and_out[1]) );
  XNOR2_X1 cell_2039_a_HPC2_and_U4 ( .A(
        cell_2039_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2039_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2039_a_HPC2_and_n8) );
  XNOR2_X1 cell_2039_a_HPC2_and_U3 ( .A(cell_2039_a_HPC2_and_n7), .B(
        cell_2039_a_HPC2_and_z_0__0_), .ZN(cell_2039_and_out[0]) );
  XNOR2_X1 cell_2039_a_HPC2_and_U2 ( .A(
        cell_2039_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2039_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2039_a_HPC2_and_n7) );
  DFF_X1 cell_2039_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2039_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2039_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2039_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2039_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2039_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2039_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2039_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2039_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2039_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2040_U4 ( .A(signal_3748), .B(cell_2040_and_out[1]), .Z(
        signal_3954) );
  XOR2_X1 cell_2040_U3 ( .A(signal_2238), .B(cell_2040_and_out[0]), .Z(
        signal_2308) );
  XOR2_X1 cell_2040_U2 ( .A(signal_3748), .B(signal_3776), .Z(
        cell_2040_and_in[1]) );
  XOR2_X1 cell_2040_U1 ( .A(signal_2238), .B(signal_2266), .Z(
        cell_2040_and_in[0]) );
  XOR2_X1 cell_2040_a_HPC2_and_U14 ( .A(Fresh[326]), .B(cell_2040_and_in[0]), 
        .Z(cell_2040_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2040_a_HPC2_and_U13 ( .A(Fresh[326]), .B(cell_2040_and_in[1]), 
        .Z(cell_2040_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2040_a_HPC2_and_U12 ( .A1(cell_2040_a_HPC2_and_a_reg[1]), .A2(
        cell_2040_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2040_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2040_a_HPC2_and_U11 ( .A1(cell_2040_a_HPC2_and_a_reg[0]), .A2(
        cell_2040_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2040_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2040_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2040_a_HPC2_and_n9), 
        .ZN(cell_2040_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2040_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2040_a_HPC2_and_n9), 
        .ZN(cell_2040_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2040_a_HPC2_and_U8 ( .A(Fresh[326]), .ZN(cell_2040_a_HPC2_and_n9) );
  AND2_X1 cell_2040_a_HPC2_and_U7 ( .A1(cell_2040_and_in[1]), .A2(n466), .ZN(
        cell_2040_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2040_a_HPC2_and_U6 ( .A1(cell_2040_and_in[0]), .A2(n462), .ZN(
        cell_2040_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2040_a_HPC2_and_U5 ( .A(cell_2040_a_HPC2_and_n8), .B(
        cell_2040_a_HPC2_and_z_1__1_), .ZN(cell_2040_and_out[1]) );
  XNOR2_X1 cell_2040_a_HPC2_and_U4 ( .A(
        cell_2040_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2040_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2040_a_HPC2_and_n8) );
  XNOR2_X1 cell_2040_a_HPC2_and_U3 ( .A(cell_2040_a_HPC2_and_n7), .B(
        cell_2040_a_HPC2_and_z_0__0_), .ZN(cell_2040_and_out[0]) );
  XNOR2_X1 cell_2040_a_HPC2_and_U2 ( .A(
        cell_2040_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2040_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2040_a_HPC2_and_n7) );
  DFF_X1 cell_2040_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2040_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2040_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2040_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2040_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2040_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2040_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2040_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2040_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2040_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2041_U4 ( .A(signal_3751), .B(cell_2041_and_out[1]), .Z(
        signal_3955) );
  XOR2_X1 cell_2041_U3 ( .A(signal_2241), .B(cell_2041_and_out[0]), .Z(
        signal_2309) );
  XOR2_X1 cell_2041_U2 ( .A(signal_3751), .B(signal_3686), .Z(
        cell_2041_and_in[1]) );
  XOR2_X1 cell_2041_U1 ( .A(signal_2241), .B(signal_2176), .Z(
        cell_2041_and_in[0]) );
  XOR2_X1 cell_2041_a_HPC2_and_U14 ( .A(Fresh[327]), .B(cell_2041_and_in[0]), 
        .Z(cell_2041_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2041_a_HPC2_and_U13 ( .A(Fresh[327]), .B(cell_2041_and_in[1]), 
        .Z(cell_2041_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2041_a_HPC2_and_U12 ( .A1(cell_2041_a_HPC2_and_a_reg[1]), .A2(
        cell_2041_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2041_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2041_a_HPC2_and_U11 ( .A1(cell_2041_a_HPC2_and_a_reg[0]), .A2(
        cell_2041_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2041_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2041_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2041_a_HPC2_and_n9), 
        .ZN(cell_2041_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2041_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2041_a_HPC2_and_n9), 
        .ZN(cell_2041_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2041_a_HPC2_and_U8 ( .A(Fresh[327]), .ZN(cell_2041_a_HPC2_and_n9) );
  AND2_X1 cell_2041_a_HPC2_and_U7 ( .A1(cell_2041_and_in[1]), .A2(n466), .ZN(
        cell_2041_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2041_a_HPC2_and_U6 ( .A1(cell_2041_and_in[0]), .A2(n462), .ZN(
        cell_2041_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2041_a_HPC2_and_U5 ( .A(cell_2041_a_HPC2_and_n8), .B(
        cell_2041_a_HPC2_and_z_1__1_), .ZN(cell_2041_and_out[1]) );
  XNOR2_X1 cell_2041_a_HPC2_and_U4 ( .A(
        cell_2041_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2041_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2041_a_HPC2_and_n8) );
  XNOR2_X1 cell_2041_a_HPC2_and_U3 ( .A(cell_2041_a_HPC2_and_n7), .B(
        cell_2041_a_HPC2_and_z_0__0_), .ZN(cell_2041_and_out[0]) );
  XNOR2_X1 cell_2041_a_HPC2_and_U2 ( .A(
        cell_2041_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2041_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2041_a_HPC2_and_n7) );
  DFF_X1 cell_2041_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2041_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2041_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2041_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2041_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2041_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2041_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2041_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2041_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2041_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2042_U4 ( .A(signal_3664), .B(cell_2042_and_out[1]), .Z(
        signal_3956) );
  XOR2_X1 cell_2042_U3 ( .A(signal_2154), .B(cell_2042_and_out[0]), .Z(
        signal_2310) );
  XOR2_X1 cell_2042_U2 ( .A(signal_3664), .B(signal_3733), .Z(
        cell_2042_and_in[1]) );
  XOR2_X1 cell_2042_U1 ( .A(signal_2154), .B(signal_2223), .Z(
        cell_2042_and_in[0]) );
  XOR2_X1 cell_2042_a_HPC2_and_U14 ( .A(Fresh[328]), .B(cell_2042_and_in[0]), 
        .Z(cell_2042_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2042_a_HPC2_and_U13 ( .A(Fresh[328]), .B(cell_2042_and_in[1]), 
        .Z(cell_2042_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2042_a_HPC2_and_U12 ( .A1(cell_2042_a_HPC2_and_a_reg[1]), .A2(
        cell_2042_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2042_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2042_a_HPC2_and_U11 ( .A1(cell_2042_a_HPC2_and_a_reg[0]), .A2(
        cell_2042_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2042_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2042_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2042_a_HPC2_and_n9), 
        .ZN(cell_2042_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2042_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2042_a_HPC2_and_n9), 
        .ZN(cell_2042_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2042_a_HPC2_and_U8 ( .A(Fresh[328]), .ZN(cell_2042_a_HPC2_and_n9) );
  AND2_X1 cell_2042_a_HPC2_and_U7 ( .A1(cell_2042_and_in[1]), .A2(n466), .ZN(
        cell_2042_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2042_a_HPC2_and_U6 ( .A1(cell_2042_and_in[0]), .A2(n462), .ZN(
        cell_2042_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2042_a_HPC2_and_U5 ( .A(cell_2042_a_HPC2_and_n8), .B(
        cell_2042_a_HPC2_and_z_1__1_), .ZN(cell_2042_and_out[1]) );
  XNOR2_X1 cell_2042_a_HPC2_and_U4 ( .A(
        cell_2042_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2042_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2042_a_HPC2_and_n8) );
  XNOR2_X1 cell_2042_a_HPC2_and_U3 ( .A(cell_2042_a_HPC2_and_n7), .B(
        cell_2042_a_HPC2_and_z_0__0_), .ZN(cell_2042_and_out[0]) );
  XNOR2_X1 cell_2042_a_HPC2_and_U2 ( .A(
        cell_2042_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2042_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2042_a_HPC2_and_n7) );
  DFF_X1 cell_2042_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2042_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2042_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2042_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2042_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2042_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2042_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2042_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2042_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2042_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2043_U4 ( .A(signal_3694), .B(cell_2043_and_out[1]), .Z(
        signal_3957) );
  XOR2_X1 cell_2043_U3 ( .A(signal_2184), .B(cell_2043_and_out[0]), .Z(
        signal_2311) );
  XOR2_X1 cell_2043_U2 ( .A(signal_3694), .B(signal_3745), .Z(
        cell_2043_and_in[1]) );
  XOR2_X1 cell_2043_U1 ( .A(signal_2184), .B(signal_2235), .Z(
        cell_2043_and_in[0]) );
  XOR2_X1 cell_2043_a_HPC2_and_U14 ( .A(Fresh[329]), .B(cell_2043_and_in[0]), 
        .Z(cell_2043_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2043_a_HPC2_and_U13 ( .A(Fresh[329]), .B(cell_2043_and_in[1]), 
        .Z(cell_2043_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2043_a_HPC2_and_U12 ( .A1(cell_2043_a_HPC2_and_a_reg[1]), .A2(
        cell_2043_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2043_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2043_a_HPC2_and_U11 ( .A1(cell_2043_a_HPC2_and_a_reg[0]), .A2(
        cell_2043_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2043_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2043_a_HPC2_and_U10 ( .A1(n466), .A2(cell_2043_a_HPC2_and_n9), 
        .ZN(cell_2043_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2043_a_HPC2_and_U9 ( .A1(n462), .A2(cell_2043_a_HPC2_and_n9), 
        .ZN(cell_2043_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2043_a_HPC2_and_U8 ( .A(Fresh[329]), .ZN(cell_2043_a_HPC2_and_n9) );
  AND2_X1 cell_2043_a_HPC2_and_U7 ( .A1(cell_2043_and_in[1]), .A2(n466), .ZN(
        cell_2043_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2043_a_HPC2_and_U6 ( .A1(cell_2043_and_in[0]), .A2(n462), .ZN(
        cell_2043_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2043_a_HPC2_and_U5 ( .A(cell_2043_a_HPC2_and_n8), .B(
        cell_2043_a_HPC2_and_z_1__1_), .ZN(cell_2043_and_out[1]) );
  XNOR2_X1 cell_2043_a_HPC2_and_U4 ( .A(
        cell_2043_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2043_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2043_a_HPC2_and_n8) );
  XNOR2_X1 cell_2043_a_HPC2_and_U3 ( .A(cell_2043_a_HPC2_and_n7), .B(
        cell_2043_a_HPC2_and_z_0__0_), .ZN(cell_2043_and_out[0]) );
  XNOR2_X1 cell_2043_a_HPC2_and_U2 ( .A(
        cell_2043_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2043_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2043_a_HPC2_and_n7) );
  DFF_X1 cell_2043_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2043_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2043_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n462), .CK(clk), 
        .Q(cell_2043_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2043_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2043_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n466), .CK(clk), 
        .Q(cell_2043_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2043_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2043_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2043_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2044_U4 ( .A(signal_3736), .B(cell_2044_and_out[1]), .Z(
        signal_3958) );
  XOR2_X1 cell_2044_U3 ( .A(signal_2226), .B(cell_2044_and_out[0]), .Z(
        signal_2312) );
  XOR2_X1 cell_2044_U2 ( .A(signal_3736), .B(signal_3683), .Z(
        cell_2044_and_in[1]) );
  XOR2_X1 cell_2044_U1 ( .A(signal_2226), .B(signal_2173), .Z(
        cell_2044_and_in[0]) );
  XOR2_X1 cell_2044_a_HPC2_and_U14 ( .A(Fresh[330]), .B(cell_2044_and_in[0]), 
        .Z(cell_2044_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2044_a_HPC2_and_U13 ( .A(Fresh[330]), .B(cell_2044_and_in[1]), 
        .Z(cell_2044_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2044_a_HPC2_and_U12 ( .A1(cell_2044_a_HPC2_and_a_reg[1]), .A2(
        cell_2044_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2044_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2044_a_HPC2_and_U11 ( .A1(cell_2044_a_HPC2_and_a_reg[0]), .A2(
        cell_2044_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2044_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2044_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2044_a_HPC2_and_n9), 
        .ZN(cell_2044_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2044_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2044_a_HPC2_and_n9), 
        .ZN(cell_2044_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2044_a_HPC2_and_U8 ( .A(Fresh[330]), .ZN(cell_2044_a_HPC2_and_n9) );
  AND2_X1 cell_2044_a_HPC2_and_U7 ( .A1(cell_2044_and_in[1]), .A2(n468), .ZN(
        cell_2044_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2044_a_HPC2_and_U6 ( .A1(cell_2044_and_in[0]), .A2(n464), .ZN(
        cell_2044_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2044_a_HPC2_and_U5 ( .A(cell_2044_a_HPC2_and_n8), .B(
        cell_2044_a_HPC2_and_z_1__1_), .ZN(cell_2044_and_out[1]) );
  XNOR2_X1 cell_2044_a_HPC2_and_U4 ( .A(
        cell_2044_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2044_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2044_a_HPC2_and_n8) );
  XNOR2_X1 cell_2044_a_HPC2_and_U3 ( .A(cell_2044_a_HPC2_and_n7), .B(
        cell_2044_a_HPC2_and_z_0__0_), .ZN(cell_2044_and_out[0]) );
  XNOR2_X1 cell_2044_a_HPC2_and_U2 ( .A(
        cell_2044_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2044_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2044_a_HPC2_and_n7) );
  DFF_X1 cell_2044_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2044_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2044_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2044_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2044_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2044_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2044_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2044_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2044_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2044_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2045_U4 ( .A(signal_3696), .B(cell_2045_and_out[1]), .Z(
        signal_3959) );
  XOR2_X1 cell_2045_U3 ( .A(signal_2186), .B(cell_2045_and_out[0]), .Z(
        signal_2313) );
  XOR2_X1 cell_2045_U2 ( .A(signal_3696), .B(signal_3719), .Z(
        cell_2045_and_in[1]) );
  XOR2_X1 cell_2045_U1 ( .A(signal_2186), .B(signal_2209), .Z(
        cell_2045_and_in[0]) );
  XOR2_X1 cell_2045_a_HPC2_and_U14 ( .A(Fresh[331]), .B(cell_2045_and_in[0]), 
        .Z(cell_2045_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2045_a_HPC2_and_U13 ( .A(Fresh[331]), .B(cell_2045_and_in[1]), 
        .Z(cell_2045_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2045_a_HPC2_and_U12 ( .A1(cell_2045_a_HPC2_and_a_reg[1]), .A2(
        cell_2045_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2045_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2045_a_HPC2_and_U11 ( .A1(cell_2045_a_HPC2_and_a_reg[0]), .A2(
        cell_2045_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2045_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2045_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2045_a_HPC2_and_n9), 
        .ZN(cell_2045_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2045_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2045_a_HPC2_and_n9), 
        .ZN(cell_2045_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2045_a_HPC2_and_U8 ( .A(Fresh[331]), .ZN(cell_2045_a_HPC2_and_n9) );
  AND2_X1 cell_2045_a_HPC2_and_U7 ( .A1(cell_2045_and_in[1]), .A2(n468), .ZN(
        cell_2045_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2045_a_HPC2_and_U6 ( .A1(cell_2045_and_in[0]), .A2(n464), .ZN(
        cell_2045_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2045_a_HPC2_and_U5 ( .A(cell_2045_a_HPC2_and_n8), .B(
        cell_2045_a_HPC2_and_z_1__1_), .ZN(cell_2045_and_out[1]) );
  XNOR2_X1 cell_2045_a_HPC2_and_U4 ( .A(
        cell_2045_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2045_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2045_a_HPC2_and_n8) );
  XNOR2_X1 cell_2045_a_HPC2_and_U3 ( .A(cell_2045_a_HPC2_and_n7), .B(
        cell_2045_a_HPC2_and_z_0__0_), .ZN(cell_2045_and_out[0]) );
  XNOR2_X1 cell_2045_a_HPC2_and_U2 ( .A(
        cell_2045_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2045_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2045_a_HPC2_and_n7) );
  DFF_X1 cell_2045_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2045_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2045_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2045_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2045_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2045_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2045_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2045_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2045_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2045_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2046_U4 ( .A(signal_3676), .B(cell_2046_and_out[1]), .Z(
        signal_3960) );
  XOR2_X1 cell_2046_U3 ( .A(signal_2166), .B(cell_2046_and_out[0]), .Z(
        signal_2314) );
  XOR2_X1 cell_2046_U2 ( .A(signal_3676), .B(signal_3685), .Z(
        cell_2046_and_in[1]) );
  XOR2_X1 cell_2046_U1 ( .A(signal_2166), .B(signal_2175), .Z(
        cell_2046_and_in[0]) );
  XOR2_X1 cell_2046_a_HPC2_and_U14 ( .A(Fresh[332]), .B(cell_2046_and_in[0]), 
        .Z(cell_2046_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2046_a_HPC2_and_U13 ( .A(Fresh[332]), .B(cell_2046_and_in[1]), 
        .Z(cell_2046_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2046_a_HPC2_and_U12 ( .A1(cell_2046_a_HPC2_and_a_reg[1]), .A2(
        cell_2046_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2046_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2046_a_HPC2_and_U11 ( .A1(cell_2046_a_HPC2_and_a_reg[0]), .A2(
        cell_2046_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2046_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2046_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2046_a_HPC2_and_n9), 
        .ZN(cell_2046_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2046_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2046_a_HPC2_and_n9), 
        .ZN(cell_2046_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2046_a_HPC2_and_U8 ( .A(Fresh[332]), .ZN(cell_2046_a_HPC2_and_n9) );
  AND2_X1 cell_2046_a_HPC2_and_U7 ( .A1(cell_2046_and_in[1]), .A2(n468), .ZN(
        cell_2046_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2046_a_HPC2_and_U6 ( .A1(cell_2046_and_in[0]), .A2(n464), .ZN(
        cell_2046_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2046_a_HPC2_and_U5 ( .A(cell_2046_a_HPC2_and_n8), .B(
        cell_2046_a_HPC2_and_z_1__1_), .ZN(cell_2046_and_out[1]) );
  XNOR2_X1 cell_2046_a_HPC2_and_U4 ( .A(
        cell_2046_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2046_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2046_a_HPC2_and_n8) );
  XNOR2_X1 cell_2046_a_HPC2_and_U3 ( .A(cell_2046_a_HPC2_and_n7), .B(
        cell_2046_a_HPC2_and_z_0__0_), .ZN(cell_2046_and_out[0]) );
  XNOR2_X1 cell_2046_a_HPC2_and_U2 ( .A(
        cell_2046_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2046_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2046_a_HPC2_and_n7) );
  DFF_X1 cell_2046_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2046_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2046_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2046_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2046_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2046_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2046_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2046_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2046_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2046_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2047_U4 ( .A(signal_3732), .B(cell_2047_and_out[1]), .Z(
        signal_3961) );
  XOR2_X1 cell_2047_U3 ( .A(signal_2222), .B(cell_2047_and_out[0]), .Z(
        signal_2315) );
  XOR2_X1 cell_2047_U2 ( .A(signal_3732), .B(signal_3752), .Z(
        cell_2047_and_in[1]) );
  XOR2_X1 cell_2047_U1 ( .A(signal_2222), .B(signal_2242), .Z(
        cell_2047_and_in[0]) );
  XOR2_X1 cell_2047_a_HPC2_and_U14 ( .A(Fresh[333]), .B(cell_2047_and_in[0]), 
        .Z(cell_2047_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2047_a_HPC2_and_U13 ( .A(Fresh[333]), .B(cell_2047_and_in[1]), 
        .Z(cell_2047_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2047_a_HPC2_and_U12 ( .A1(cell_2047_a_HPC2_and_a_reg[1]), .A2(
        cell_2047_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2047_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2047_a_HPC2_and_U11 ( .A1(cell_2047_a_HPC2_and_a_reg[0]), .A2(
        cell_2047_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2047_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2047_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2047_a_HPC2_and_n9), 
        .ZN(cell_2047_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2047_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2047_a_HPC2_and_n9), 
        .ZN(cell_2047_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2047_a_HPC2_and_U8 ( .A(Fresh[333]), .ZN(cell_2047_a_HPC2_and_n9) );
  AND2_X1 cell_2047_a_HPC2_and_U7 ( .A1(cell_2047_and_in[1]), .A2(n468), .ZN(
        cell_2047_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2047_a_HPC2_and_U6 ( .A1(cell_2047_and_in[0]), .A2(n464), .ZN(
        cell_2047_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2047_a_HPC2_and_U5 ( .A(cell_2047_a_HPC2_and_n8), .B(
        cell_2047_a_HPC2_and_z_1__1_), .ZN(cell_2047_and_out[1]) );
  XNOR2_X1 cell_2047_a_HPC2_and_U4 ( .A(
        cell_2047_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2047_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2047_a_HPC2_and_n8) );
  XNOR2_X1 cell_2047_a_HPC2_and_U3 ( .A(cell_2047_a_HPC2_and_n7), .B(
        cell_2047_a_HPC2_and_z_0__0_), .ZN(cell_2047_and_out[0]) );
  XNOR2_X1 cell_2047_a_HPC2_and_U2 ( .A(
        cell_2047_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2047_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2047_a_HPC2_and_n7) );
  DFF_X1 cell_2047_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2047_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2047_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2047_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2047_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2047_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2047_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2047_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2047_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2047_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2048_U4 ( .A(signal_3734), .B(cell_2048_and_out[1]), .Z(
        signal_3962) );
  XOR2_X1 cell_2048_U3 ( .A(signal_2224), .B(cell_2048_and_out[0]), .Z(
        signal_2316) );
  XOR2_X1 cell_2048_U2 ( .A(signal_3734), .B(signal_3700), .Z(
        cell_2048_and_in[1]) );
  XOR2_X1 cell_2048_U1 ( .A(signal_2224), .B(signal_2190), .Z(
        cell_2048_and_in[0]) );
  XOR2_X1 cell_2048_a_HPC2_and_U14 ( .A(Fresh[334]), .B(cell_2048_and_in[0]), 
        .Z(cell_2048_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2048_a_HPC2_and_U13 ( .A(Fresh[334]), .B(cell_2048_and_in[1]), 
        .Z(cell_2048_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2048_a_HPC2_and_U12 ( .A1(cell_2048_a_HPC2_and_a_reg[1]), .A2(
        cell_2048_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2048_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2048_a_HPC2_and_U11 ( .A1(cell_2048_a_HPC2_and_a_reg[0]), .A2(
        cell_2048_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2048_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2048_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2048_a_HPC2_and_n9), 
        .ZN(cell_2048_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2048_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2048_a_HPC2_and_n9), 
        .ZN(cell_2048_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2048_a_HPC2_and_U8 ( .A(Fresh[334]), .ZN(cell_2048_a_HPC2_and_n9) );
  AND2_X1 cell_2048_a_HPC2_and_U7 ( .A1(cell_2048_and_in[1]), .A2(n468), .ZN(
        cell_2048_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2048_a_HPC2_and_U6 ( .A1(cell_2048_and_in[0]), .A2(n464), .ZN(
        cell_2048_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2048_a_HPC2_and_U5 ( .A(cell_2048_a_HPC2_and_n8), .B(
        cell_2048_a_HPC2_and_z_1__1_), .ZN(cell_2048_and_out[1]) );
  XNOR2_X1 cell_2048_a_HPC2_and_U4 ( .A(
        cell_2048_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2048_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2048_a_HPC2_and_n8) );
  XNOR2_X1 cell_2048_a_HPC2_and_U3 ( .A(cell_2048_a_HPC2_and_n7), .B(
        cell_2048_a_HPC2_and_z_0__0_), .ZN(cell_2048_and_out[0]) );
  XNOR2_X1 cell_2048_a_HPC2_and_U2 ( .A(
        cell_2048_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2048_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2048_a_HPC2_and_n7) );
  DFF_X1 cell_2048_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2048_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2048_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2048_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2048_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2048_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2048_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2048_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2048_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2048_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2049_U4 ( .A(signal_3684), .B(cell_2049_and_out[1]), .Z(
        signal_3963) );
  XOR2_X1 cell_2049_U3 ( .A(signal_2174), .B(cell_2049_and_out[0]), .Z(
        signal_2317) );
  XOR2_X1 cell_2049_U2 ( .A(signal_3684), .B(signal_3762), .Z(
        cell_2049_and_in[1]) );
  XOR2_X1 cell_2049_U1 ( .A(signal_2174), .B(signal_2252), .Z(
        cell_2049_and_in[0]) );
  XOR2_X1 cell_2049_a_HPC2_and_U14 ( .A(Fresh[335]), .B(cell_2049_and_in[0]), 
        .Z(cell_2049_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2049_a_HPC2_and_U13 ( .A(Fresh[335]), .B(cell_2049_and_in[1]), 
        .Z(cell_2049_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2049_a_HPC2_and_U12 ( .A1(cell_2049_a_HPC2_and_a_reg[1]), .A2(
        cell_2049_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2049_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2049_a_HPC2_and_U11 ( .A1(cell_2049_a_HPC2_and_a_reg[0]), .A2(
        cell_2049_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2049_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2049_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2049_a_HPC2_and_n9), 
        .ZN(cell_2049_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2049_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2049_a_HPC2_and_n9), 
        .ZN(cell_2049_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2049_a_HPC2_and_U8 ( .A(Fresh[335]), .ZN(cell_2049_a_HPC2_and_n9) );
  AND2_X1 cell_2049_a_HPC2_and_U7 ( .A1(cell_2049_and_in[1]), .A2(n468), .ZN(
        cell_2049_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2049_a_HPC2_and_U6 ( .A1(cell_2049_and_in[0]), .A2(n464), .ZN(
        cell_2049_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2049_a_HPC2_and_U5 ( .A(cell_2049_a_HPC2_and_n8), .B(
        cell_2049_a_HPC2_and_z_1__1_), .ZN(cell_2049_and_out[1]) );
  XNOR2_X1 cell_2049_a_HPC2_and_U4 ( .A(
        cell_2049_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2049_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2049_a_HPC2_and_n8) );
  XNOR2_X1 cell_2049_a_HPC2_and_U3 ( .A(cell_2049_a_HPC2_and_n7), .B(
        cell_2049_a_HPC2_and_z_0__0_), .ZN(cell_2049_and_out[0]) );
  XNOR2_X1 cell_2049_a_HPC2_and_U2 ( .A(
        cell_2049_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2049_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2049_a_HPC2_and_n7) );
  DFF_X1 cell_2049_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2049_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2049_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2049_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2049_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2049_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2049_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2049_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2049_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2049_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2050_U4 ( .A(signal_3704), .B(cell_2050_and_out[1]), .Z(
        signal_3964) );
  XOR2_X1 cell_2050_U3 ( .A(signal_2194), .B(cell_2050_and_out[0]), .Z(
        signal_2318) );
  XOR2_X1 cell_2050_U2 ( .A(signal_3704), .B(signal_3680), .Z(
        cell_2050_and_in[1]) );
  XOR2_X1 cell_2050_U1 ( .A(signal_2194), .B(signal_2170), .Z(
        cell_2050_and_in[0]) );
  XOR2_X1 cell_2050_a_HPC2_and_U14 ( .A(Fresh[336]), .B(cell_2050_and_in[0]), 
        .Z(cell_2050_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2050_a_HPC2_and_U13 ( .A(Fresh[336]), .B(cell_2050_and_in[1]), 
        .Z(cell_2050_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2050_a_HPC2_and_U12 ( .A1(cell_2050_a_HPC2_and_a_reg[1]), .A2(
        cell_2050_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2050_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2050_a_HPC2_and_U11 ( .A1(cell_2050_a_HPC2_and_a_reg[0]), .A2(
        cell_2050_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2050_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2050_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2050_a_HPC2_and_n9), 
        .ZN(cell_2050_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2050_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2050_a_HPC2_and_n9), 
        .ZN(cell_2050_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2050_a_HPC2_and_U8 ( .A(Fresh[336]), .ZN(cell_2050_a_HPC2_and_n9) );
  AND2_X1 cell_2050_a_HPC2_and_U7 ( .A1(cell_2050_and_in[1]), .A2(n468), .ZN(
        cell_2050_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2050_a_HPC2_and_U6 ( .A1(cell_2050_and_in[0]), .A2(n464), .ZN(
        cell_2050_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2050_a_HPC2_and_U5 ( .A(cell_2050_a_HPC2_and_n8), .B(
        cell_2050_a_HPC2_and_z_1__1_), .ZN(cell_2050_and_out[1]) );
  XNOR2_X1 cell_2050_a_HPC2_and_U4 ( .A(
        cell_2050_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2050_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2050_a_HPC2_and_n8) );
  XNOR2_X1 cell_2050_a_HPC2_and_U3 ( .A(cell_2050_a_HPC2_and_n7), .B(
        cell_2050_a_HPC2_and_z_0__0_), .ZN(cell_2050_and_out[0]) );
  XNOR2_X1 cell_2050_a_HPC2_and_U2 ( .A(
        cell_2050_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2050_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2050_a_HPC2_and_n7) );
  DFF_X1 cell_2050_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2050_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2050_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2050_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2050_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2050_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2050_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2050_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2050_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2050_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2051_U4 ( .A(signal_3671), .B(cell_2051_and_out[1]), .Z(
        signal_3965) );
  XOR2_X1 cell_2051_U3 ( .A(signal_2161), .B(cell_2051_and_out[0]), .Z(
        signal_2319) );
  XOR2_X1 cell_2051_U2 ( .A(signal_3671), .B(signal_3757), .Z(
        cell_2051_and_in[1]) );
  XOR2_X1 cell_2051_U1 ( .A(signal_2161), .B(signal_2247), .Z(
        cell_2051_and_in[0]) );
  XOR2_X1 cell_2051_a_HPC2_and_U14 ( .A(Fresh[337]), .B(cell_2051_and_in[0]), 
        .Z(cell_2051_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2051_a_HPC2_and_U13 ( .A(Fresh[337]), .B(cell_2051_and_in[1]), 
        .Z(cell_2051_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2051_a_HPC2_and_U12 ( .A1(cell_2051_a_HPC2_and_a_reg[1]), .A2(
        cell_2051_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2051_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2051_a_HPC2_and_U11 ( .A1(cell_2051_a_HPC2_and_a_reg[0]), .A2(
        cell_2051_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2051_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2051_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2051_a_HPC2_and_n9), 
        .ZN(cell_2051_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2051_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2051_a_HPC2_and_n9), 
        .ZN(cell_2051_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2051_a_HPC2_and_U8 ( .A(Fresh[337]), .ZN(cell_2051_a_HPC2_and_n9) );
  AND2_X1 cell_2051_a_HPC2_and_U7 ( .A1(cell_2051_and_in[1]), .A2(n468), .ZN(
        cell_2051_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2051_a_HPC2_and_U6 ( .A1(cell_2051_and_in[0]), .A2(n464), .ZN(
        cell_2051_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2051_a_HPC2_and_U5 ( .A(cell_2051_a_HPC2_and_n8), .B(
        cell_2051_a_HPC2_and_z_1__1_), .ZN(cell_2051_and_out[1]) );
  XNOR2_X1 cell_2051_a_HPC2_and_U4 ( .A(
        cell_2051_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2051_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2051_a_HPC2_and_n8) );
  XNOR2_X1 cell_2051_a_HPC2_and_U3 ( .A(cell_2051_a_HPC2_and_n7), .B(
        cell_2051_a_HPC2_and_z_0__0_), .ZN(cell_2051_and_out[0]) );
  XNOR2_X1 cell_2051_a_HPC2_and_U2 ( .A(
        cell_2051_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2051_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2051_a_HPC2_and_n7) );
  DFF_X1 cell_2051_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2051_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2051_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2051_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2051_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2051_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2051_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2051_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2051_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2051_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2052_U4 ( .A(signal_3720), .B(cell_2052_and_out[1]), .Z(
        signal_3966) );
  XOR2_X1 cell_2052_U3 ( .A(signal_2210), .B(cell_2052_and_out[0]), .Z(
        signal_2320) );
  XOR2_X1 cell_2052_U2 ( .A(signal_3720), .B(signal_3714), .Z(
        cell_2052_and_in[1]) );
  XOR2_X1 cell_2052_U1 ( .A(signal_2210), .B(signal_2204), .Z(
        cell_2052_and_in[0]) );
  XOR2_X1 cell_2052_a_HPC2_and_U14 ( .A(Fresh[338]), .B(cell_2052_and_in[0]), 
        .Z(cell_2052_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2052_a_HPC2_and_U13 ( .A(Fresh[338]), .B(cell_2052_and_in[1]), 
        .Z(cell_2052_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2052_a_HPC2_and_U12 ( .A1(cell_2052_a_HPC2_and_a_reg[1]), .A2(
        cell_2052_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2052_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2052_a_HPC2_and_U11 ( .A1(cell_2052_a_HPC2_and_a_reg[0]), .A2(
        cell_2052_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2052_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2052_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2052_a_HPC2_and_n9), 
        .ZN(cell_2052_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2052_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2052_a_HPC2_and_n9), 
        .ZN(cell_2052_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2052_a_HPC2_and_U8 ( .A(Fresh[338]), .ZN(cell_2052_a_HPC2_and_n9) );
  AND2_X1 cell_2052_a_HPC2_and_U7 ( .A1(cell_2052_and_in[1]), .A2(n468), .ZN(
        cell_2052_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2052_a_HPC2_and_U6 ( .A1(cell_2052_and_in[0]), .A2(n464), .ZN(
        cell_2052_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2052_a_HPC2_and_U5 ( .A(cell_2052_a_HPC2_and_n8), .B(
        cell_2052_a_HPC2_and_z_1__1_), .ZN(cell_2052_and_out[1]) );
  XNOR2_X1 cell_2052_a_HPC2_and_U4 ( .A(
        cell_2052_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2052_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2052_a_HPC2_and_n8) );
  XNOR2_X1 cell_2052_a_HPC2_and_U3 ( .A(cell_2052_a_HPC2_and_n7), .B(
        cell_2052_a_HPC2_and_z_0__0_), .ZN(cell_2052_and_out[0]) );
  XNOR2_X1 cell_2052_a_HPC2_and_U2 ( .A(
        cell_2052_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2052_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2052_a_HPC2_and_n7) );
  DFF_X1 cell_2052_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2052_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2052_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2052_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2052_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2052_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2052_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2052_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2052_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2052_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2053_U4 ( .A(signal_3739), .B(cell_2053_and_out[1]), .Z(
        signal_3967) );
  XOR2_X1 cell_2053_U3 ( .A(signal_2229), .B(cell_2053_and_out[0]), .Z(
        signal_2321) );
  XOR2_X1 cell_2053_U2 ( .A(signal_3739), .B(signal_3672), .Z(
        cell_2053_and_in[1]) );
  XOR2_X1 cell_2053_U1 ( .A(signal_2229), .B(signal_2162), .Z(
        cell_2053_and_in[0]) );
  XOR2_X1 cell_2053_a_HPC2_and_U14 ( .A(Fresh[339]), .B(cell_2053_and_in[0]), 
        .Z(cell_2053_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2053_a_HPC2_and_U13 ( .A(Fresh[339]), .B(cell_2053_and_in[1]), 
        .Z(cell_2053_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2053_a_HPC2_and_U12 ( .A1(cell_2053_a_HPC2_and_a_reg[1]), .A2(
        cell_2053_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2053_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2053_a_HPC2_and_U11 ( .A1(cell_2053_a_HPC2_and_a_reg[0]), .A2(
        cell_2053_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2053_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2053_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2053_a_HPC2_and_n9), 
        .ZN(cell_2053_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2053_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2053_a_HPC2_and_n9), 
        .ZN(cell_2053_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2053_a_HPC2_and_U8 ( .A(Fresh[339]), .ZN(cell_2053_a_HPC2_and_n9) );
  AND2_X1 cell_2053_a_HPC2_and_U7 ( .A1(cell_2053_and_in[1]), .A2(n468), .ZN(
        cell_2053_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2053_a_HPC2_and_U6 ( .A1(cell_2053_and_in[0]), .A2(n464), .ZN(
        cell_2053_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2053_a_HPC2_and_U5 ( .A(cell_2053_a_HPC2_and_n8), .B(
        cell_2053_a_HPC2_and_z_1__1_), .ZN(cell_2053_and_out[1]) );
  XNOR2_X1 cell_2053_a_HPC2_and_U4 ( .A(
        cell_2053_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2053_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2053_a_HPC2_and_n8) );
  XNOR2_X1 cell_2053_a_HPC2_and_U3 ( .A(cell_2053_a_HPC2_and_n7), .B(
        cell_2053_a_HPC2_and_z_0__0_), .ZN(cell_2053_and_out[0]) );
  XNOR2_X1 cell_2053_a_HPC2_and_U2 ( .A(
        cell_2053_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2053_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2053_a_HPC2_and_n7) );
  DFF_X1 cell_2053_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2053_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2053_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2053_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2053_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2053_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2053_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2053_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2053_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2053_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2054_U4 ( .A(signal_3666), .B(cell_2054_and_out[1]), .Z(
        signal_3968) );
  XOR2_X1 cell_2054_U3 ( .A(signal_2156), .B(cell_2054_and_out[0]), .Z(
        signal_2322) );
  XOR2_X1 cell_2054_U2 ( .A(signal_3666), .B(signal_3744), .Z(
        cell_2054_and_in[1]) );
  XOR2_X1 cell_2054_U1 ( .A(signal_2156), .B(signal_2234), .Z(
        cell_2054_and_in[0]) );
  XOR2_X1 cell_2054_a_HPC2_and_U14 ( .A(Fresh[340]), .B(cell_2054_and_in[0]), 
        .Z(cell_2054_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2054_a_HPC2_and_U13 ( .A(Fresh[340]), .B(cell_2054_and_in[1]), 
        .Z(cell_2054_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2054_a_HPC2_and_U12 ( .A1(cell_2054_a_HPC2_and_a_reg[1]), .A2(
        cell_2054_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2054_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2054_a_HPC2_and_U11 ( .A1(cell_2054_a_HPC2_and_a_reg[0]), .A2(
        cell_2054_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2054_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2054_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2054_a_HPC2_and_n9), 
        .ZN(cell_2054_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2054_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2054_a_HPC2_and_n9), 
        .ZN(cell_2054_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2054_a_HPC2_and_U8 ( .A(Fresh[340]), .ZN(cell_2054_a_HPC2_and_n9) );
  AND2_X1 cell_2054_a_HPC2_and_U7 ( .A1(cell_2054_and_in[1]), .A2(n468), .ZN(
        cell_2054_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2054_a_HPC2_and_U6 ( .A1(cell_2054_and_in[0]), .A2(n464), .ZN(
        cell_2054_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2054_a_HPC2_and_U5 ( .A(cell_2054_a_HPC2_and_n8), .B(
        cell_2054_a_HPC2_and_z_1__1_), .ZN(cell_2054_and_out[1]) );
  XNOR2_X1 cell_2054_a_HPC2_and_U4 ( .A(
        cell_2054_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2054_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2054_a_HPC2_and_n8) );
  XNOR2_X1 cell_2054_a_HPC2_and_U3 ( .A(cell_2054_a_HPC2_and_n7), .B(
        cell_2054_a_HPC2_and_z_0__0_), .ZN(cell_2054_and_out[0]) );
  XNOR2_X1 cell_2054_a_HPC2_and_U2 ( .A(
        cell_2054_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2054_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2054_a_HPC2_and_n7) );
  DFF_X1 cell_2054_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2054_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2054_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2054_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2054_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2054_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2054_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2054_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2054_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2054_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2055_U4 ( .A(signal_3713), .B(cell_2055_and_out[1]), .Z(
        signal_3969) );
  XOR2_X1 cell_2055_U3 ( .A(signal_2203), .B(cell_2055_and_out[0]), .Z(
        signal_2323) );
  XOR2_X1 cell_2055_U2 ( .A(signal_3713), .B(signal_3702), .Z(
        cell_2055_and_in[1]) );
  XOR2_X1 cell_2055_U1 ( .A(signal_2203), .B(signal_2192), .Z(
        cell_2055_and_in[0]) );
  XOR2_X1 cell_2055_a_HPC2_and_U14 ( .A(Fresh[341]), .B(cell_2055_and_in[0]), 
        .Z(cell_2055_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2055_a_HPC2_and_U13 ( .A(Fresh[341]), .B(cell_2055_and_in[1]), 
        .Z(cell_2055_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2055_a_HPC2_and_U12 ( .A1(cell_2055_a_HPC2_and_a_reg[1]), .A2(
        cell_2055_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2055_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2055_a_HPC2_and_U11 ( .A1(cell_2055_a_HPC2_and_a_reg[0]), .A2(
        cell_2055_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2055_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2055_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2055_a_HPC2_and_n9), 
        .ZN(cell_2055_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2055_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2055_a_HPC2_and_n9), 
        .ZN(cell_2055_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2055_a_HPC2_and_U8 ( .A(Fresh[341]), .ZN(cell_2055_a_HPC2_and_n9) );
  AND2_X1 cell_2055_a_HPC2_and_U7 ( .A1(cell_2055_and_in[1]), .A2(n468), .ZN(
        cell_2055_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2055_a_HPC2_and_U6 ( .A1(cell_2055_and_in[0]), .A2(n464), .ZN(
        cell_2055_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2055_a_HPC2_and_U5 ( .A(cell_2055_a_HPC2_and_n8), .B(
        cell_2055_a_HPC2_and_z_1__1_), .ZN(cell_2055_and_out[1]) );
  XNOR2_X1 cell_2055_a_HPC2_and_U4 ( .A(
        cell_2055_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2055_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2055_a_HPC2_and_n8) );
  XNOR2_X1 cell_2055_a_HPC2_and_U3 ( .A(cell_2055_a_HPC2_and_n7), .B(
        cell_2055_a_HPC2_and_z_0__0_), .ZN(cell_2055_and_out[0]) );
  XNOR2_X1 cell_2055_a_HPC2_and_U2 ( .A(
        cell_2055_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2055_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2055_a_HPC2_and_n7) );
  DFF_X1 cell_2055_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2055_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2055_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2055_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2055_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2055_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2055_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2055_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2055_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2055_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2056_U4 ( .A(signal_3673), .B(cell_2056_and_out[1]), .Z(
        signal_3970) );
  XOR2_X1 cell_2056_U3 ( .A(signal_2163), .B(cell_2056_and_out[0]), .Z(
        signal_2324) );
  XOR2_X1 cell_2056_U2 ( .A(signal_3673), .B(signal_3721), .Z(
        cell_2056_and_in[1]) );
  XOR2_X1 cell_2056_U1 ( .A(signal_2163), .B(signal_2211), .Z(
        cell_2056_and_in[0]) );
  XOR2_X1 cell_2056_a_HPC2_and_U14 ( .A(Fresh[342]), .B(cell_2056_and_in[0]), 
        .Z(cell_2056_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2056_a_HPC2_and_U13 ( .A(Fresh[342]), .B(cell_2056_and_in[1]), 
        .Z(cell_2056_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2056_a_HPC2_and_U12 ( .A1(cell_2056_a_HPC2_and_a_reg[1]), .A2(
        cell_2056_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2056_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2056_a_HPC2_and_U11 ( .A1(cell_2056_a_HPC2_and_a_reg[0]), .A2(
        cell_2056_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2056_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2056_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2056_a_HPC2_and_n9), 
        .ZN(cell_2056_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2056_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2056_a_HPC2_and_n9), 
        .ZN(cell_2056_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2056_a_HPC2_and_U8 ( .A(Fresh[342]), .ZN(cell_2056_a_HPC2_and_n9) );
  AND2_X1 cell_2056_a_HPC2_and_U7 ( .A1(cell_2056_and_in[1]), .A2(n469), .ZN(
        cell_2056_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2056_a_HPC2_and_U6 ( .A1(cell_2056_and_in[0]), .A2(n465), .ZN(
        cell_2056_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2056_a_HPC2_and_U5 ( .A(cell_2056_a_HPC2_and_n8), .B(
        cell_2056_a_HPC2_and_z_1__1_), .ZN(cell_2056_and_out[1]) );
  XNOR2_X1 cell_2056_a_HPC2_and_U4 ( .A(
        cell_2056_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2056_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2056_a_HPC2_and_n8) );
  XNOR2_X1 cell_2056_a_HPC2_and_U3 ( .A(cell_2056_a_HPC2_and_n7), .B(
        cell_2056_a_HPC2_and_z_0__0_), .ZN(cell_2056_and_out[0]) );
  XNOR2_X1 cell_2056_a_HPC2_and_U2 ( .A(
        cell_2056_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2056_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2056_a_HPC2_and_n7) );
  DFF_X1 cell_2056_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2056_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2056_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2056_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2056_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2056_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2056_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2056_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2056_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2056_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2057_U4 ( .A(signal_3689), .B(cell_2057_and_out[1]), .Z(
        signal_3971) );
  XOR2_X1 cell_2057_U3 ( .A(signal_2179), .B(cell_2057_and_out[0]), .Z(
        signal_2325) );
  XOR2_X1 cell_2057_U2 ( .A(signal_3689), .B(signal_3687), .Z(
        cell_2057_and_in[1]) );
  XOR2_X1 cell_2057_U1 ( .A(signal_2179), .B(signal_2177), .Z(
        cell_2057_and_in[0]) );
  XOR2_X1 cell_2057_a_HPC2_and_U14 ( .A(Fresh[343]), .B(cell_2057_and_in[0]), 
        .Z(cell_2057_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2057_a_HPC2_and_U13 ( .A(Fresh[343]), .B(cell_2057_and_in[1]), 
        .Z(cell_2057_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2057_a_HPC2_and_U12 ( .A1(cell_2057_a_HPC2_and_a_reg[1]), .A2(
        cell_2057_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2057_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2057_a_HPC2_and_U11 ( .A1(cell_2057_a_HPC2_and_a_reg[0]), .A2(
        cell_2057_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2057_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2057_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2057_a_HPC2_and_n9), 
        .ZN(cell_2057_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2057_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2057_a_HPC2_and_n9), 
        .ZN(cell_2057_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2057_a_HPC2_and_U8 ( .A(Fresh[343]), .ZN(cell_2057_a_HPC2_and_n9) );
  AND2_X1 cell_2057_a_HPC2_and_U7 ( .A1(cell_2057_and_in[1]), .A2(n469), .ZN(
        cell_2057_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2057_a_HPC2_and_U6 ( .A1(cell_2057_and_in[0]), .A2(n465), .ZN(
        cell_2057_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2057_a_HPC2_and_U5 ( .A(cell_2057_a_HPC2_and_n8), .B(
        cell_2057_a_HPC2_and_z_1__1_), .ZN(cell_2057_and_out[1]) );
  XNOR2_X1 cell_2057_a_HPC2_and_U4 ( .A(
        cell_2057_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2057_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2057_a_HPC2_and_n8) );
  XNOR2_X1 cell_2057_a_HPC2_and_U3 ( .A(cell_2057_a_HPC2_and_n7), .B(
        cell_2057_a_HPC2_and_z_0__0_), .ZN(cell_2057_and_out[0]) );
  XNOR2_X1 cell_2057_a_HPC2_and_U2 ( .A(
        cell_2057_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2057_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2057_a_HPC2_and_n7) );
  DFF_X1 cell_2057_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2057_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2057_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2057_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2057_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2057_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2057_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2057_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2057_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2057_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2058_U4 ( .A(signal_3675), .B(cell_2058_and_out[1]), .Z(
        signal_3972) );
  XOR2_X1 cell_2058_U3 ( .A(signal_2165), .B(cell_2058_and_out[0]), .Z(
        signal_2326) );
  XOR2_X1 cell_2058_U2 ( .A(signal_3675), .B(signal_3761), .Z(
        cell_2058_and_in[1]) );
  XOR2_X1 cell_2058_U1 ( .A(signal_2165), .B(signal_2251), .Z(
        cell_2058_and_in[0]) );
  XOR2_X1 cell_2058_a_HPC2_and_U14 ( .A(Fresh[344]), .B(cell_2058_and_in[0]), 
        .Z(cell_2058_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2058_a_HPC2_and_U13 ( .A(Fresh[344]), .B(cell_2058_and_in[1]), 
        .Z(cell_2058_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2058_a_HPC2_and_U12 ( .A1(cell_2058_a_HPC2_and_a_reg[1]), .A2(
        cell_2058_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2058_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2058_a_HPC2_and_U11 ( .A1(cell_2058_a_HPC2_and_a_reg[0]), .A2(
        cell_2058_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2058_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2058_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2058_a_HPC2_and_n9), 
        .ZN(cell_2058_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2058_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2058_a_HPC2_and_n9), 
        .ZN(cell_2058_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2058_a_HPC2_and_U8 ( .A(Fresh[344]), .ZN(cell_2058_a_HPC2_and_n9) );
  AND2_X1 cell_2058_a_HPC2_and_U7 ( .A1(cell_2058_and_in[1]), .A2(n469), .ZN(
        cell_2058_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2058_a_HPC2_and_U6 ( .A1(cell_2058_and_in[0]), .A2(n465), .ZN(
        cell_2058_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2058_a_HPC2_and_U5 ( .A(cell_2058_a_HPC2_and_n8), .B(
        cell_2058_a_HPC2_and_z_1__1_), .ZN(cell_2058_and_out[1]) );
  XNOR2_X1 cell_2058_a_HPC2_and_U4 ( .A(
        cell_2058_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2058_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2058_a_HPC2_and_n8) );
  XNOR2_X1 cell_2058_a_HPC2_and_U3 ( .A(cell_2058_a_HPC2_and_n7), .B(
        cell_2058_a_HPC2_and_z_0__0_), .ZN(cell_2058_and_out[0]) );
  XNOR2_X1 cell_2058_a_HPC2_and_U2 ( .A(
        cell_2058_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2058_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2058_a_HPC2_and_n7) );
  DFF_X1 cell_2058_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2058_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2058_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2058_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2058_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2058_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2058_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2058_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2058_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2058_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2059_U4 ( .A(signal_3728), .B(cell_2059_and_out[1]), .Z(
        signal_3973) );
  XOR2_X1 cell_2059_U3 ( .A(signal_2218), .B(cell_2059_and_out[0]), .Z(
        signal_2327) );
  XOR2_X1 cell_2059_U2 ( .A(signal_3728), .B(signal_3735), .Z(
        cell_2059_and_in[1]) );
  XOR2_X1 cell_2059_U1 ( .A(signal_2218), .B(signal_2225), .Z(
        cell_2059_and_in[0]) );
  XOR2_X1 cell_2059_a_HPC2_and_U14 ( .A(Fresh[345]), .B(cell_2059_and_in[0]), 
        .Z(cell_2059_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2059_a_HPC2_and_U13 ( .A(Fresh[345]), .B(cell_2059_and_in[1]), 
        .Z(cell_2059_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2059_a_HPC2_and_U12 ( .A1(cell_2059_a_HPC2_and_a_reg[1]), .A2(
        cell_2059_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2059_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2059_a_HPC2_and_U11 ( .A1(cell_2059_a_HPC2_and_a_reg[0]), .A2(
        cell_2059_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2059_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2059_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2059_a_HPC2_and_n9), 
        .ZN(cell_2059_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2059_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2059_a_HPC2_and_n9), 
        .ZN(cell_2059_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2059_a_HPC2_and_U8 ( .A(Fresh[345]), .ZN(cell_2059_a_HPC2_and_n9) );
  AND2_X1 cell_2059_a_HPC2_and_U7 ( .A1(cell_2059_and_in[1]), .A2(n469), .ZN(
        cell_2059_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2059_a_HPC2_and_U6 ( .A1(cell_2059_and_in[0]), .A2(n465), .ZN(
        cell_2059_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2059_a_HPC2_and_U5 ( .A(cell_2059_a_HPC2_and_n8), .B(
        cell_2059_a_HPC2_and_z_1__1_), .ZN(cell_2059_and_out[1]) );
  XNOR2_X1 cell_2059_a_HPC2_and_U4 ( .A(
        cell_2059_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2059_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2059_a_HPC2_and_n8) );
  XNOR2_X1 cell_2059_a_HPC2_and_U3 ( .A(cell_2059_a_HPC2_and_n7), .B(
        cell_2059_a_HPC2_and_z_0__0_), .ZN(cell_2059_and_out[0]) );
  XNOR2_X1 cell_2059_a_HPC2_and_U2 ( .A(
        cell_2059_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2059_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2059_a_HPC2_and_n7) );
  DFF_X1 cell_2059_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2059_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2059_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2059_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2059_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2059_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2059_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2059_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2059_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2059_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2060_U4 ( .A(signal_3758), .B(cell_2060_and_out[1]), .Z(
        signal_3974) );
  XOR2_X1 cell_2060_U3 ( .A(signal_2248), .B(cell_2060_and_out[0]), .Z(
        signal_2328) );
  XOR2_X1 cell_2060_U2 ( .A(signal_3758), .B(signal_3767), .Z(
        cell_2060_and_in[1]) );
  XOR2_X1 cell_2060_U1 ( .A(signal_2248), .B(signal_2257), .Z(
        cell_2060_and_in[0]) );
  XOR2_X1 cell_2060_a_HPC2_and_U14 ( .A(Fresh[346]), .B(cell_2060_and_in[0]), 
        .Z(cell_2060_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2060_a_HPC2_and_U13 ( .A(Fresh[346]), .B(cell_2060_and_in[1]), 
        .Z(cell_2060_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2060_a_HPC2_and_U12 ( .A1(cell_2060_a_HPC2_and_a_reg[1]), .A2(
        cell_2060_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2060_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2060_a_HPC2_and_U11 ( .A1(cell_2060_a_HPC2_and_a_reg[0]), .A2(
        cell_2060_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2060_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2060_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2060_a_HPC2_and_n9), 
        .ZN(cell_2060_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2060_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2060_a_HPC2_and_n9), 
        .ZN(cell_2060_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2060_a_HPC2_and_U8 ( .A(Fresh[346]), .ZN(cell_2060_a_HPC2_and_n9) );
  AND2_X1 cell_2060_a_HPC2_and_U7 ( .A1(cell_2060_and_in[1]), .A2(n469), .ZN(
        cell_2060_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2060_a_HPC2_and_U6 ( .A1(cell_2060_and_in[0]), .A2(n465), .ZN(
        cell_2060_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2060_a_HPC2_and_U5 ( .A(cell_2060_a_HPC2_and_n8), .B(
        cell_2060_a_HPC2_and_z_1__1_), .ZN(cell_2060_and_out[1]) );
  XNOR2_X1 cell_2060_a_HPC2_and_U4 ( .A(
        cell_2060_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2060_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2060_a_HPC2_and_n8) );
  XNOR2_X1 cell_2060_a_HPC2_and_U3 ( .A(cell_2060_a_HPC2_and_n7), .B(
        cell_2060_a_HPC2_and_z_0__0_), .ZN(cell_2060_and_out[0]) );
  XNOR2_X1 cell_2060_a_HPC2_and_U2 ( .A(
        cell_2060_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2060_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2060_a_HPC2_and_n7) );
  DFF_X1 cell_2060_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2060_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2060_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2060_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2060_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2060_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2060_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2060_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2060_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2060_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2061_U4 ( .A(signal_3518), .B(cell_2061_and_out[1]), .Z(
        signal_3975) );
  XOR2_X1 cell_2061_U3 ( .A(signal_2080), .B(cell_2061_and_out[0]), .Z(
        signal_2329) );
  XOR2_X1 cell_2061_U2 ( .A(signal_3518), .B(signal_3738), .Z(
        cell_2061_and_in[1]) );
  XOR2_X1 cell_2061_U1 ( .A(signal_2080), .B(signal_2228), .Z(
        cell_2061_and_in[0]) );
  XOR2_X1 cell_2061_a_HPC2_and_U14 ( .A(Fresh[347]), .B(cell_2061_and_in[0]), 
        .Z(cell_2061_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2061_a_HPC2_and_U13 ( .A(Fresh[347]), .B(cell_2061_and_in[1]), 
        .Z(cell_2061_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2061_a_HPC2_and_U12 ( .A1(cell_2061_a_HPC2_and_a_reg[1]), .A2(
        cell_2061_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2061_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2061_a_HPC2_and_U11 ( .A1(cell_2061_a_HPC2_and_a_reg[0]), .A2(
        cell_2061_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2061_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2061_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2061_a_HPC2_and_n9), 
        .ZN(cell_2061_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2061_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2061_a_HPC2_and_n9), 
        .ZN(cell_2061_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2061_a_HPC2_and_U8 ( .A(Fresh[347]), .ZN(cell_2061_a_HPC2_and_n9) );
  AND2_X1 cell_2061_a_HPC2_and_U7 ( .A1(cell_2061_and_in[1]), .A2(n469), .ZN(
        cell_2061_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2061_a_HPC2_and_U6 ( .A1(cell_2061_and_in[0]), .A2(n465), .ZN(
        cell_2061_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2061_a_HPC2_and_U5 ( .A(cell_2061_a_HPC2_and_n8), .B(
        cell_2061_a_HPC2_and_z_1__1_), .ZN(cell_2061_and_out[1]) );
  XNOR2_X1 cell_2061_a_HPC2_and_U4 ( .A(
        cell_2061_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2061_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2061_a_HPC2_and_n8) );
  XNOR2_X1 cell_2061_a_HPC2_and_U3 ( .A(cell_2061_a_HPC2_and_n7), .B(
        cell_2061_a_HPC2_and_z_0__0_), .ZN(cell_2061_and_out[0]) );
  XNOR2_X1 cell_2061_a_HPC2_and_U2 ( .A(
        cell_2061_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2061_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2061_a_HPC2_and_n7) );
  DFF_X1 cell_2061_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2061_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2061_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2061_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2061_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2061_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2061_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2061_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2061_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2061_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2062_U4 ( .A(signal_3693), .B(cell_2062_and_out[1]), .Z(
        signal_3976) );
  XOR2_X1 cell_2062_U3 ( .A(signal_2183), .B(cell_2062_and_out[0]), .Z(
        signal_2330) );
  XOR2_X1 cell_2062_U2 ( .A(signal_3693), .B(signal_3773), .Z(
        cell_2062_and_in[1]) );
  XOR2_X1 cell_2062_U1 ( .A(signal_2183), .B(signal_2263), .Z(
        cell_2062_and_in[0]) );
  XOR2_X1 cell_2062_a_HPC2_and_U14 ( .A(Fresh[348]), .B(cell_2062_and_in[0]), 
        .Z(cell_2062_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2062_a_HPC2_and_U13 ( .A(Fresh[348]), .B(cell_2062_and_in[1]), 
        .Z(cell_2062_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2062_a_HPC2_and_U12 ( .A1(cell_2062_a_HPC2_and_a_reg[1]), .A2(
        cell_2062_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2062_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2062_a_HPC2_and_U11 ( .A1(cell_2062_a_HPC2_and_a_reg[0]), .A2(
        cell_2062_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2062_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2062_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2062_a_HPC2_and_n9), 
        .ZN(cell_2062_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2062_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2062_a_HPC2_and_n9), 
        .ZN(cell_2062_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2062_a_HPC2_and_U8 ( .A(Fresh[348]), .ZN(cell_2062_a_HPC2_and_n9) );
  AND2_X1 cell_2062_a_HPC2_and_U7 ( .A1(cell_2062_and_in[1]), .A2(n469), .ZN(
        cell_2062_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2062_a_HPC2_and_U6 ( .A1(cell_2062_and_in[0]), .A2(n465), .ZN(
        cell_2062_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2062_a_HPC2_and_U5 ( .A(cell_2062_a_HPC2_and_n8), .B(
        cell_2062_a_HPC2_and_z_1__1_), .ZN(cell_2062_and_out[1]) );
  XNOR2_X1 cell_2062_a_HPC2_and_U4 ( .A(
        cell_2062_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2062_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2062_a_HPC2_and_n8) );
  XNOR2_X1 cell_2062_a_HPC2_and_U3 ( .A(cell_2062_a_HPC2_and_n7), .B(
        cell_2062_a_HPC2_and_z_0__0_), .ZN(cell_2062_and_out[0]) );
  XNOR2_X1 cell_2062_a_HPC2_and_U2 ( .A(
        cell_2062_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2062_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2062_a_HPC2_and_n7) );
  DFF_X1 cell_2062_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2062_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2062_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2062_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2062_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2062_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2062_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2062_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2062_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2062_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2063_U4 ( .A(signal_3690), .B(cell_2063_and_out[1]), .Z(
        signal_3977) );
  XOR2_X1 cell_2063_U3 ( .A(signal_2180), .B(cell_2063_and_out[0]), .Z(
        signal_2331) );
  XOR2_X1 cell_2063_U2 ( .A(signal_3690), .B(signal_3679), .Z(
        cell_2063_and_in[1]) );
  XOR2_X1 cell_2063_U1 ( .A(signal_2180), .B(signal_2169), .Z(
        cell_2063_and_in[0]) );
  XOR2_X1 cell_2063_a_HPC2_and_U14 ( .A(Fresh[349]), .B(cell_2063_and_in[0]), 
        .Z(cell_2063_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2063_a_HPC2_and_U13 ( .A(Fresh[349]), .B(cell_2063_and_in[1]), 
        .Z(cell_2063_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2063_a_HPC2_and_U12 ( .A1(cell_2063_a_HPC2_and_a_reg[1]), .A2(
        cell_2063_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2063_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2063_a_HPC2_and_U11 ( .A1(cell_2063_a_HPC2_and_a_reg[0]), .A2(
        cell_2063_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2063_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2063_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2063_a_HPC2_and_n9), 
        .ZN(cell_2063_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2063_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2063_a_HPC2_and_n9), 
        .ZN(cell_2063_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2063_a_HPC2_and_U8 ( .A(Fresh[349]), .ZN(cell_2063_a_HPC2_and_n9) );
  AND2_X1 cell_2063_a_HPC2_and_U7 ( .A1(cell_2063_and_in[1]), .A2(n469), .ZN(
        cell_2063_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2063_a_HPC2_and_U6 ( .A1(cell_2063_and_in[0]), .A2(n465), .ZN(
        cell_2063_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2063_a_HPC2_and_U5 ( .A(cell_2063_a_HPC2_and_n8), .B(
        cell_2063_a_HPC2_and_z_1__1_), .ZN(cell_2063_and_out[1]) );
  XNOR2_X1 cell_2063_a_HPC2_and_U4 ( .A(
        cell_2063_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2063_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2063_a_HPC2_and_n8) );
  XNOR2_X1 cell_2063_a_HPC2_and_U3 ( .A(cell_2063_a_HPC2_and_n7), .B(
        cell_2063_a_HPC2_and_z_0__0_), .ZN(cell_2063_and_out[0]) );
  XNOR2_X1 cell_2063_a_HPC2_and_U2 ( .A(
        cell_2063_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2063_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2063_a_HPC2_and_n7) );
  DFF_X1 cell_2063_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2063_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2063_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2063_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2063_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2063_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2063_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2063_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2063_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2063_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2064_U4 ( .A(signal_3782), .B(cell_2064_and_out[1]), .Z(
        signal_3978) );
  XOR2_X1 cell_2064_U3 ( .A(signal_2272), .B(cell_2064_and_out[0]), .Z(
        signal_2332) );
  XOR2_X1 cell_2064_U2 ( .A(signal_3782), .B(signal_3763), .Z(
        cell_2064_and_in[1]) );
  XOR2_X1 cell_2064_U1 ( .A(signal_2272), .B(signal_2253), .Z(
        cell_2064_and_in[0]) );
  XOR2_X1 cell_2064_a_HPC2_and_U14 ( .A(Fresh[350]), .B(cell_2064_and_in[0]), 
        .Z(cell_2064_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2064_a_HPC2_and_U13 ( .A(Fresh[350]), .B(cell_2064_and_in[1]), 
        .Z(cell_2064_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2064_a_HPC2_and_U12 ( .A1(cell_2064_a_HPC2_and_a_reg[1]), .A2(
        cell_2064_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2064_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2064_a_HPC2_and_U11 ( .A1(cell_2064_a_HPC2_and_a_reg[0]), .A2(
        cell_2064_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2064_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2064_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2064_a_HPC2_and_n9), 
        .ZN(cell_2064_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2064_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2064_a_HPC2_and_n9), 
        .ZN(cell_2064_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2064_a_HPC2_and_U8 ( .A(Fresh[350]), .ZN(cell_2064_a_HPC2_and_n9) );
  AND2_X1 cell_2064_a_HPC2_and_U7 ( .A1(cell_2064_and_in[1]), .A2(n469), .ZN(
        cell_2064_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2064_a_HPC2_and_U6 ( .A1(cell_2064_and_in[0]), .A2(n465), .ZN(
        cell_2064_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2064_a_HPC2_and_U5 ( .A(cell_2064_a_HPC2_and_n8), .B(
        cell_2064_a_HPC2_and_z_1__1_), .ZN(cell_2064_and_out[1]) );
  XNOR2_X1 cell_2064_a_HPC2_and_U4 ( .A(
        cell_2064_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2064_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2064_a_HPC2_and_n8) );
  XNOR2_X1 cell_2064_a_HPC2_and_U3 ( .A(cell_2064_a_HPC2_and_n7), .B(
        cell_2064_a_HPC2_and_z_0__0_), .ZN(cell_2064_and_out[0]) );
  XNOR2_X1 cell_2064_a_HPC2_and_U2 ( .A(
        cell_2064_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2064_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2064_a_HPC2_and_n7) );
  DFF_X1 cell_2064_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2064_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2064_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2064_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2064_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2064_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2064_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2064_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2064_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2064_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2065_U4 ( .A(signal_3777), .B(cell_2065_and_out[1]), .Z(
        signal_3979) );
  XOR2_X1 cell_2065_U3 ( .A(signal_2267), .B(cell_2065_and_out[0]), .Z(
        signal_2333) );
  XOR2_X1 cell_2065_U2 ( .A(signal_3777), .B(signal_3749), .Z(
        cell_2065_and_in[1]) );
  XOR2_X1 cell_2065_U1 ( .A(signal_2267), .B(signal_2239), .Z(
        cell_2065_and_in[0]) );
  XOR2_X1 cell_2065_a_HPC2_and_U14 ( .A(Fresh[351]), .B(cell_2065_and_in[0]), 
        .Z(cell_2065_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2065_a_HPC2_and_U13 ( .A(Fresh[351]), .B(cell_2065_and_in[1]), 
        .Z(cell_2065_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2065_a_HPC2_and_U12 ( .A1(cell_2065_a_HPC2_and_a_reg[1]), .A2(
        cell_2065_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2065_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2065_a_HPC2_and_U11 ( .A1(cell_2065_a_HPC2_and_a_reg[0]), .A2(
        cell_2065_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2065_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2065_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2065_a_HPC2_and_n9), 
        .ZN(cell_2065_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2065_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2065_a_HPC2_and_n9), 
        .ZN(cell_2065_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2065_a_HPC2_and_U8 ( .A(Fresh[351]), .ZN(cell_2065_a_HPC2_and_n9) );
  AND2_X1 cell_2065_a_HPC2_and_U7 ( .A1(cell_2065_and_in[1]), .A2(n469), .ZN(
        cell_2065_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2065_a_HPC2_and_U6 ( .A1(cell_2065_and_in[0]), .A2(n465), .ZN(
        cell_2065_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2065_a_HPC2_and_U5 ( .A(cell_2065_a_HPC2_and_n8), .B(
        cell_2065_a_HPC2_and_z_1__1_), .ZN(cell_2065_and_out[1]) );
  XNOR2_X1 cell_2065_a_HPC2_and_U4 ( .A(
        cell_2065_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2065_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2065_a_HPC2_and_n8) );
  XNOR2_X1 cell_2065_a_HPC2_and_U3 ( .A(cell_2065_a_HPC2_and_n7), .B(
        cell_2065_a_HPC2_and_z_0__0_), .ZN(cell_2065_and_out[0]) );
  XNOR2_X1 cell_2065_a_HPC2_and_U2 ( .A(
        cell_2065_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2065_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2065_a_HPC2_and_n7) );
  DFF_X1 cell_2065_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2065_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2065_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2065_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2065_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2065_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2065_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2065_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2065_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2065_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2066_U4 ( .A(signal_3559), .B(cell_2066_and_out[1]), .Z(
        signal_3980) );
  XOR2_X1 cell_2066_U3 ( .A(signal_2121), .B(cell_2066_and_out[0]), .Z(
        signal_2334) );
  XOR2_X1 cell_2066_U2 ( .A(signal_3559), .B(signal_3756), .Z(
        cell_2066_and_in[1]) );
  XOR2_X1 cell_2066_U1 ( .A(signal_2121), .B(signal_2246), .Z(
        cell_2066_and_in[0]) );
  XOR2_X1 cell_2066_a_HPC2_and_U14 ( .A(Fresh[352]), .B(cell_2066_and_in[0]), 
        .Z(cell_2066_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2066_a_HPC2_and_U13 ( .A(Fresh[352]), .B(cell_2066_and_in[1]), 
        .Z(cell_2066_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2066_a_HPC2_and_U12 ( .A1(cell_2066_a_HPC2_and_a_reg[1]), .A2(
        cell_2066_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2066_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2066_a_HPC2_and_U11 ( .A1(cell_2066_a_HPC2_and_a_reg[0]), .A2(
        cell_2066_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2066_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2066_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2066_a_HPC2_and_n9), 
        .ZN(cell_2066_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2066_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2066_a_HPC2_and_n9), 
        .ZN(cell_2066_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2066_a_HPC2_and_U8 ( .A(Fresh[352]), .ZN(cell_2066_a_HPC2_and_n9) );
  AND2_X1 cell_2066_a_HPC2_and_U7 ( .A1(cell_2066_and_in[1]), .A2(n469), .ZN(
        cell_2066_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2066_a_HPC2_and_U6 ( .A1(cell_2066_and_in[0]), .A2(n465), .ZN(
        cell_2066_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2066_a_HPC2_and_U5 ( .A(cell_2066_a_HPC2_and_n8), .B(
        cell_2066_a_HPC2_and_z_1__1_), .ZN(cell_2066_and_out[1]) );
  XNOR2_X1 cell_2066_a_HPC2_and_U4 ( .A(
        cell_2066_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2066_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2066_a_HPC2_and_n8) );
  XNOR2_X1 cell_2066_a_HPC2_and_U3 ( .A(cell_2066_a_HPC2_and_n7), .B(
        cell_2066_a_HPC2_and_z_0__0_), .ZN(cell_2066_and_out[0]) );
  XNOR2_X1 cell_2066_a_HPC2_and_U2 ( .A(
        cell_2066_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2066_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2066_a_HPC2_and_n7) );
  DFF_X1 cell_2066_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2066_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2066_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2066_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2066_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2066_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2066_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2066_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2066_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2066_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2067_U4 ( .A(signal_3701), .B(cell_2067_and_out[1]), .Z(
        signal_3981) );
  XOR2_X1 cell_2067_U3 ( .A(signal_2191), .B(cell_2067_and_out[0]), .Z(
        signal_2335) );
  XOR2_X1 cell_2067_U2 ( .A(signal_3701), .B(signal_3709), .Z(
        cell_2067_and_in[1]) );
  XOR2_X1 cell_2067_U1 ( .A(signal_2191), .B(signal_2199), .Z(
        cell_2067_and_in[0]) );
  XOR2_X1 cell_2067_a_HPC2_and_U14 ( .A(Fresh[353]), .B(cell_2067_and_in[0]), 
        .Z(cell_2067_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2067_a_HPC2_and_U13 ( .A(Fresh[353]), .B(cell_2067_and_in[1]), 
        .Z(cell_2067_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2067_a_HPC2_and_U12 ( .A1(cell_2067_a_HPC2_and_a_reg[1]), .A2(
        cell_2067_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2067_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2067_a_HPC2_and_U11 ( .A1(cell_2067_a_HPC2_and_a_reg[0]), .A2(
        cell_2067_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2067_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2067_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2067_a_HPC2_and_n9), 
        .ZN(cell_2067_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2067_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2067_a_HPC2_and_n9), 
        .ZN(cell_2067_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2067_a_HPC2_and_U8 ( .A(Fresh[353]), .ZN(cell_2067_a_HPC2_and_n9) );
  AND2_X1 cell_2067_a_HPC2_and_U7 ( .A1(cell_2067_and_in[1]), .A2(n469), .ZN(
        cell_2067_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2067_a_HPC2_and_U6 ( .A1(cell_2067_and_in[0]), .A2(n465), .ZN(
        cell_2067_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2067_a_HPC2_and_U5 ( .A(cell_2067_a_HPC2_and_n8), .B(
        cell_2067_a_HPC2_and_z_1__1_), .ZN(cell_2067_and_out[1]) );
  XNOR2_X1 cell_2067_a_HPC2_and_U4 ( .A(
        cell_2067_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2067_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2067_a_HPC2_and_n8) );
  XNOR2_X1 cell_2067_a_HPC2_and_U3 ( .A(cell_2067_a_HPC2_and_n7), .B(
        cell_2067_a_HPC2_and_z_0__0_), .ZN(cell_2067_and_out[0]) );
  XNOR2_X1 cell_2067_a_HPC2_and_U2 ( .A(
        cell_2067_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2067_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2067_a_HPC2_and_n7) );
  DFF_X1 cell_2067_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2067_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2067_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2067_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2067_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2067_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2067_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2067_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2067_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2067_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2068_U4 ( .A(signal_3688), .B(cell_2068_and_out[1]), .Z(
        signal_3982) );
  XOR2_X1 cell_2068_U3 ( .A(signal_2178), .B(cell_2068_and_out[0]), .Z(
        signal_2336) );
  XOR2_X1 cell_2068_U2 ( .A(signal_3688), .B(signal_3670), .Z(
        cell_2068_and_in[1]) );
  XOR2_X1 cell_2068_U1 ( .A(signal_2178), .B(signal_2160), .Z(
        cell_2068_and_in[0]) );
  XOR2_X1 cell_2068_a_HPC2_and_U14 ( .A(Fresh[354]), .B(cell_2068_and_in[0]), 
        .Z(cell_2068_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2068_a_HPC2_and_U13 ( .A(Fresh[354]), .B(cell_2068_and_in[1]), 
        .Z(cell_2068_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2068_a_HPC2_and_U12 ( .A1(cell_2068_a_HPC2_and_a_reg[1]), .A2(
        cell_2068_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2068_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2068_a_HPC2_and_U11 ( .A1(cell_2068_a_HPC2_and_a_reg[0]), .A2(
        cell_2068_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2068_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2068_a_HPC2_and_U10 ( .A1(n467), .A2(cell_2068_a_HPC2_and_n9), 
        .ZN(cell_2068_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2068_a_HPC2_and_U9 ( .A1(n463), .A2(cell_2068_a_HPC2_and_n9), 
        .ZN(cell_2068_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2068_a_HPC2_and_U8 ( .A(Fresh[354]), .ZN(cell_2068_a_HPC2_and_n9) );
  AND2_X1 cell_2068_a_HPC2_and_U7 ( .A1(cell_2068_and_in[1]), .A2(n467), .ZN(
        cell_2068_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2068_a_HPC2_and_U6 ( .A1(cell_2068_and_in[0]), .A2(n463), .ZN(
        cell_2068_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2068_a_HPC2_and_U5 ( .A(cell_2068_a_HPC2_and_n8), .B(
        cell_2068_a_HPC2_and_z_1__1_), .ZN(cell_2068_and_out[1]) );
  XNOR2_X1 cell_2068_a_HPC2_and_U4 ( .A(
        cell_2068_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2068_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2068_a_HPC2_and_n8) );
  XNOR2_X1 cell_2068_a_HPC2_and_U3 ( .A(cell_2068_a_HPC2_and_n7), .B(
        cell_2068_a_HPC2_and_z_0__0_), .ZN(cell_2068_and_out[0]) );
  XNOR2_X1 cell_2068_a_HPC2_and_U2 ( .A(
        cell_2068_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2068_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2068_a_HPC2_and_n7) );
  DFF_X1 cell_2068_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2068_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2068_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n463), .CK(clk), 
        .Q(cell_2068_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2068_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2068_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n467), .CK(clk), 
        .Q(cell_2068_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2068_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2068_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2068_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2069_U4 ( .A(signal_3716), .B(cell_2069_and_out[1]), .Z(
        signal_3983) );
  XOR2_X1 cell_2069_U3 ( .A(signal_2206), .B(cell_2069_and_out[0]), .Z(
        signal_2337) );
  XOR2_X1 cell_2069_U2 ( .A(signal_3716), .B(signal_3698), .Z(
        cell_2069_and_in[1]) );
  XOR2_X1 cell_2069_U1 ( .A(signal_2206), .B(signal_2188), .Z(
        cell_2069_and_in[0]) );
  XOR2_X1 cell_2069_a_HPC2_and_U14 ( .A(Fresh[355]), .B(cell_2069_and_in[0]), 
        .Z(cell_2069_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2069_a_HPC2_and_U13 ( .A(Fresh[355]), .B(cell_2069_and_in[1]), 
        .Z(cell_2069_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2069_a_HPC2_and_U12 ( .A1(cell_2069_a_HPC2_and_a_reg[1]), .A2(
        cell_2069_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2069_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2069_a_HPC2_and_U11 ( .A1(cell_2069_a_HPC2_and_a_reg[0]), .A2(
        cell_2069_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2069_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2069_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2069_a_HPC2_and_n9), 
        .ZN(cell_2069_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2069_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2069_a_HPC2_and_n9), 
        .ZN(cell_2069_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2069_a_HPC2_and_U8 ( .A(Fresh[355]), .ZN(cell_2069_a_HPC2_and_n9) );
  AND2_X1 cell_2069_a_HPC2_and_U7 ( .A1(cell_2069_and_in[1]), .A2(n469), .ZN(
        cell_2069_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2069_a_HPC2_and_U6 ( .A1(cell_2069_and_in[0]), .A2(n465), .ZN(
        cell_2069_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2069_a_HPC2_and_U5 ( .A(cell_2069_a_HPC2_and_n8), .B(
        cell_2069_a_HPC2_and_z_1__1_), .ZN(cell_2069_and_out[1]) );
  XNOR2_X1 cell_2069_a_HPC2_and_U4 ( .A(
        cell_2069_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2069_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2069_a_HPC2_and_n8) );
  XNOR2_X1 cell_2069_a_HPC2_and_U3 ( .A(cell_2069_a_HPC2_and_n7), .B(
        cell_2069_a_HPC2_and_z_0__0_), .ZN(cell_2069_and_out[0]) );
  XNOR2_X1 cell_2069_a_HPC2_and_U2 ( .A(
        cell_2069_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2069_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2069_a_HPC2_and_n7) );
  DFF_X1 cell_2069_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2069_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2069_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2069_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2069_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2069_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2069_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2069_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2069_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2069_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2070_U4 ( .A(signal_3746), .B(cell_2070_and_out[1]), .Z(
        signal_3984) );
  XOR2_X1 cell_2070_U3 ( .A(signal_2236), .B(cell_2070_and_out[0]), .Z(
        signal_2338) );
  XOR2_X1 cell_2070_U2 ( .A(signal_3746), .B(signal_3711), .Z(
        cell_2070_and_in[1]) );
  XOR2_X1 cell_2070_U1 ( .A(signal_2236), .B(signal_2201), .Z(
        cell_2070_and_in[0]) );
  XOR2_X1 cell_2070_a_HPC2_and_U14 ( .A(Fresh[356]), .B(cell_2070_and_in[0]), 
        .Z(cell_2070_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2070_a_HPC2_and_U13 ( .A(Fresh[356]), .B(cell_2070_and_in[1]), 
        .Z(cell_2070_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2070_a_HPC2_and_U12 ( .A1(cell_2070_a_HPC2_and_a_reg[1]), .A2(
        cell_2070_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2070_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2070_a_HPC2_and_U11 ( .A1(cell_2070_a_HPC2_and_a_reg[0]), .A2(
        cell_2070_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2070_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2070_a_HPC2_and_U10 ( .A1(n468), .A2(cell_2070_a_HPC2_and_n9), 
        .ZN(cell_2070_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2070_a_HPC2_and_U9 ( .A1(n464), .A2(cell_2070_a_HPC2_and_n9), 
        .ZN(cell_2070_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2070_a_HPC2_and_U8 ( .A(Fresh[356]), .ZN(cell_2070_a_HPC2_and_n9) );
  AND2_X1 cell_2070_a_HPC2_and_U7 ( .A1(cell_2070_and_in[1]), .A2(n468), .ZN(
        cell_2070_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2070_a_HPC2_and_U6 ( .A1(cell_2070_and_in[0]), .A2(n464), .ZN(
        cell_2070_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2070_a_HPC2_and_U5 ( .A(cell_2070_a_HPC2_and_n8), .B(
        cell_2070_a_HPC2_and_z_1__1_), .ZN(cell_2070_and_out[1]) );
  XNOR2_X1 cell_2070_a_HPC2_and_U4 ( .A(
        cell_2070_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2070_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2070_a_HPC2_and_n8) );
  XNOR2_X1 cell_2070_a_HPC2_and_U3 ( .A(cell_2070_a_HPC2_and_n7), .B(
        cell_2070_a_HPC2_and_z_0__0_), .ZN(cell_2070_and_out[0]) );
  XNOR2_X1 cell_2070_a_HPC2_and_U2 ( .A(
        cell_2070_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2070_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2070_a_HPC2_and_n7) );
  DFF_X1 cell_2070_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2070_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2070_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n464), .CK(clk), 
        .Q(cell_2070_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2070_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2070_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n468), .CK(clk), 
        .Q(cell_2070_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2070_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2070_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2070_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2071_U4 ( .A(signal_3740), .B(cell_2071_and_out[1]), .Z(
        signal_3985) );
  XOR2_X1 cell_2071_U3 ( .A(signal_2230), .B(cell_2071_and_out[0]), .Z(
        signal_2339) );
  XOR2_X1 cell_2071_U2 ( .A(signal_3740), .B(signal_3695), .Z(
        cell_2071_and_in[1]) );
  XOR2_X1 cell_2071_U1 ( .A(signal_2230), .B(signal_2185), .Z(
        cell_2071_and_in[0]) );
  XOR2_X1 cell_2071_a_HPC2_and_U14 ( .A(Fresh[357]), .B(cell_2071_and_in[0]), 
        .Z(cell_2071_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2071_a_HPC2_and_U13 ( .A(Fresh[357]), .B(cell_2071_and_in[1]), 
        .Z(cell_2071_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2071_a_HPC2_and_U12 ( .A1(cell_2071_a_HPC2_and_a_reg[1]), .A2(
        cell_2071_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2071_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2071_a_HPC2_and_U11 ( .A1(cell_2071_a_HPC2_and_a_reg[0]), .A2(
        cell_2071_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2071_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2071_a_HPC2_and_U10 ( .A1(n469), .A2(cell_2071_a_HPC2_and_n9), 
        .ZN(cell_2071_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2071_a_HPC2_and_U9 ( .A1(n465), .A2(cell_2071_a_HPC2_and_n9), 
        .ZN(cell_2071_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2071_a_HPC2_and_U8 ( .A(Fresh[357]), .ZN(cell_2071_a_HPC2_and_n9) );
  AND2_X1 cell_2071_a_HPC2_and_U7 ( .A1(cell_2071_and_in[1]), .A2(n469), .ZN(
        cell_2071_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2071_a_HPC2_and_U6 ( .A1(cell_2071_and_in[0]), .A2(n465), .ZN(
        cell_2071_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2071_a_HPC2_and_U5 ( .A(cell_2071_a_HPC2_and_n8), .B(
        cell_2071_a_HPC2_and_z_1__1_), .ZN(cell_2071_and_out[1]) );
  XNOR2_X1 cell_2071_a_HPC2_and_U4 ( .A(
        cell_2071_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2071_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2071_a_HPC2_and_n8) );
  XNOR2_X1 cell_2071_a_HPC2_and_U3 ( .A(cell_2071_a_HPC2_and_n7), .B(
        cell_2071_a_HPC2_and_z_0__0_), .ZN(cell_2071_and_out[0]) );
  XNOR2_X1 cell_2071_a_HPC2_and_U2 ( .A(
        cell_2071_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2071_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2071_a_HPC2_and_n7) );
  DFF_X1 cell_2071_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2071_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2071_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n465), .CK(clk), 
        .Q(cell_2071_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2071_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2071_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n469), .CK(clk), 
        .Q(cell_2071_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2071_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2071_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2071_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2072_U4 ( .A(signal_3944), .B(cell_2072_and_out[1]), .Z(
        signal_4090) );
  XOR2_X1 cell_2072_U3 ( .A(signal_2298), .B(cell_2072_and_out[0]), .Z(
        signal_2340) );
  XOR2_X1 cell_2072_U2 ( .A(signal_3944), .B(signal_3929), .Z(
        cell_2072_and_in[1]) );
  XOR2_X1 cell_2072_U1 ( .A(signal_2298), .B(signal_2283), .Z(
        cell_2072_and_in[0]) );
  XOR2_X1 cell_2072_a_HPC2_and_U14 ( .A(Fresh[358]), .B(cell_2072_and_in[0]), 
        .Z(cell_2072_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2072_a_HPC2_and_U13 ( .A(Fresh[358]), .B(cell_2072_and_in[1]), 
        .Z(cell_2072_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2072_a_HPC2_and_U12 ( .A1(cell_2072_a_HPC2_and_a_reg[1]), .A2(
        cell_2072_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2072_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2072_a_HPC2_and_U11 ( .A1(cell_2072_a_HPC2_and_a_reg[0]), .A2(
        cell_2072_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2072_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2072_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2072_a_HPC2_and_n9), 
        .ZN(cell_2072_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2072_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2072_a_HPC2_and_n9), 
        .ZN(cell_2072_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2072_a_HPC2_and_U8 ( .A(Fresh[358]), .ZN(cell_2072_a_HPC2_and_n9) );
  AND2_X1 cell_2072_a_HPC2_and_U7 ( .A1(cell_2072_and_in[1]), .A2(n459), .ZN(
        cell_2072_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2072_a_HPC2_and_U6 ( .A1(cell_2072_and_in[0]), .A2(n456), .ZN(
        cell_2072_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2072_a_HPC2_and_U5 ( .A(cell_2072_a_HPC2_and_n8), .B(
        cell_2072_a_HPC2_and_z_1__1_), .ZN(cell_2072_and_out[1]) );
  XNOR2_X1 cell_2072_a_HPC2_and_U4 ( .A(
        cell_2072_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2072_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2072_a_HPC2_and_n8) );
  XNOR2_X1 cell_2072_a_HPC2_and_U3 ( .A(cell_2072_a_HPC2_and_n7), .B(
        cell_2072_a_HPC2_and_z_0__0_), .ZN(cell_2072_and_out[0]) );
  XNOR2_X1 cell_2072_a_HPC2_and_U2 ( .A(
        cell_2072_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2072_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2072_a_HPC2_and_n7) );
  DFF_X1 cell_2072_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2072_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2072_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2072_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2072_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2072_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2072_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2072_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2072_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2072_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2073_U4 ( .A(signal_3942), .B(cell_2073_and_out[1]), .Z(
        signal_4091) );
  XOR2_X1 cell_2073_U3 ( .A(signal_2296), .B(cell_2073_and_out[0]), .Z(
        signal_2341) );
  XOR2_X1 cell_2073_U2 ( .A(signal_3942), .B(signal_3968), .Z(
        cell_2073_and_in[1]) );
  XOR2_X1 cell_2073_U1 ( .A(signal_2296), .B(signal_2322), .Z(
        cell_2073_and_in[0]) );
  XOR2_X1 cell_2073_a_HPC2_and_U14 ( .A(Fresh[359]), .B(cell_2073_and_in[0]), 
        .Z(cell_2073_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2073_a_HPC2_and_U13 ( .A(Fresh[359]), .B(cell_2073_and_in[1]), 
        .Z(cell_2073_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2073_a_HPC2_and_U12 ( .A1(cell_2073_a_HPC2_and_a_reg[1]), .A2(
        cell_2073_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2073_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2073_a_HPC2_and_U11 ( .A1(cell_2073_a_HPC2_and_a_reg[0]), .A2(
        cell_2073_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2073_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2073_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2073_a_HPC2_and_n9), 
        .ZN(cell_2073_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2073_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2073_a_HPC2_and_n9), 
        .ZN(cell_2073_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2073_a_HPC2_and_U8 ( .A(Fresh[359]), .ZN(cell_2073_a_HPC2_and_n9) );
  AND2_X1 cell_2073_a_HPC2_and_U7 ( .A1(cell_2073_and_in[1]), .A2(n460), .ZN(
        cell_2073_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2073_a_HPC2_and_U6 ( .A1(cell_2073_and_in[0]), .A2(n457), .ZN(
        cell_2073_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2073_a_HPC2_and_U5 ( .A(cell_2073_a_HPC2_and_n8), .B(
        cell_2073_a_HPC2_and_z_1__1_), .ZN(cell_2073_and_out[1]) );
  XNOR2_X1 cell_2073_a_HPC2_and_U4 ( .A(
        cell_2073_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2073_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2073_a_HPC2_and_n8) );
  XNOR2_X1 cell_2073_a_HPC2_and_U3 ( .A(cell_2073_a_HPC2_and_n7), .B(
        cell_2073_a_HPC2_and_z_0__0_), .ZN(cell_2073_and_out[0]) );
  XNOR2_X1 cell_2073_a_HPC2_and_U2 ( .A(
        cell_2073_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2073_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2073_a_HPC2_and_n7) );
  DFF_X1 cell_2073_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2073_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2073_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2073_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2073_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2073_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2073_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2073_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2073_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2073_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2074_U4 ( .A(signal_3972), .B(cell_2074_and_out[1]), .Z(
        signal_4092) );
  XOR2_X1 cell_2074_U3 ( .A(signal_2326), .B(cell_2074_and_out[0]), .Z(
        signal_2342) );
  XOR2_X1 cell_2074_U2 ( .A(signal_3972), .B(signal_3928), .Z(
        cell_2074_and_in[1]) );
  XOR2_X1 cell_2074_U1 ( .A(signal_2326), .B(signal_2282), .Z(
        cell_2074_and_in[0]) );
  XOR2_X1 cell_2074_a_HPC2_and_U14 ( .A(Fresh[360]), .B(cell_2074_and_in[0]), 
        .Z(cell_2074_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2074_a_HPC2_and_U13 ( .A(Fresh[360]), .B(cell_2074_and_in[1]), 
        .Z(cell_2074_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2074_a_HPC2_and_U12 ( .A1(cell_2074_a_HPC2_and_a_reg[1]), .A2(
        cell_2074_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2074_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2074_a_HPC2_and_U11 ( .A1(cell_2074_a_HPC2_and_a_reg[0]), .A2(
        cell_2074_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2074_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2074_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2074_a_HPC2_and_n9), 
        .ZN(cell_2074_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2074_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2074_a_HPC2_and_n9), 
        .ZN(cell_2074_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2074_a_HPC2_and_U8 ( .A(Fresh[360]), .ZN(cell_2074_a_HPC2_and_n9) );
  AND2_X1 cell_2074_a_HPC2_and_U7 ( .A1(cell_2074_and_in[1]), .A2(n461), .ZN(
        cell_2074_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2074_a_HPC2_and_U6 ( .A1(cell_2074_and_in[0]), .A2(n458), .ZN(
        cell_2074_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2074_a_HPC2_and_U5 ( .A(cell_2074_a_HPC2_and_n8), .B(
        cell_2074_a_HPC2_and_z_1__1_), .ZN(cell_2074_and_out[1]) );
  XNOR2_X1 cell_2074_a_HPC2_and_U4 ( .A(
        cell_2074_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2074_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2074_a_HPC2_and_n8) );
  XNOR2_X1 cell_2074_a_HPC2_and_U3 ( .A(cell_2074_a_HPC2_and_n7), .B(
        cell_2074_a_HPC2_and_z_0__0_), .ZN(cell_2074_and_out[0]) );
  XNOR2_X1 cell_2074_a_HPC2_and_U2 ( .A(
        cell_2074_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2074_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2074_a_HPC2_and_n7) );
  DFF_X1 cell_2074_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2074_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2074_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2074_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2074_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2074_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2074_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2074_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2074_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2074_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2075_U4 ( .A(signal_3980), .B(cell_2075_and_out[1]), .Z(
        signal_4093) );
  XOR2_X1 cell_2075_U3 ( .A(signal_2334), .B(cell_2075_and_out[0]), .Z(
        signal_2343) );
  XOR2_X1 cell_2075_U2 ( .A(signal_3980), .B(signal_3958), .Z(
        cell_2075_and_in[1]) );
  XOR2_X1 cell_2075_U1 ( .A(signal_2334), .B(signal_2312), .Z(
        cell_2075_and_in[0]) );
  XOR2_X1 cell_2075_a_HPC2_and_U14 ( .A(Fresh[361]), .B(cell_2075_and_in[0]), 
        .Z(cell_2075_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2075_a_HPC2_and_U13 ( .A(Fresh[361]), .B(cell_2075_and_in[1]), 
        .Z(cell_2075_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2075_a_HPC2_and_U12 ( .A1(cell_2075_a_HPC2_and_a_reg[1]), .A2(
        cell_2075_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2075_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2075_a_HPC2_and_U11 ( .A1(cell_2075_a_HPC2_and_a_reg[0]), .A2(
        cell_2075_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2075_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2075_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2075_a_HPC2_and_n9), .ZN(cell_2075_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2075_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2075_a_HPC2_and_n9), .ZN(cell_2075_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2075_a_HPC2_and_U8 ( .A(Fresh[361]), .ZN(cell_2075_a_HPC2_and_n9) );
  AND2_X1 cell_2075_a_HPC2_and_U7 ( .A1(cell_2075_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2075_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2075_a_HPC2_and_U6 ( .A1(cell_2075_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2075_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2075_a_HPC2_and_U5 ( .A(cell_2075_a_HPC2_and_n8), .B(
        cell_2075_a_HPC2_and_z_1__1_), .ZN(cell_2075_and_out[1]) );
  XNOR2_X1 cell_2075_a_HPC2_and_U4 ( .A(
        cell_2075_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2075_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2075_a_HPC2_and_n8) );
  XNOR2_X1 cell_2075_a_HPC2_and_U3 ( .A(cell_2075_a_HPC2_and_n7), .B(
        cell_2075_a_HPC2_and_z_0__0_), .ZN(cell_2075_and_out[0]) );
  XNOR2_X1 cell_2075_a_HPC2_and_U2 ( .A(
        cell_2075_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2075_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2075_a_HPC2_and_n7) );
  DFF_X1 cell_2075_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2075_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2075_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2075_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2075_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2075_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2075_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2075_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2075_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2075_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2076_U4 ( .A(signal_3978), .B(cell_2076_and_out[1]), .Z(
        signal_4094) );
  XOR2_X1 cell_2076_U3 ( .A(signal_2332), .B(cell_2076_and_out[0]), .Z(
        signal_2344) );
  XOR2_X1 cell_2076_U2 ( .A(signal_3978), .B(signal_3931), .Z(
        cell_2076_and_in[1]) );
  XOR2_X1 cell_2076_U1 ( .A(signal_2332), .B(signal_2285), .Z(
        cell_2076_and_in[0]) );
  XOR2_X1 cell_2076_a_HPC2_and_U14 ( .A(Fresh[362]), .B(cell_2076_and_in[0]), 
        .Z(cell_2076_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2076_a_HPC2_and_U13 ( .A(Fresh[362]), .B(cell_2076_and_in[1]), 
        .Z(cell_2076_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2076_a_HPC2_and_U12 ( .A1(cell_2076_a_HPC2_and_a_reg[1]), .A2(
        cell_2076_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2076_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2076_a_HPC2_and_U11 ( .A1(cell_2076_a_HPC2_and_a_reg[0]), .A2(
        cell_2076_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2076_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2076_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2076_a_HPC2_and_n9), .ZN(cell_2076_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2076_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2076_a_HPC2_and_n9), .ZN(cell_2076_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2076_a_HPC2_and_U8 ( .A(Fresh[362]), .ZN(cell_2076_a_HPC2_and_n9) );
  AND2_X1 cell_2076_a_HPC2_and_U7 ( .A1(cell_2076_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2076_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2076_a_HPC2_and_U6 ( .A1(cell_2076_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2076_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2076_a_HPC2_and_U5 ( .A(cell_2076_a_HPC2_and_n8), .B(
        cell_2076_a_HPC2_and_z_1__1_), .ZN(cell_2076_and_out[1]) );
  XNOR2_X1 cell_2076_a_HPC2_and_U4 ( .A(
        cell_2076_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2076_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2076_a_HPC2_and_n8) );
  XNOR2_X1 cell_2076_a_HPC2_and_U3 ( .A(cell_2076_a_HPC2_and_n7), .B(
        cell_2076_a_HPC2_and_z_0__0_), .ZN(cell_2076_and_out[0]) );
  XNOR2_X1 cell_2076_a_HPC2_and_U2 ( .A(
        cell_2076_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2076_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2076_a_HPC2_and_n7) );
  DFF_X1 cell_2076_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2076_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2076_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2076_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2076_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2076_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2076_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2076_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2076_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2076_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2077_U4 ( .A(signal_3985), .B(cell_2077_and_out[1]), .Z(
        signal_4095) );
  XOR2_X1 cell_2077_U3 ( .A(signal_2339), .B(cell_2077_and_out[0]), .Z(
        signal_2345) );
  XOR2_X1 cell_2077_U2 ( .A(signal_3985), .B(signal_3979), .Z(
        cell_2077_and_in[1]) );
  XOR2_X1 cell_2077_U1 ( .A(signal_2339), .B(signal_2333), .Z(
        cell_2077_and_in[0]) );
  XOR2_X1 cell_2077_a_HPC2_and_U14 ( .A(Fresh[363]), .B(cell_2077_and_in[0]), 
        .Z(cell_2077_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2077_a_HPC2_and_U13 ( .A(Fresh[363]), .B(cell_2077_and_in[1]), 
        .Z(cell_2077_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2077_a_HPC2_and_U12 ( .A1(cell_2077_a_HPC2_and_a_reg[1]), .A2(
        cell_2077_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2077_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2077_a_HPC2_and_U11 ( .A1(cell_2077_a_HPC2_and_a_reg[0]), .A2(
        cell_2077_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2077_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2077_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2077_a_HPC2_and_n9), .ZN(cell_2077_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2077_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2077_a_HPC2_and_n9), .ZN(cell_2077_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2077_a_HPC2_and_U8 ( .A(Fresh[363]), .ZN(cell_2077_a_HPC2_and_n9) );
  AND2_X1 cell_2077_a_HPC2_and_U7 ( .A1(cell_2077_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2077_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2077_a_HPC2_and_U6 ( .A1(cell_2077_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2077_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2077_a_HPC2_and_U5 ( .A(cell_2077_a_HPC2_and_n8), .B(
        cell_2077_a_HPC2_and_z_1__1_), .ZN(cell_2077_and_out[1]) );
  XNOR2_X1 cell_2077_a_HPC2_and_U4 ( .A(
        cell_2077_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2077_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2077_a_HPC2_and_n8) );
  XNOR2_X1 cell_2077_a_HPC2_and_U3 ( .A(cell_2077_a_HPC2_and_n7), .B(
        cell_2077_a_HPC2_and_z_0__0_), .ZN(cell_2077_and_out[0]) );
  XNOR2_X1 cell_2077_a_HPC2_and_U2 ( .A(
        cell_2077_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2077_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2077_a_HPC2_and_n7) );
  DFF_X1 cell_2077_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2077_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2077_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2077_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2077_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2077_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2077_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2077_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2077_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2077_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2078_U4 ( .A(signal_3966), .B(cell_2078_and_out[1]), .Z(
        signal_4096) );
  XOR2_X1 cell_2078_U3 ( .A(signal_2320), .B(cell_2078_and_out[0]), .Z(
        signal_2346) );
  XOR2_X1 cell_2078_U2 ( .A(signal_3966), .B(signal_3933), .Z(
        cell_2078_and_in[1]) );
  XOR2_X1 cell_2078_U1 ( .A(signal_2320), .B(signal_2287), .Z(
        cell_2078_and_in[0]) );
  XOR2_X1 cell_2078_a_HPC2_and_U14 ( .A(Fresh[364]), .B(cell_2078_and_in[0]), 
        .Z(cell_2078_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2078_a_HPC2_and_U13 ( .A(Fresh[364]), .B(cell_2078_and_in[1]), 
        .Z(cell_2078_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2078_a_HPC2_and_U12 ( .A1(cell_2078_a_HPC2_and_a_reg[1]), .A2(
        cell_2078_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2078_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2078_a_HPC2_and_U11 ( .A1(cell_2078_a_HPC2_and_a_reg[0]), .A2(
        cell_2078_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2078_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2078_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2078_a_HPC2_and_n9), .ZN(cell_2078_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2078_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2078_a_HPC2_and_n9), .ZN(cell_2078_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2078_a_HPC2_and_U8 ( .A(Fresh[364]), .ZN(cell_2078_a_HPC2_and_n9) );
  AND2_X1 cell_2078_a_HPC2_and_U7 ( .A1(cell_2078_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2078_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2078_a_HPC2_and_U6 ( .A1(cell_2078_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2078_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2078_a_HPC2_and_U5 ( .A(cell_2078_a_HPC2_and_n8), .B(
        cell_2078_a_HPC2_and_z_1__1_), .ZN(cell_2078_and_out[1]) );
  XNOR2_X1 cell_2078_a_HPC2_and_U4 ( .A(
        cell_2078_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2078_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2078_a_HPC2_and_n8) );
  XNOR2_X1 cell_2078_a_HPC2_and_U3 ( .A(cell_2078_a_HPC2_and_n7), .B(
        cell_2078_a_HPC2_and_z_0__0_), .ZN(cell_2078_and_out[0]) );
  XNOR2_X1 cell_2078_a_HPC2_and_U2 ( .A(
        cell_2078_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2078_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2078_a_HPC2_and_n7) );
  DFF_X1 cell_2078_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2078_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2078_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2078_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2078_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2078_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2078_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2078_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2078_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2078_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2079_U4 ( .A(signal_3951), .B(cell_2079_and_out[1]), .Z(
        signal_4097) );
  XOR2_X1 cell_2079_U3 ( .A(signal_2305), .B(cell_2079_and_out[0]), .Z(
        signal_2347) );
  XOR2_X1 cell_2079_U2 ( .A(signal_3951), .B(signal_3964), .Z(
        cell_2079_and_in[1]) );
  XOR2_X1 cell_2079_U1 ( .A(signal_2305), .B(signal_2318), .Z(
        cell_2079_and_in[0]) );
  XOR2_X1 cell_2079_a_HPC2_and_U14 ( .A(Fresh[365]), .B(cell_2079_and_in[0]), 
        .Z(cell_2079_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2079_a_HPC2_and_U13 ( .A(Fresh[365]), .B(cell_2079_and_in[1]), 
        .Z(cell_2079_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2079_a_HPC2_and_U12 ( .A1(cell_2079_a_HPC2_and_a_reg[1]), .A2(
        cell_2079_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2079_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2079_a_HPC2_and_U11 ( .A1(cell_2079_a_HPC2_and_a_reg[0]), .A2(
        cell_2079_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2079_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2079_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2079_a_HPC2_and_n9), 
        .ZN(cell_2079_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2079_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2079_a_HPC2_and_n9), 
        .ZN(cell_2079_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2079_a_HPC2_and_U8 ( .A(Fresh[365]), .ZN(cell_2079_a_HPC2_and_n9) );
  AND2_X1 cell_2079_a_HPC2_and_U7 ( .A1(cell_2079_and_in[1]), .A2(n459), .ZN(
        cell_2079_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2079_a_HPC2_and_U6 ( .A1(cell_2079_and_in[0]), .A2(n456), .ZN(
        cell_2079_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2079_a_HPC2_and_U5 ( .A(cell_2079_a_HPC2_and_n8), .B(
        cell_2079_a_HPC2_and_z_1__1_), .ZN(cell_2079_and_out[1]) );
  XNOR2_X1 cell_2079_a_HPC2_and_U4 ( .A(
        cell_2079_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2079_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2079_a_HPC2_and_n8) );
  XNOR2_X1 cell_2079_a_HPC2_and_U3 ( .A(cell_2079_a_HPC2_and_n7), .B(
        cell_2079_a_HPC2_and_z_0__0_), .ZN(cell_2079_and_out[0]) );
  XNOR2_X1 cell_2079_a_HPC2_and_U2 ( .A(
        cell_2079_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2079_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2079_a_HPC2_and_n7) );
  DFF_X1 cell_2079_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2079_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2079_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2079_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2079_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2079_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2079_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2079_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2079_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2079_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2080_U4 ( .A(signal_3924), .B(cell_2080_and_out[1]), .Z(
        signal_4098) );
  XOR2_X1 cell_2080_U3 ( .A(signal_2278), .B(cell_2080_and_out[0]), .Z(
        signal_2348) );
  XOR2_X1 cell_2080_U2 ( .A(signal_3924), .B(signal_3930), .Z(
        cell_2080_and_in[1]) );
  XOR2_X1 cell_2080_U1 ( .A(signal_2278), .B(signal_2284), .Z(
        cell_2080_and_in[0]) );
  XOR2_X1 cell_2080_a_HPC2_and_U14 ( .A(Fresh[366]), .B(cell_2080_and_in[0]), 
        .Z(cell_2080_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2080_a_HPC2_and_U13 ( .A(Fresh[366]), .B(cell_2080_and_in[1]), 
        .Z(cell_2080_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2080_a_HPC2_and_U12 ( .A1(cell_2080_a_HPC2_and_a_reg[1]), .A2(
        cell_2080_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2080_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2080_a_HPC2_and_U11 ( .A1(cell_2080_a_HPC2_and_a_reg[0]), .A2(
        cell_2080_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2080_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2080_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2080_a_HPC2_and_n9), 
        .ZN(cell_2080_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2080_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2080_a_HPC2_and_n9), 
        .ZN(cell_2080_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2080_a_HPC2_and_U8 ( .A(Fresh[366]), .ZN(cell_2080_a_HPC2_and_n9) );
  AND2_X1 cell_2080_a_HPC2_and_U7 ( .A1(cell_2080_and_in[1]), .A2(n459), .ZN(
        cell_2080_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2080_a_HPC2_and_U6 ( .A1(cell_2080_and_in[0]), .A2(n456), .ZN(
        cell_2080_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2080_a_HPC2_and_U5 ( .A(cell_2080_a_HPC2_and_n8), .B(
        cell_2080_a_HPC2_and_z_1__1_), .ZN(cell_2080_and_out[1]) );
  XNOR2_X1 cell_2080_a_HPC2_and_U4 ( .A(
        cell_2080_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2080_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2080_a_HPC2_and_n8) );
  XNOR2_X1 cell_2080_a_HPC2_and_U3 ( .A(cell_2080_a_HPC2_and_n7), .B(
        cell_2080_a_HPC2_and_z_0__0_), .ZN(cell_2080_and_out[0]) );
  XNOR2_X1 cell_2080_a_HPC2_and_U2 ( .A(
        cell_2080_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2080_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2080_a_HPC2_and_n7) );
  DFF_X1 cell_2080_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2080_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2080_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2080_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2080_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2080_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2080_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2080_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2080_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2080_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2081_U4 ( .A(signal_3922), .B(cell_2081_and_out[1]), .Z(
        signal_4099) );
  XOR2_X1 cell_2081_U3 ( .A(signal_2276), .B(cell_2081_and_out[0]), .Z(
        signal_2349) );
  XOR2_X1 cell_2081_U2 ( .A(signal_3922), .B(signal_3975), .Z(
        cell_2081_and_in[1]) );
  XOR2_X1 cell_2081_U1 ( .A(signal_2276), .B(signal_2329), .Z(
        cell_2081_and_in[0]) );
  XOR2_X1 cell_2081_a_HPC2_and_U14 ( .A(Fresh[367]), .B(cell_2081_and_in[0]), 
        .Z(cell_2081_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2081_a_HPC2_and_U13 ( .A(Fresh[367]), .B(cell_2081_and_in[1]), 
        .Z(cell_2081_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2081_a_HPC2_and_U12 ( .A1(cell_2081_a_HPC2_and_a_reg[1]), .A2(
        cell_2081_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2081_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2081_a_HPC2_and_U11 ( .A1(cell_2081_a_HPC2_and_a_reg[0]), .A2(
        cell_2081_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2081_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2081_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2081_a_HPC2_and_n9), 
        .ZN(cell_2081_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2081_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2081_a_HPC2_and_n9), 
        .ZN(cell_2081_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2081_a_HPC2_and_U8 ( .A(Fresh[367]), .ZN(cell_2081_a_HPC2_and_n9) );
  AND2_X1 cell_2081_a_HPC2_and_U7 ( .A1(cell_2081_and_in[1]), .A2(n459), .ZN(
        cell_2081_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2081_a_HPC2_and_U6 ( .A1(cell_2081_and_in[0]), .A2(n456), .ZN(
        cell_2081_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2081_a_HPC2_and_U5 ( .A(cell_2081_a_HPC2_and_n8), .B(
        cell_2081_a_HPC2_and_z_1__1_), .ZN(cell_2081_and_out[1]) );
  XNOR2_X1 cell_2081_a_HPC2_and_U4 ( .A(
        cell_2081_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2081_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2081_a_HPC2_and_n8) );
  XNOR2_X1 cell_2081_a_HPC2_and_U3 ( .A(cell_2081_a_HPC2_and_n7), .B(
        cell_2081_a_HPC2_and_z_0__0_), .ZN(cell_2081_and_out[0]) );
  XNOR2_X1 cell_2081_a_HPC2_and_U2 ( .A(
        cell_2081_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2081_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2081_a_HPC2_and_n7) );
  DFF_X1 cell_2081_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2081_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2081_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2081_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2081_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2081_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2081_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2081_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2081_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2081_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2082_U4 ( .A(signal_3927), .B(cell_2082_and_out[1]), .Z(
        signal_4100) );
  XOR2_X1 cell_2082_U3 ( .A(signal_2281), .B(cell_2082_and_out[0]), .Z(
        signal_2350) );
  XOR2_X1 cell_2082_U2 ( .A(signal_3927), .B(signal_3971), .Z(
        cell_2082_and_in[1]) );
  XOR2_X1 cell_2082_U1 ( .A(signal_2281), .B(signal_2325), .Z(
        cell_2082_and_in[0]) );
  XOR2_X1 cell_2082_a_HPC2_and_U14 ( .A(Fresh[368]), .B(cell_2082_and_in[0]), 
        .Z(cell_2082_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2082_a_HPC2_and_U13 ( .A(Fresh[368]), .B(cell_2082_and_in[1]), 
        .Z(cell_2082_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2082_a_HPC2_and_U12 ( .A1(cell_2082_a_HPC2_and_a_reg[1]), .A2(
        cell_2082_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2082_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2082_a_HPC2_and_U11 ( .A1(cell_2082_a_HPC2_and_a_reg[0]), .A2(
        cell_2082_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2082_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2082_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2082_a_HPC2_and_n9), 
        .ZN(cell_2082_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2082_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2082_a_HPC2_and_n9), 
        .ZN(cell_2082_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2082_a_HPC2_and_U8 ( .A(Fresh[368]), .ZN(cell_2082_a_HPC2_and_n9) );
  AND2_X1 cell_2082_a_HPC2_and_U7 ( .A1(cell_2082_and_in[1]), .A2(n459), .ZN(
        cell_2082_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2082_a_HPC2_and_U6 ( .A1(cell_2082_and_in[0]), .A2(n456), .ZN(
        cell_2082_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2082_a_HPC2_and_U5 ( .A(cell_2082_a_HPC2_and_n8), .B(
        cell_2082_a_HPC2_and_z_1__1_), .ZN(cell_2082_and_out[1]) );
  XNOR2_X1 cell_2082_a_HPC2_and_U4 ( .A(
        cell_2082_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2082_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2082_a_HPC2_and_n8) );
  XNOR2_X1 cell_2082_a_HPC2_and_U3 ( .A(cell_2082_a_HPC2_and_n7), .B(
        cell_2082_a_HPC2_and_z_0__0_), .ZN(cell_2082_and_out[0]) );
  XNOR2_X1 cell_2082_a_HPC2_and_U2 ( .A(
        cell_2082_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2082_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2082_a_HPC2_and_n7) );
  DFF_X1 cell_2082_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2082_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2082_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2082_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2082_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2082_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2082_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2082_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2082_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2082_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2083_U4 ( .A(signal_3938), .B(cell_2083_and_out[1]), .Z(
        signal_4101) );
  XOR2_X1 cell_2083_U3 ( .A(signal_2292), .B(cell_2083_and_out[0]), .Z(
        signal_2351) );
  XOR2_X1 cell_2083_U2 ( .A(signal_3938), .B(signal_3926), .Z(
        cell_2083_and_in[1]) );
  XOR2_X1 cell_2083_U1 ( .A(signal_2292), .B(signal_2280), .Z(
        cell_2083_and_in[0]) );
  XOR2_X1 cell_2083_a_HPC2_and_U14 ( .A(Fresh[369]), .B(cell_2083_and_in[0]), 
        .Z(cell_2083_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2083_a_HPC2_and_U13 ( .A(Fresh[369]), .B(cell_2083_and_in[1]), 
        .Z(cell_2083_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2083_a_HPC2_and_U12 ( .A1(cell_2083_a_HPC2_and_a_reg[1]), .A2(
        cell_2083_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2083_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2083_a_HPC2_and_U11 ( .A1(cell_2083_a_HPC2_and_a_reg[0]), .A2(
        cell_2083_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2083_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2083_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2083_a_HPC2_and_n9), 
        .ZN(cell_2083_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2083_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2083_a_HPC2_and_n9), 
        .ZN(cell_2083_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2083_a_HPC2_and_U8 ( .A(Fresh[369]), .ZN(cell_2083_a_HPC2_and_n9) );
  AND2_X1 cell_2083_a_HPC2_and_U7 ( .A1(cell_2083_and_in[1]), .A2(n459), .ZN(
        cell_2083_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2083_a_HPC2_and_U6 ( .A1(cell_2083_and_in[0]), .A2(n456), .ZN(
        cell_2083_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2083_a_HPC2_and_U5 ( .A(cell_2083_a_HPC2_and_n8), .B(
        cell_2083_a_HPC2_and_z_1__1_), .ZN(cell_2083_and_out[1]) );
  XNOR2_X1 cell_2083_a_HPC2_and_U4 ( .A(
        cell_2083_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2083_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2083_a_HPC2_and_n8) );
  XNOR2_X1 cell_2083_a_HPC2_and_U3 ( .A(cell_2083_a_HPC2_and_n7), .B(
        cell_2083_a_HPC2_and_z_0__0_), .ZN(cell_2083_and_out[0]) );
  XNOR2_X1 cell_2083_a_HPC2_and_U2 ( .A(
        cell_2083_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2083_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2083_a_HPC2_and_n7) );
  DFF_X1 cell_2083_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2083_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2083_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2083_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2083_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2083_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2083_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2083_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2083_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2083_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2084_U4 ( .A(signal_3936), .B(cell_2084_and_out[1]), .Z(
        signal_4102) );
  XOR2_X1 cell_2084_U3 ( .A(signal_2290), .B(cell_2084_and_out[0]), .Z(
        signal_2352) );
  XOR2_X1 cell_2084_U2 ( .A(signal_3936), .B(signal_3970), .Z(
        cell_2084_and_in[1]) );
  XOR2_X1 cell_2084_U1 ( .A(signal_2290), .B(signal_2324), .Z(
        cell_2084_and_in[0]) );
  XOR2_X1 cell_2084_a_HPC2_and_U14 ( .A(Fresh[370]), .B(cell_2084_and_in[0]), 
        .Z(cell_2084_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2084_a_HPC2_and_U13 ( .A(Fresh[370]), .B(cell_2084_and_in[1]), 
        .Z(cell_2084_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2084_a_HPC2_and_U12 ( .A1(cell_2084_a_HPC2_and_a_reg[1]), .A2(
        cell_2084_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2084_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2084_a_HPC2_and_U11 ( .A1(cell_2084_a_HPC2_and_a_reg[0]), .A2(
        cell_2084_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2084_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2084_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2084_a_HPC2_and_n9), 
        .ZN(cell_2084_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2084_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2084_a_HPC2_and_n9), 
        .ZN(cell_2084_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2084_a_HPC2_and_U8 ( .A(Fresh[370]), .ZN(cell_2084_a_HPC2_and_n9) );
  AND2_X1 cell_2084_a_HPC2_and_U7 ( .A1(cell_2084_and_in[1]), .A2(n459), .ZN(
        cell_2084_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2084_a_HPC2_and_U6 ( .A1(cell_2084_and_in[0]), .A2(n456), .ZN(
        cell_2084_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2084_a_HPC2_and_U5 ( .A(cell_2084_a_HPC2_and_n8), .B(
        cell_2084_a_HPC2_and_z_1__1_), .ZN(cell_2084_and_out[1]) );
  XNOR2_X1 cell_2084_a_HPC2_and_U4 ( .A(
        cell_2084_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2084_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2084_a_HPC2_and_n8) );
  XNOR2_X1 cell_2084_a_HPC2_and_U3 ( .A(cell_2084_a_HPC2_and_n7), .B(
        cell_2084_a_HPC2_and_z_0__0_), .ZN(cell_2084_and_out[0]) );
  XNOR2_X1 cell_2084_a_HPC2_and_U2 ( .A(
        cell_2084_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2084_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2084_a_HPC2_and_n7) );
  DFF_X1 cell_2084_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2084_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2084_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2084_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2084_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2084_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2084_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2084_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2084_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2084_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2085_U4 ( .A(signal_3939), .B(cell_2085_and_out[1]), .Z(
        signal_4103) );
  XOR2_X1 cell_2085_U3 ( .A(signal_2293), .B(cell_2085_and_out[0]), .Z(
        signal_2353) );
  XOR2_X1 cell_2085_U2 ( .A(signal_3939), .B(signal_3956), .Z(
        cell_2085_and_in[1]) );
  XOR2_X1 cell_2085_U1 ( .A(signal_2293), .B(signal_2310), .Z(
        cell_2085_and_in[0]) );
  XOR2_X1 cell_2085_a_HPC2_and_U14 ( .A(Fresh[371]), .B(cell_2085_and_in[0]), 
        .Z(cell_2085_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2085_a_HPC2_and_U13 ( .A(Fresh[371]), .B(cell_2085_and_in[1]), 
        .Z(cell_2085_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2085_a_HPC2_and_U12 ( .A1(cell_2085_a_HPC2_and_a_reg[1]), .A2(
        cell_2085_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2085_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2085_a_HPC2_and_U11 ( .A1(cell_2085_a_HPC2_and_a_reg[0]), .A2(
        cell_2085_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2085_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2085_a_HPC2_and_U10 ( .A1(n459), .A2(cell_2085_a_HPC2_and_n9), 
        .ZN(cell_2085_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2085_a_HPC2_and_U9 ( .A1(n456), .A2(cell_2085_a_HPC2_and_n9), 
        .ZN(cell_2085_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2085_a_HPC2_and_U8 ( .A(Fresh[371]), .ZN(cell_2085_a_HPC2_and_n9) );
  AND2_X1 cell_2085_a_HPC2_and_U7 ( .A1(cell_2085_and_in[1]), .A2(n459), .ZN(
        cell_2085_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2085_a_HPC2_and_U6 ( .A1(cell_2085_and_in[0]), .A2(n456), .ZN(
        cell_2085_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2085_a_HPC2_and_U5 ( .A(cell_2085_a_HPC2_and_n8), .B(
        cell_2085_a_HPC2_and_z_1__1_), .ZN(cell_2085_and_out[1]) );
  XNOR2_X1 cell_2085_a_HPC2_and_U4 ( .A(
        cell_2085_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2085_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2085_a_HPC2_and_n8) );
  XNOR2_X1 cell_2085_a_HPC2_and_U3 ( .A(cell_2085_a_HPC2_and_n7), .B(
        cell_2085_a_HPC2_and_z_0__0_), .ZN(cell_2085_and_out[0]) );
  XNOR2_X1 cell_2085_a_HPC2_and_U2 ( .A(
        cell_2085_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2085_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2085_a_HPC2_and_n7) );
  DFF_X1 cell_2085_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2085_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2085_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n456), .CK(clk), 
        .Q(cell_2085_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2085_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2085_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n459), .CK(clk), 
        .Q(cell_2085_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2085_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2085_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2085_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2086_U4 ( .A(signal_3947), .B(cell_2086_and_out[1]), .Z(
        signal_4104) );
  XOR2_X1 cell_2086_U3 ( .A(signal_2301), .B(cell_2086_and_out[0]), .Z(
        signal_2354) );
  XOR2_X1 cell_2086_U2 ( .A(signal_3947), .B(signal_3961), .Z(
        cell_2086_and_in[1]) );
  XOR2_X1 cell_2086_U1 ( .A(signal_2301), .B(signal_2315), .Z(
        cell_2086_and_in[0]) );
  XOR2_X1 cell_2086_a_HPC2_and_U14 ( .A(Fresh[372]), .B(cell_2086_and_in[0]), 
        .Z(cell_2086_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2086_a_HPC2_and_U13 ( .A(Fresh[372]), .B(cell_2086_and_in[1]), 
        .Z(cell_2086_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2086_a_HPC2_and_U12 ( .A1(cell_2086_a_HPC2_and_a_reg[1]), .A2(
        cell_2086_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2086_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2086_a_HPC2_and_U11 ( .A1(cell_2086_a_HPC2_and_a_reg[0]), .A2(
        cell_2086_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2086_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2086_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2086_a_HPC2_and_n9), 
        .ZN(cell_2086_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2086_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2086_a_HPC2_and_n9), 
        .ZN(cell_2086_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2086_a_HPC2_and_U8 ( .A(Fresh[372]), .ZN(cell_2086_a_HPC2_and_n9) );
  AND2_X1 cell_2086_a_HPC2_and_U7 ( .A1(cell_2086_and_in[1]), .A2(n460), .ZN(
        cell_2086_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2086_a_HPC2_and_U6 ( .A1(cell_2086_and_in[0]), .A2(n457), .ZN(
        cell_2086_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2086_a_HPC2_and_U5 ( .A(cell_2086_a_HPC2_and_n8), .B(
        cell_2086_a_HPC2_and_z_1__1_), .ZN(cell_2086_and_out[1]) );
  XNOR2_X1 cell_2086_a_HPC2_and_U4 ( .A(
        cell_2086_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2086_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2086_a_HPC2_and_n8) );
  XNOR2_X1 cell_2086_a_HPC2_and_U3 ( .A(cell_2086_a_HPC2_and_n7), .B(
        cell_2086_a_HPC2_and_z_0__0_), .ZN(cell_2086_and_out[0]) );
  XNOR2_X1 cell_2086_a_HPC2_and_U2 ( .A(
        cell_2086_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2086_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2086_a_HPC2_and_n7) );
  DFF_X1 cell_2086_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2086_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2086_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2086_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2086_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2086_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2086_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2086_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2086_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2086_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2087_U4 ( .A(signal_3981), .B(cell_2087_and_out[1]), .Z(
        signal_4105) );
  XOR2_X1 cell_2087_U3 ( .A(signal_2335), .B(cell_2087_and_out[0]), .Z(
        signal_2355) );
  XOR2_X1 cell_2087_U2 ( .A(signal_3981), .B(signal_3983), .Z(
        cell_2087_and_in[1]) );
  XOR2_X1 cell_2087_U1 ( .A(signal_2335), .B(signal_2337), .Z(
        cell_2087_and_in[0]) );
  XOR2_X1 cell_2087_a_HPC2_and_U14 ( .A(Fresh[373]), .B(cell_2087_and_in[0]), 
        .Z(cell_2087_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2087_a_HPC2_and_U13 ( .A(Fresh[373]), .B(cell_2087_and_in[1]), 
        .Z(cell_2087_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2087_a_HPC2_and_U12 ( .A1(cell_2087_a_HPC2_and_a_reg[1]), .A2(
        cell_2087_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2087_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2087_a_HPC2_and_U11 ( .A1(cell_2087_a_HPC2_and_a_reg[0]), .A2(
        cell_2087_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2087_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2087_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2087_a_HPC2_and_n9), 
        .ZN(cell_2087_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2087_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2087_a_HPC2_and_n9), 
        .ZN(cell_2087_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2087_a_HPC2_and_U8 ( .A(Fresh[373]), .ZN(cell_2087_a_HPC2_and_n9) );
  AND2_X1 cell_2087_a_HPC2_and_U7 ( .A1(cell_2087_and_in[1]), .A2(n460), .ZN(
        cell_2087_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2087_a_HPC2_and_U6 ( .A1(cell_2087_and_in[0]), .A2(n457), .ZN(
        cell_2087_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2087_a_HPC2_and_U5 ( .A(cell_2087_a_HPC2_and_n8), .B(
        cell_2087_a_HPC2_and_z_1__1_), .ZN(cell_2087_and_out[1]) );
  XNOR2_X1 cell_2087_a_HPC2_and_U4 ( .A(
        cell_2087_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2087_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2087_a_HPC2_and_n8) );
  XNOR2_X1 cell_2087_a_HPC2_and_U3 ( .A(cell_2087_a_HPC2_and_n7), .B(
        cell_2087_a_HPC2_and_z_0__0_), .ZN(cell_2087_and_out[0]) );
  XNOR2_X1 cell_2087_a_HPC2_and_U2 ( .A(
        cell_2087_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2087_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2087_a_HPC2_and_n7) );
  DFF_X1 cell_2087_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2087_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2087_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2087_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2087_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2087_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2087_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2087_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2087_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2087_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2088_U4 ( .A(signal_3949), .B(cell_2088_and_out[1]), .Z(
        signal_4106) );
  XOR2_X1 cell_2088_U3 ( .A(signal_2303), .B(cell_2088_and_out[0]), .Z(
        signal_2356) );
  XOR2_X1 cell_2088_U2 ( .A(signal_3949), .B(signal_3974), .Z(
        cell_2088_and_in[1]) );
  XOR2_X1 cell_2088_U1 ( .A(signal_2303), .B(signal_2328), .Z(
        cell_2088_and_in[0]) );
  XOR2_X1 cell_2088_a_HPC2_and_U14 ( .A(Fresh[374]), .B(cell_2088_and_in[0]), 
        .Z(cell_2088_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2088_a_HPC2_and_U13 ( .A(Fresh[374]), .B(cell_2088_and_in[1]), 
        .Z(cell_2088_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2088_a_HPC2_and_U12 ( .A1(cell_2088_a_HPC2_and_a_reg[1]), .A2(
        cell_2088_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2088_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2088_a_HPC2_and_U11 ( .A1(cell_2088_a_HPC2_and_a_reg[0]), .A2(
        cell_2088_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2088_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2088_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2088_a_HPC2_and_n9), 
        .ZN(cell_2088_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2088_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2088_a_HPC2_and_n9), 
        .ZN(cell_2088_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2088_a_HPC2_and_U8 ( .A(Fresh[374]), .ZN(cell_2088_a_HPC2_and_n9) );
  AND2_X1 cell_2088_a_HPC2_and_U7 ( .A1(cell_2088_and_in[1]), .A2(n460), .ZN(
        cell_2088_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2088_a_HPC2_and_U6 ( .A1(cell_2088_and_in[0]), .A2(n457), .ZN(
        cell_2088_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2088_a_HPC2_and_U5 ( .A(cell_2088_a_HPC2_and_n8), .B(
        cell_2088_a_HPC2_and_z_1__1_), .ZN(cell_2088_and_out[1]) );
  XNOR2_X1 cell_2088_a_HPC2_and_U4 ( .A(
        cell_2088_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2088_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2088_a_HPC2_and_n8) );
  XNOR2_X1 cell_2088_a_HPC2_and_U3 ( .A(cell_2088_a_HPC2_and_n7), .B(
        cell_2088_a_HPC2_and_z_0__0_), .ZN(cell_2088_and_out[0]) );
  XNOR2_X1 cell_2088_a_HPC2_and_U2 ( .A(
        cell_2088_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2088_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2088_a_HPC2_and_n7) );
  DFF_X1 cell_2088_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2088_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2088_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2088_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2088_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2088_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2088_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2088_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2088_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2088_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2089_U4 ( .A(signal_3960), .B(cell_2089_and_out[1]), .Z(
        signal_4107) );
  XOR2_X1 cell_2089_U3 ( .A(signal_2314), .B(cell_2089_and_out[0]), .Z(
        signal_2357) );
  XOR2_X1 cell_2089_U2 ( .A(signal_3960), .B(signal_3937), .Z(
        cell_2089_and_in[1]) );
  XOR2_X1 cell_2089_U1 ( .A(signal_2314), .B(signal_2291), .Z(
        cell_2089_and_in[0]) );
  XOR2_X1 cell_2089_a_HPC2_and_U14 ( .A(Fresh[375]), .B(cell_2089_and_in[0]), 
        .Z(cell_2089_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2089_a_HPC2_and_U13 ( .A(Fresh[375]), .B(cell_2089_and_in[1]), 
        .Z(cell_2089_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2089_a_HPC2_and_U12 ( .A1(cell_2089_a_HPC2_and_a_reg[1]), .A2(
        cell_2089_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2089_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2089_a_HPC2_and_U11 ( .A1(cell_2089_a_HPC2_and_a_reg[0]), .A2(
        cell_2089_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2089_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2089_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2089_a_HPC2_and_n9), 
        .ZN(cell_2089_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2089_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2089_a_HPC2_and_n9), 
        .ZN(cell_2089_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2089_a_HPC2_and_U8 ( .A(Fresh[375]), .ZN(cell_2089_a_HPC2_and_n9) );
  AND2_X1 cell_2089_a_HPC2_and_U7 ( .A1(cell_2089_and_in[1]), .A2(n460), .ZN(
        cell_2089_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2089_a_HPC2_and_U6 ( .A1(cell_2089_and_in[0]), .A2(n457), .ZN(
        cell_2089_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2089_a_HPC2_and_U5 ( .A(cell_2089_a_HPC2_and_n8), .B(
        cell_2089_a_HPC2_and_z_1__1_), .ZN(cell_2089_and_out[1]) );
  XNOR2_X1 cell_2089_a_HPC2_and_U4 ( .A(
        cell_2089_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2089_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2089_a_HPC2_and_n8) );
  XNOR2_X1 cell_2089_a_HPC2_and_U3 ( .A(cell_2089_a_HPC2_and_n7), .B(
        cell_2089_a_HPC2_and_z_0__0_), .ZN(cell_2089_and_out[0]) );
  XNOR2_X1 cell_2089_a_HPC2_and_U2 ( .A(
        cell_2089_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2089_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2089_a_HPC2_and_n7) );
  DFF_X1 cell_2089_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2089_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2089_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2089_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2089_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2089_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2089_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2089_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2089_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2089_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2090_U4 ( .A(signal_3969), .B(cell_2090_and_out[1]), .Z(
        signal_4108) );
  XOR2_X1 cell_2090_U3 ( .A(signal_2323), .B(cell_2090_and_out[0]), .Z(
        signal_2358) );
  XOR2_X1 cell_2090_U2 ( .A(signal_3969), .B(signal_3946), .Z(
        cell_2090_and_in[1]) );
  XOR2_X1 cell_2090_U1 ( .A(signal_2323), .B(signal_2300), .Z(
        cell_2090_and_in[0]) );
  XOR2_X1 cell_2090_a_HPC2_and_U14 ( .A(Fresh[376]), .B(cell_2090_and_in[0]), 
        .Z(cell_2090_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2090_a_HPC2_and_U13 ( .A(Fresh[376]), .B(cell_2090_and_in[1]), 
        .Z(cell_2090_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2090_a_HPC2_and_U12 ( .A1(cell_2090_a_HPC2_and_a_reg[1]), .A2(
        cell_2090_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2090_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2090_a_HPC2_and_U11 ( .A1(cell_2090_a_HPC2_and_a_reg[0]), .A2(
        cell_2090_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2090_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2090_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2090_a_HPC2_and_n9), 
        .ZN(cell_2090_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2090_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2090_a_HPC2_and_n9), 
        .ZN(cell_2090_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2090_a_HPC2_and_U8 ( .A(Fresh[376]), .ZN(cell_2090_a_HPC2_and_n9) );
  AND2_X1 cell_2090_a_HPC2_and_U7 ( .A1(cell_2090_and_in[1]), .A2(n460), .ZN(
        cell_2090_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2090_a_HPC2_and_U6 ( .A1(cell_2090_and_in[0]), .A2(n457), .ZN(
        cell_2090_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2090_a_HPC2_and_U5 ( .A(cell_2090_a_HPC2_and_n8), .B(
        cell_2090_a_HPC2_and_z_1__1_), .ZN(cell_2090_and_out[1]) );
  XNOR2_X1 cell_2090_a_HPC2_and_U4 ( .A(
        cell_2090_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2090_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2090_a_HPC2_and_n8) );
  XNOR2_X1 cell_2090_a_HPC2_and_U3 ( .A(cell_2090_a_HPC2_and_n7), .B(
        cell_2090_a_HPC2_and_z_0__0_), .ZN(cell_2090_and_out[0]) );
  XNOR2_X1 cell_2090_a_HPC2_and_U2 ( .A(
        cell_2090_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2090_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2090_a_HPC2_and_n7) );
  DFF_X1 cell_2090_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2090_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2090_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2090_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2090_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2090_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2090_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2090_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2090_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2090_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2091_U4 ( .A(signal_3963), .B(cell_2091_and_out[1]), .Z(
        signal_4109) );
  XOR2_X1 cell_2091_U3 ( .A(signal_2317), .B(cell_2091_and_out[0]), .Z(
        signal_2359) );
  XOR2_X1 cell_2091_U2 ( .A(signal_3963), .B(signal_3935), .Z(
        cell_2091_and_in[1]) );
  XOR2_X1 cell_2091_U1 ( .A(signal_2317), .B(signal_2289), .Z(
        cell_2091_and_in[0]) );
  XOR2_X1 cell_2091_a_HPC2_and_U14 ( .A(Fresh[377]), .B(cell_2091_and_in[0]), 
        .Z(cell_2091_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2091_a_HPC2_and_U13 ( .A(Fresh[377]), .B(cell_2091_and_in[1]), 
        .Z(cell_2091_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2091_a_HPC2_and_U12 ( .A1(cell_2091_a_HPC2_and_a_reg[1]), .A2(
        cell_2091_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2091_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2091_a_HPC2_and_U11 ( .A1(cell_2091_a_HPC2_and_a_reg[0]), .A2(
        cell_2091_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2091_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2091_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2091_a_HPC2_and_n9), 
        .ZN(cell_2091_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2091_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2091_a_HPC2_and_n9), 
        .ZN(cell_2091_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2091_a_HPC2_and_U8 ( .A(Fresh[377]), .ZN(cell_2091_a_HPC2_and_n9) );
  AND2_X1 cell_2091_a_HPC2_and_U7 ( .A1(cell_2091_and_in[1]), .A2(n460), .ZN(
        cell_2091_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2091_a_HPC2_and_U6 ( .A1(cell_2091_and_in[0]), .A2(n457), .ZN(
        cell_2091_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2091_a_HPC2_and_U5 ( .A(cell_2091_a_HPC2_and_n8), .B(
        cell_2091_a_HPC2_and_z_1__1_), .ZN(cell_2091_and_out[1]) );
  XNOR2_X1 cell_2091_a_HPC2_and_U4 ( .A(
        cell_2091_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2091_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2091_a_HPC2_and_n8) );
  XNOR2_X1 cell_2091_a_HPC2_and_U3 ( .A(cell_2091_a_HPC2_and_n7), .B(
        cell_2091_a_HPC2_and_z_0__0_), .ZN(cell_2091_and_out[0]) );
  XNOR2_X1 cell_2091_a_HPC2_and_U2 ( .A(
        cell_2091_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2091_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2091_a_HPC2_and_n7) );
  DFF_X1 cell_2091_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2091_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2091_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2091_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2091_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2091_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2091_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2091_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2091_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2091_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2092_U4 ( .A(signal_3984), .B(cell_2092_and_out[1]), .Z(
        signal_4110) );
  XOR2_X1 cell_2092_U3 ( .A(signal_2338), .B(cell_2092_and_out[0]), .Z(
        signal_2360) );
  XOR2_X1 cell_2092_U2 ( .A(signal_3984), .B(signal_3982), .Z(
        cell_2092_and_in[1]) );
  XOR2_X1 cell_2092_U1 ( .A(signal_2338), .B(signal_2336), .Z(
        cell_2092_and_in[0]) );
  XOR2_X1 cell_2092_a_HPC2_and_U14 ( .A(Fresh[378]), .B(cell_2092_and_in[0]), 
        .Z(cell_2092_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2092_a_HPC2_and_U13 ( .A(Fresh[378]), .B(cell_2092_and_in[1]), 
        .Z(cell_2092_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2092_a_HPC2_and_U12 ( .A1(cell_2092_a_HPC2_and_a_reg[1]), .A2(
        cell_2092_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2092_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2092_a_HPC2_and_U11 ( .A1(cell_2092_a_HPC2_and_a_reg[0]), .A2(
        cell_2092_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2092_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2092_a_HPC2_and_U10 ( .A1(n460), .A2(cell_2092_a_HPC2_and_n9), 
        .ZN(cell_2092_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2092_a_HPC2_and_U9 ( .A1(n457), .A2(cell_2092_a_HPC2_and_n9), 
        .ZN(cell_2092_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2092_a_HPC2_and_U8 ( .A(Fresh[378]), .ZN(cell_2092_a_HPC2_and_n9) );
  AND2_X1 cell_2092_a_HPC2_and_U7 ( .A1(cell_2092_and_in[1]), .A2(n460), .ZN(
        cell_2092_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2092_a_HPC2_and_U6 ( .A1(cell_2092_and_in[0]), .A2(n457), .ZN(
        cell_2092_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2092_a_HPC2_and_U5 ( .A(cell_2092_a_HPC2_and_n8), .B(
        cell_2092_a_HPC2_and_z_1__1_), .ZN(cell_2092_and_out[1]) );
  XNOR2_X1 cell_2092_a_HPC2_and_U4 ( .A(
        cell_2092_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2092_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2092_a_HPC2_and_n8) );
  XNOR2_X1 cell_2092_a_HPC2_and_U3 ( .A(cell_2092_a_HPC2_and_n7), .B(
        cell_2092_a_HPC2_and_z_0__0_), .ZN(cell_2092_and_out[0]) );
  XNOR2_X1 cell_2092_a_HPC2_and_U2 ( .A(
        cell_2092_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2092_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2092_a_HPC2_and_n7) );
  DFF_X1 cell_2092_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2092_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2092_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n457), .CK(clk), 
        .Q(cell_2092_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2092_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2092_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n460), .CK(clk), 
        .Q(cell_2092_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2092_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2092_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2092_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2093_U4 ( .A(signal_3934), .B(cell_2093_and_out[1]), .Z(
        signal_4111) );
  XOR2_X1 cell_2093_U3 ( .A(signal_2288), .B(cell_2093_and_out[0]), .Z(
        signal_2361) );
  XOR2_X1 cell_2093_U2 ( .A(signal_3934), .B(signal_3976), .Z(
        cell_2093_and_in[1]) );
  XOR2_X1 cell_2093_U1 ( .A(signal_2288), .B(signal_2330), .Z(
        cell_2093_and_in[0]) );
  XOR2_X1 cell_2093_a_HPC2_and_U14 ( .A(Fresh[379]), .B(cell_2093_and_in[0]), 
        .Z(cell_2093_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2093_a_HPC2_and_U13 ( .A(Fresh[379]), .B(cell_2093_and_in[1]), 
        .Z(cell_2093_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2093_a_HPC2_and_U12 ( .A1(cell_2093_a_HPC2_and_a_reg[1]), .A2(
        cell_2093_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2093_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2093_a_HPC2_and_U11 ( .A1(cell_2093_a_HPC2_and_a_reg[0]), .A2(
        cell_2093_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2093_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2093_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2093_a_HPC2_and_n9), 
        .ZN(cell_2093_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2093_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2093_a_HPC2_and_n9), 
        .ZN(cell_2093_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2093_a_HPC2_and_U8 ( .A(Fresh[379]), .ZN(cell_2093_a_HPC2_and_n9) );
  AND2_X1 cell_2093_a_HPC2_and_U7 ( .A1(cell_2093_and_in[1]), .A2(n461), .ZN(
        cell_2093_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2093_a_HPC2_and_U6 ( .A1(cell_2093_and_in[0]), .A2(n458), .ZN(
        cell_2093_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2093_a_HPC2_and_U5 ( .A(cell_2093_a_HPC2_and_n8), .B(
        cell_2093_a_HPC2_and_z_1__1_), .ZN(cell_2093_and_out[1]) );
  XNOR2_X1 cell_2093_a_HPC2_and_U4 ( .A(
        cell_2093_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2093_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2093_a_HPC2_and_n8) );
  XNOR2_X1 cell_2093_a_HPC2_and_U3 ( .A(cell_2093_a_HPC2_and_n7), .B(
        cell_2093_a_HPC2_and_z_0__0_), .ZN(cell_2093_and_out[0]) );
  XNOR2_X1 cell_2093_a_HPC2_and_U2 ( .A(
        cell_2093_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2093_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2093_a_HPC2_and_n7) );
  DFF_X1 cell_2093_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2093_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2093_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2093_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2093_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2093_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2093_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2093_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2093_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2093_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2094_U4 ( .A(signal_3959), .B(cell_2094_and_out[1]), .Z(
        signal_4112) );
  XOR2_X1 cell_2094_U3 ( .A(signal_2313), .B(cell_2094_and_out[0]), .Z(
        signal_2362) );
  XOR2_X1 cell_2094_U2 ( .A(signal_3959), .B(signal_3945), .Z(
        cell_2094_and_in[1]) );
  XOR2_X1 cell_2094_U1 ( .A(signal_2313), .B(signal_2299), .Z(
        cell_2094_and_in[0]) );
  XOR2_X1 cell_2094_a_HPC2_and_U14 ( .A(Fresh[380]), .B(cell_2094_and_in[0]), 
        .Z(cell_2094_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2094_a_HPC2_and_U13 ( .A(Fresh[380]), .B(cell_2094_and_in[1]), 
        .Z(cell_2094_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2094_a_HPC2_and_U12 ( .A1(cell_2094_a_HPC2_and_a_reg[1]), .A2(
        cell_2094_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2094_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2094_a_HPC2_and_U11 ( .A1(cell_2094_a_HPC2_and_a_reg[0]), .A2(
        cell_2094_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2094_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2094_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2094_a_HPC2_and_n9), 
        .ZN(cell_2094_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2094_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2094_a_HPC2_and_n9), 
        .ZN(cell_2094_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2094_a_HPC2_and_U8 ( .A(Fresh[380]), .ZN(cell_2094_a_HPC2_and_n9) );
  AND2_X1 cell_2094_a_HPC2_and_U7 ( .A1(cell_2094_and_in[1]), .A2(n461), .ZN(
        cell_2094_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2094_a_HPC2_and_U6 ( .A1(cell_2094_and_in[0]), .A2(n458), .ZN(
        cell_2094_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2094_a_HPC2_and_U5 ( .A(cell_2094_a_HPC2_and_n8), .B(
        cell_2094_a_HPC2_and_z_1__1_), .ZN(cell_2094_and_out[1]) );
  XNOR2_X1 cell_2094_a_HPC2_and_U4 ( .A(
        cell_2094_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2094_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2094_a_HPC2_and_n8) );
  XNOR2_X1 cell_2094_a_HPC2_and_U3 ( .A(cell_2094_a_HPC2_and_n7), .B(
        cell_2094_a_HPC2_and_z_0__0_), .ZN(cell_2094_and_out[0]) );
  XNOR2_X1 cell_2094_a_HPC2_and_U2 ( .A(
        cell_2094_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2094_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2094_a_HPC2_and_n7) );
  DFF_X1 cell_2094_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2094_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2094_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2094_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2094_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2094_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2094_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2094_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2094_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2094_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2095_U4 ( .A(signal_3952), .B(cell_2095_and_out[1]), .Z(
        signal_4113) );
  XOR2_X1 cell_2095_U3 ( .A(signal_2306), .B(cell_2095_and_out[0]), .Z(
        signal_2363) );
  XOR2_X1 cell_2095_U2 ( .A(signal_3952), .B(signal_3941), .Z(
        cell_2095_and_in[1]) );
  XOR2_X1 cell_2095_U1 ( .A(signal_2306), .B(signal_2295), .Z(
        cell_2095_and_in[0]) );
  XOR2_X1 cell_2095_a_HPC2_and_U14 ( .A(Fresh[381]), .B(cell_2095_and_in[0]), 
        .Z(cell_2095_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2095_a_HPC2_and_U13 ( .A(Fresh[381]), .B(cell_2095_and_in[1]), 
        .Z(cell_2095_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2095_a_HPC2_and_U12 ( .A1(cell_2095_a_HPC2_and_a_reg[1]), .A2(
        cell_2095_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2095_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2095_a_HPC2_and_U11 ( .A1(cell_2095_a_HPC2_and_a_reg[0]), .A2(
        cell_2095_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2095_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2095_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2095_a_HPC2_and_n9), 
        .ZN(cell_2095_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2095_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2095_a_HPC2_and_n9), 
        .ZN(cell_2095_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2095_a_HPC2_and_U8 ( .A(Fresh[381]), .ZN(cell_2095_a_HPC2_and_n9) );
  AND2_X1 cell_2095_a_HPC2_and_U7 ( .A1(cell_2095_and_in[1]), .A2(n461), .ZN(
        cell_2095_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2095_a_HPC2_and_U6 ( .A1(cell_2095_and_in[0]), .A2(n458), .ZN(
        cell_2095_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2095_a_HPC2_and_U5 ( .A(cell_2095_a_HPC2_and_n8), .B(
        cell_2095_a_HPC2_and_z_1__1_), .ZN(cell_2095_and_out[1]) );
  XNOR2_X1 cell_2095_a_HPC2_and_U4 ( .A(
        cell_2095_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2095_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2095_a_HPC2_and_n8) );
  XNOR2_X1 cell_2095_a_HPC2_and_U3 ( .A(cell_2095_a_HPC2_and_n7), .B(
        cell_2095_a_HPC2_and_z_0__0_), .ZN(cell_2095_and_out[0]) );
  XNOR2_X1 cell_2095_a_HPC2_and_U2 ( .A(
        cell_2095_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2095_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2095_a_HPC2_and_n7) );
  DFF_X1 cell_2095_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2095_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2095_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2095_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2095_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2095_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2095_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2095_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2095_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2095_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2096_U4 ( .A(signal_3923), .B(cell_2096_and_out[1]), .Z(
        signal_4114) );
  XOR2_X1 cell_2096_U3 ( .A(signal_2277), .B(cell_2096_and_out[0]), .Z(
        signal_2364) );
  XOR2_X1 cell_2096_U2 ( .A(signal_3923), .B(signal_3948), .Z(
        cell_2096_and_in[1]) );
  XOR2_X1 cell_2096_U1 ( .A(signal_2277), .B(signal_2302), .Z(
        cell_2096_and_in[0]) );
  XOR2_X1 cell_2096_a_HPC2_and_U14 ( .A(Fresh[382]), .B(cell_2096_and_in[0]), 
        .Z(cell_2096_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2096_a_HPC2_and_U13 ( .A(Fresh[382]), .B(cell_2096_and_in[1]), 
        .Z(cell_2096_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2096_a_HPC2_and_U12 ( .A1(cell_2096_a_HPC2_and_a_reg[1]), .A2(
        cell_2096_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2096_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2096_a_HPC2_and_U11 ( .A1(cell_2096_a_HPC2_and_a_reg[0]), .A2(
        cell_2096_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2096_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2096_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2096_a_HPC2_and_n9), 
        .ZN(cell_2096_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2096_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2096_a_HPC2_and_n9), 
        .ZN(cell_2096_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2096_a_HPC2_and_U8 ( .A(Fresh[382]), .ZN(cell_2096_a_HPC2_and_n9) );
  AND2_X1 cell_2096_a_HPC2_and_U7 ( .A1(cell_2096_and_in[1]), .A2(n461), .ZN(
        cell_2096_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2096_a_HPC2_and_U6 ( .A1(cell_2096_and_in[0]), .A2(n458), .ZN(
        cell_2096_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2096_a_HPC2_and_U5 ( .A(cell_2096_a_HPC2_and_n8), .B(
        cell_2096_a_HPC2_and_z_1__1_), .ZN(cell_2096_and_out[1]) );
  XNOR2_X1 cell_2096_a_HPC2_and_U4 ( .A(
        cell_2096_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2096_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2096_a_HPC2_and_n8) );
  XNOR2_X1 cell_2096_a_HPC2_and_U3 ( .A(cell_2096_a_HPC2_and_n7), .B(
        cell_2096_a_HPC2_and_z_0__0_), .ZN(cell_2096_and_out[0]) );
  XNOR2_X1 cell_2096_a_HPC2_and_U2 ( .A(
        cell_2096_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2096_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2096_a_HPC2_and_n7) );
  DFF_X1 cell_2096_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2096_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2096_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2096_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2096_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2096_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2096_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2096_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2096_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2096_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2097_U4 ( .A(signal_3954), .B(cell_2097_and_out[1]), .Z(
        signal_4115) );
  XOR2_X1 cell_2097_U3 ( .A(signal_2308), .B(cell_2097_and_out[0]), .Z(
        signal_2365) );
  XOR2_X1 cell_2097_U2 ( .A(signal_3954), .B(signal_3967), .Z(
        cell_2097_and_in[1]) );
  XOR2_X1 cell_2097_U1 ( .A(signal_2308), .B(signal_2321), .Z(
        cell_2097_and_in[0]) );
  XOR2_X1 cell_2097_a_HPC2_and_U14 ( .A(Fresh[383]), .B(cell_2097_and_in[0]), 
        .Z(cell_2097_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2097_a_HPC2_and_U13 ( .A(Fresh[383]), .B(cell_2097_and_in[1]), 
        .Z(cell_2097_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2097_a_HPC2_and_U12 ( .A1(cell_2097_a_HPC2_and_a_reg[1]), .A2(
        cell_2097_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2097_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2097_a_HPC2_and_U11 ( .A1(cell_2097_a_HPC2_and_a_reg[0]), .A2(
        cell_2097_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2097_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2097_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2097_a_HPC2_and_n9), 
        .ZN(cell_2097_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2097_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2097_a_HPC2_and_n9), 
        .ZN(cell_2097_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2097_a_HPC2_and_U8 ( .A(Fresh[383]), .ZN(cell_2097_a_HPC2_and_n9) );
  AND2_X1 cell_2097_a_HPC2_and_U7 ( .A1(cell_2097_and_in[1]), .A2(n461), .ZN(
        cell_2097_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2097_a_HPC2_and_U6 ( .A1(cell_2097_and_in[0]), .A2(n458), .ZN(
        cell_2097_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2097_a_HPC2_and_U5 ( .A(cell_2097_a_HPC2_and_n8), .B(
        cell_2097_a_HPC2_and_z_1__1_), .ZN(cell_2097_and_out[1]) );
  XNOR2_X1 cell_2097_a_HPC2_and_U4 ( .A(
        cell_2097_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2097_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2097_a_HPC2_and_n8) );
  XNOR2_X1 cell_2097_a_HPC2_and_U3 ( .A(cell_2097_a_HPC2_and_n7), .B(
        cell_2097_a_HPC2_and_z_0__0_), .ZN(cell_2097_and_out[0]) );
  XNOR2_X1 cell_2097_a_HPC2_and_U2 ( .A(
        cell_2097_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2097_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2097_a_HPC2_and_n7) );
  DFF_X1 cell_2097_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2097_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2097_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2097_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2097_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2097_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2097_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2097_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2097_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2097_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2098_U4 ( .A(signal_3965), .B(cell_2098_and_out[1]), .Z(
        signal_4116) );
  XOR2_X1 cell_2098_U3 ( .A(signal_2319), .B(cell_2098_and_out[0]), .Z(
        signal_2366) );
  XOR2_X1 cell_2098_U2 ( .A(signal_3965), .B(signal_3950), .Z(
        cell_2098_and_in[1]) );
  XOR2_X1 cell_2098_U1 ( .A(signal_2319), .B(signal_2304), .Z(
        cell_2098_and_in[0]) );
  XOR2_X1 cell_2098_a_HPC2_and_U14 ( .A(Fresh[384]), .B(cell_2098_and_in[0]), 
        .Z(cell_2098_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2098_a_HPC2_and_U13 ( .A(Fresh[384]), .B(cell_2098_and_in[1]), 
        .Z(cell_2098_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2098_a_HPC2_and_U12 ( .A1(cell_2098_a_HPC2_and_a_reg[1]), .A2(
        cell_2098_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2098_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2098_a_HPC2_and_U11 ( .A1(cell_2098_a_HPC2_and_a_reg[0]), .A2(
        cell_2098_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2098_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2098_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2098_a_HPC2_and_n9), 
        .ZN(cell_2098_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2098_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2098_a_HPC2_and_n9), 
        .ZN(cell_2098_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2098_a_HPC2_and_U8 ( .A(Fresh[384]), .ZN(cell_2098_a_HPC2_and_n9) );
  AND2_X1 cell_2098_a_HPC2_and_U7 ( .A1(cell_2098_and_in[1]), .A2(n461), .ZN(
        cell_2098_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2098_a_HPC2_and_U6 ( .A1(cell_2098_and_in[0]), .A2(n458), .ZN(
        cell_2098_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2098_a_HPC2_and_U5 ( .A(cell_2098_a_HPC2_and_n8), .B(
        cell_2098_a_HPC2_and_z_1__1_), .ZN(cell_2098_and_out[1]) );
  XNOR2_X1 cell_2098_a_HPC2_and_U4 ( .A(
        cell_2098_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2098_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2098_a_HPC2_and_n8) );
  XNOR2_X1 cell_2098_a_HPC2_and_U3 ( .A(cell_2098_a_HPC2_and_n7), .B(
        cell_2098_a_HPC2_and_z_0__0_), .ZN(cell_2098_and_out[0]) );
  XNOR2_X1 cell_2098_a_HPC2_and_U2 ( .A(
        cell_2098_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2098_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2098_a_HPC2_and_n7) );
  DFF_X1 cell_2098_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2098_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2098_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2098_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2098_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2098_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2098_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2098_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2098_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2098_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2099_U4 ( .A(signal_3943), .B(cell_2099_and_out[1]), .Z(
        signal_4117) );
  XOR2_X1 cell_2099_U3 ( .A(signal_2297), .B(cell_2099_and_out[0]), .Z(
        signal_2367) );
  XOR2_X1 cell_2099_U2 ( .A(signal_3943), .B(signal_3957), .Z(
        cell_2099_and_in[1]) );
  XOR2_X1 cell_2099_U1 ( .A(signal_2297), .B(signal_2311), .Z(
        cell_2099_and_in[0]) );
  XOR2_X1 cell_2099_a_HPC2_and_U14 ( .A(Fresh[385]), .B(cell_2099_and_in[0]), 
        .Z(cell_2099_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2099_a_HPC2_and_U13 ( .A(Fresh[385]), .B(cell_2099_and_in[1]), 
        .Z(cell_2099_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2099_a_HPC2_and_U12 ( .A1(cell_2099_a_HPC2_and_a_reg[1]), .A2(
        cell_2099_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2099_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2099_a_HPC2_and_U11 ( .A1(cell_2099_a_HPC2_and_a_reg[0]), .A2(
        cell_2099_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2099_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2099_a_HPC2_and_U10 ( .A1(n461), .A2(cell_2099_a_HPC2_and_n9), 
        .ZN(cell_2099_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2099_a_HPC2_and_U9 ( .A1(n458), .A2(cell_2099_a_HPC2_and_n9), 
        .ZN(cell_2099_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2099_a_HPC2_and_U8 ( .A(Fresh[385]), .ZN(cell_2099_a_HPC2_and_n9) );
  AND2_X1 cell_2099_a_HPC2_and_U7 ( .A1(cell_2099_and_in[1]), .A2(n461), .ZN(
        cell_2099_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2099_a_HPC2_and_U6 ( .A1(cell_2099_and_in[0]), .A2(n458), .ZN(
        cell_2099_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2099_a_HPC2_and_U5 ( .A(cell_2099_a_HPC2_and_n8), .B(
        cell_2099_a_HPC2_and_z_1__1_), .ZN(cell_2099_and_out[1]) );
  XNOR2_X1 cell_2099_a_HPC2_and_U4 ( .A(
        cell_2099_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2099_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2099_a_HPC2_and_n8) );
  XNOR2_X1 cell_2099_a_HPC2_and_U3 ( .A(cell_2099_a_HPC2_and_n7), .B(
        cell_2099_a_HPC2_and_z_0__0_), .ZN(cell_2099_and_out[0]) );
  XNOR2_X1 cell_2099_a_HPC2_and_U2 ( .A(
        cell_2099_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2099_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2099_a_HPC2_and_n7) );
  DFF_X1 cell_2099_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2099_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2099_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n458), .CK(clk), 
        .Q(cell_2099_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2099_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2099_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n461), .CK(clk), 
        .Q(cell_2099_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2099_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2099_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2099_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2100_U4 ( .A(signal_3940), .B(cell_2100_and_out[1]), .Z(
        signal_4118) );
  XOR2_X1 cell_2100_U3 ( .A(signal_2294), .B(cell_2100_and_out[0]), .Z(
        signal_2368) );
  XOR2_X1 cell_2100_U2 ( .A(signal_3940), .B(signal_3932), .Z(
        cell_2100_and_in[1]) );
  XOR2_X1 cell_2100_U1 ( .A(signal_2294), .B(signal_2286), .Z(
        cell_2100_and_in[0]) );
  XOR2_X1 cell_2100_a_HPC2_and_U14 ( .A(Fresh[386]), .B(cell_2100_and_in[0]), 
        .Z(cell_2100_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2100_a_HPC2_and_U13 ( .A(Fresh[386]), .B(cell_2100_and_in[1]), 
        .Z(cell_2100_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2100_a_HPC2_and_U12 ( .A1(cell_2100_a_HPC2_and_a_reg[1]), .A2(
        cell_2100_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2100_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2100_a_HPC2_and_U11 ( .A1(cell_2100_a_HPC2_and_a_reg[0]), .A2(
        cell_2100_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2100_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2100_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2100_a_HPC2_and_n9), .ZN(cell_2100_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2100_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2100_a_HPC2_and_n9), .ZN(cell_2100_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2100_a_HPC2_and_U8 ( .A(Fresh[386]), .ZN(cell_2100_a_HPC2_and_n9) );
  AND2_X1 cell_2100_a_HPC2_and_U7 ( .A1(cell_2100_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2100_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2100_a_HPC2_and_U6 ( .A1(cell_2100_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2100_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2100_a_HPC2_and_U5 ( .A(cell_2100_a_HPC2_and_n8), .B(
        cell_2100_a_HPC2_and_z_1__1_), .ZN(cell_2100_and_out[1]) );
  XNOR2_X1 cell_2100_a_HPC2_and_U4 ( .A(
        cell_2100_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2100_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2100_a_HPC2_and_n8) );
  XNOR2_X1 cell_2100_a_HPC2_and_U3 ( .A(cell_2100_a_HPC2_and_n7), .B(
        cell_2100_a_HPC2_and_z_0__0_), .ZN(cell_2100_and_out[0]) );
  XNOR2_X1 cell_2100_a_HPC2_and_U2 ( .A(
        cell_2100_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2100_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2100_a_HPC2_and_n7) );
  DFF_X1 cell_2100_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2100_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2100_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2100_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2100_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2100_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2100_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2100_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2100_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2100_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2101_U4 ( .A(signal_3955), .B(cell_2101_and_out[1]), .Z(
        signal_4119) );
  XOR2_X1 cell_2101_U3 ( .A(signal_2309), .B(cell_2101_and_out[0]), .Z(
        signal_2369) );
  XOR2_X1 cell_2101_U2 ( .A(signal_3955), .B(signal_3953), .Z(
        cell_2101_and_in[1]) );
  XOR2_X1 cell_2101_U1 ( .A(signal_2309), .B(signal_2307), .Z(
        cell_2101_and_in[0]) );
  XOR2_X1 cell_2101_a_HPC2_and_U14 ( .A(Fresh[387]), .B(cell_2101_and_in[0]), 
        .Z(cell_2101_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2101_a_HPC2_and_U13 ( .A(Fresh[387]), .B(cell_2101_and_in[1]), 
        .Z(cell_2101_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2101_a_HPC2_and_U12 ( .A1(cell_2101_a_HPC2_and_a_reg[1]), .A2(
        cell_2101_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2101_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2101_a_HPC2_and_U11 ( .A1(cell_2101_a_HPC2_and_a_reg[0]), .A2(
        cell_2101_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2101_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2101_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2101_a_HPC2_and_n9), .ZN(cell_2101_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2101_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2101_a_HPC2_and_n9), .ZN(cell_2101_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2101_a_HPC2_and_U8 ( .A(Fresh[387]), .ZN(cell_2101_a_HPC2_and_n9) );
  AND2_X1 cell_2101_a_HPC2_and_U7 ( .A1(cell_2101_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2101_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2101_a_HPC2_and_U6 ( .A1(cell_2101_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2101_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2101_a_HPC2_and_U5 ( .A(cell_2101_a_HPC2_and_n8), .B(
        cell_2101_a_HPC2_and_z_1__1_), .ZN(cell_2101_and_out[1]) );
  XNOR2_X1 cell_2101_a_HPC2_and_U4 ( .A(
        cell_2101_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2101_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2101_a_HPC2_and_n8) );
  XNOR2_X1 cell_2101_a_HPC2_and_U3 ( .A(cell_2101_a_HPC2_and_n7), .B(
        cell_2101_a_HPC2_and_z_0__0_), .ZN(cell_2101_and_out[0]) );
  XNOR2_X1 cell_2101_a_HPC2_and_U2 ( .A(
        cell_2101_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2101_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2101_a_HPC2_and_n7) );
  DFF_X1 cell_2101_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2101_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2101_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2101_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2101_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2101_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2101_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2101_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2101_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2101_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2102_U4 ( .A(signal_3925), .B(cell_2102_and_out[1]), .Z(
        signal_4120) );
  XOR2_X1 cell_2102_U3 ( .A(signal_2279), .B(cell_2102_and_out[0]), .Z(
        signal_2370) );
  XOR2_X1 cell_2102_U2 ( .A(signal_3925), .B(signal_3973), .Z(
        cell_2102_and_in[1]) );
  XOR2_X1 cell_2102_U1 ( .A(signal_2279), .B(signal_2327), .Z(
        cell_2102_and_in[0]) );
  XOR2_X1 cell_2102_a_HPC2_and_U14 ( .A(Fresh[388]), .B(cell_2102_and_in[0]), 
        .Z(cell_2102_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2102_a_HPC2_and_U13 ( .A(Fresh[388]), .B(cell_2102_and_in[1]), 
        .Z(cell_2102_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2102_a_HPC2_and_U12 ( .A1(cell_2102_a_HPC2_and_a_reg[1]), .A2(
        cell_2102_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2102_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2102_a_HPC2_and_U11 ( .A1(cell_2102_a_HPC2_and_a_reg[0]), .A2(
        cell_2102_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2102_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2102_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2102_a_HPC2_and_n9), .ZN(cell_2102_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2102_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2102_a_HPC2_and_n9), .ZN(cell_2102_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2102_a_HPC2_and_U8 ( .A(Fresh[388]), .ZN(cell_2102_a_HPC2_and_n9) );
  AND2_X1 cell_2102_a_HPC2_and_U7 ( .A1(cell_2102_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2102_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2102_a_HPC2_and_U6 ( .A1(cell_2102_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2102_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2102_a_HPC2_and_U5 ( .A(cell_2102_a_HPC2_and_n8), .B(
        cell_2102_a_HPC2_and_z_1__1_), .ZN(cell_2102_and_out[1]) );
  XNOR2_X1 cell_2102_a_HPC2_and_U4 ( .A(
        cell_2102_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2102_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2102_a_HPC2_and_n8) );
  XNOR2_X1 cell_2102_a_HPC2_and_U3 ( .A(cell_2102_a_HPC2_and_n7), .B(
        cell_2102_a_HPC2_and_z_0__0_), .ZN(cell_2102_and_out[0]) );
  XNOR2_X1 cell_2102_a_HPC2_and_U2 ( .A(
        cell_2102_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2102_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2102_a_HPC2_and_n7) );
  DFF_X1 cell_2102_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2102_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2102_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2102_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2102_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2102_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2102_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2102_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2102_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2102_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2103_U4 ( .A(signal_3977), .B(cell_2103_and_out[1]), .Z(
        signal_4121) );
  XOR2_X1 cell_2103_U3 ( .A(signal_2331), .B(cell_2103_and_out[0]), .Z(
        signal_2371) );
  XOR2_X1 cell_2103_U2 ( .A(signal_3977), .B(signal_3962), .Z(
        cell_2103_and_in[1]) );
  XOR2_X1 cell_2103_U1 ( .A(signal_2331), .B(signal_2316), .Z(
        cell_2103_and_in[0]) );
  XOR2_X1 cell_2103_a_HPC2_and_U14 ( .A(Fresh[389]), .B(cell_2103_and_in[0]), 
        .Z(cell_2103_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2103_a_HPC2_and_U13 ( .A(Fresh[389]), .B(cell_2103_and_in[1]), 
        .Z(cell_2103_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2103_a_HPC2_and_U12 ( .A1(cell_2103_a_HPC2_and_a_reg[1]), .A2(
        cell_2103_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2103_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2103_a_HPC2_and_U11 ( .A1(cell_2103_a_HPC2_and_a_reg[0]), .A2(
        cell_2103_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2103_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2103_a_HPC2_and_U10 ( .A1(signal_3234), .A2(
        cell_2103_a_HPC2_and_n9), .ZN(cell_2103_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2103_a_HPC2_and_U9 ( .A1(signal_1515), .A2(
        cell_2103_a_HPC2_and_n9), .ZN(cell_2103_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2103_a_HPC2_and_U8 ( .A(Fresh[389]), .ZN(cell_2103_a_HPC2_and_n9) );
  AND2_X1 cell_2103_a_HPC2_and_U7 ( .A1(cell_2103_and_in[1]), .A2(signal_3234), 
        .ZN(cell_2103_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2103_a_HPC2_and_U6 ( .A1(cell_2103_and_in[0]), .A2(signal_1515), 
        .ZN(cell_2103_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2103_a_HPC2_and_U5 ( .A(cell_2103_a_HPC2_and_n8), .B(
        cell_2103_a_HPC2_and_z_1__1_), .ZN(cell_2103_and_out[1]) );
  XNOR2_X1 cell_2103_a_HPC2_and_U4 ( .A(
        cell_2103_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2103_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2103_a_HPC2_and_n8) );
  XNOR2_X1 cell_2103_a_HPC2_and_U3 ( .A(cell_2103_a_HPC2_and_n7), .B(
        cell_2103_a_HPC2_and_z_0__0_), .ZN(cell_2103_and_out[0]) );
  XNOR2_X1 cell_2103_a_HPC2_and_U2 ( .A(
        cell_2103_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2103_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2103_a_HPC2_and_n7) );
  DFF_X1 cell_2103_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2103_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2103_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1515), 
        .CK(clk), .Q(cell_2103_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2103_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2103_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3234), 
        .CK(clk), .Q(cell_2103_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2103_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2103_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2103_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2104_U4 ( .A(signal_4119), .B(cell_2104_and_out[1]), .Z(
        signal_4130) );
  XOR2_X1 cell_2104_U3 ( .A(signal_2369), .B(cell_2104_and_out[0]), .Z(
        signal_2372) );
  XOR2_X1 cell_2104_U2 ( .A(signal_4119), .B(signal_4111), .Z(
        cell_2104_and_in[1]) );
  XOR2_X1 cell_2104_U1 ( .A(signal_2369), .B(signal_2361), .Z(
        cell_2104_and_in[0]) );
  XOR2_X1 cell_2104_a_HPC2_and_U14 ( .A(Fresh[390]), .B(cell_2104_and_in[0]), 
        .Z(cell_2104_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2104_a_HPC2_and_U13 ( .A(Fresh[390]), .B(cell_2104_and_in[1]), 
        .Z(cell_2104_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2104_a_HPC2_and_U12 ( .A1(cell_2104_a_HPC2_and_a_reg[1]), .A2(
        cell_2104_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2104_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2104_a_HPC2_and_U11 ( .A1(cell_2104_a_HPC2_and_a_reg[0]), .A2(
        cell_2104_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2104_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2104_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2104_a_HPC2_and_n9), .ZN(cell_2104_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2104_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2104_a_HPC2_and_n9), .ZN(cell_2104_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2104_a_HPC2_and_U8 ( .A(Fresh[390]), .ZN(cell_2104_a_HPC2_and_n9) );
  AND2_X1 cell_2104_a_HPC2_and_U7 ( .A1(cell_2104_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2104_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2104_a_HPC2_and_U6 ( .A1(cell_2104_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2104_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2104_a_HPC2_and_U5 ( .A(cell_2104_a_HPC2_and_n8), .B(
        cell_2104_a_HPC2_and_z_1__1_), .ZN(cell_2104_and_out[1]) );
  XNOR2_X1 cell_2104_a_HPC2_and_U4 ( .A(
        cell_2104_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2104_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2104_a_HPC2_and_n8) );
  XNOR2_X1 cell_2104_a_HPC2_and_U3 ( .A(cell_2104_a_HPC2_and_n7), .B(
        cell_2104_a_HPC2_and_z_0__0_), .ZN(cell_2104_and_out[0]) );
  XNOR2_X1 cell_2104_a_HPC2_and_U2 ( .A(
        cell_2104_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2104_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2104_a_HPC2_and_n7) );
  DFF_X1 cell_2104_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2104_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2104_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2104_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2104_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2104_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2104_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2104_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2104_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2104_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2105_U4 ( .A(signal_4099), .B(cell_2105_and_out[1]), .Z(
        signal_4131) );
  XOR2_X1 cell_2105_U3 ( .A(signal_2349), .B(cell_2105_and_out[0]), .Z(
        signal_2373) );
  XOR2_X1 cell_2105_U2 ( .A(signal_4099), .B(signal_4091), .Z(
        cell_2105_and_in[1]) );
  XOR2_X1 cell_2105_U1 ( .A(signal_2349), .B(signal_2341), .Z(
        cell_2105_and_in[0]) );
  XOR2_X1 cell_2105_a_HPC2_and_U14 ( .A(Fresh[391]), .B(cell_2105_and_in[0]), 
        .Z(cell_2105_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2105_a_HPC2_and_U13 ( .A(Fresh[391]), .B(cell_2105_and_in[1]), 
        .Z(cell_2105_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2105_a_HPC2_and_U12 ( .A1(cell_2105_a_HPC2_and_a_reg[1]), .A2(
        cell_2105_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2105_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2105_a_HPC2_and_U11 ( .A1(cell_2105_a_HPC2_and_a_reg[0]), .A2(
        cell_2105_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2105_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2105_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2105_a_HPC2_and_n9), .ZN(cell_2105_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2105_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2105_a_HPC2_and_n9), .ZN(cell_2105_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2105_a_HPC2_and_U8 ( .A(Fresh[391]), .ZN(cell_2105_a_HPC2_and_n9) );
  AND2_X1 cell_2105_a_HPC2_and_U7 ( .A1(cell_2105_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2105_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2105_a_HPC2_and_U6 ( .A1(cell_2105_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2105_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2105_a_HPC2_and_U5 ( .A(cell_2105_a_HPC2_and_n8), .B(
        cell_2105_a_HPC2_and_z_1__1_), .ZN(cell_2105_and_out[1]) );
  XNOR2_X1 cell_2105_a_HPC2_and_U4 ( .A(
        cell_2105_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2105_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2105_a_HPC2_and_n8) );
  XNOR2_X1 cell_2105_a_HPC2_and_U3 ( .A(cell_2105_a_HPC2_and_n7), .B(
        cell_2105_a_HPC2_and_z_0__0_), .ZN(cell_2105_and_out[0]) );
  XNOR2_X1 cell_2105_a_HPC2_and_U2 ( .A(
        cell_2105_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2105_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2105_a_HPC2_and_n7) );
  DFF_X1 cell_2105_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2105_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2105_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2105_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2105_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2105_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2105_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2105_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2105_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2105_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2106_U4 ( .A(signal_4114), .B(cell_2106_and_out[1]), .Z(
        signal_4132) );
  XOR2_X1 cell_2106_U3 ( .A(signal_2364), .B(cell_2106_and_out[0]), .Z(
        signal_2374) );
  XOR2_X1 cell_2106_U2 ( .A(signal_4114), .B(signal_4121), .Z(
        cell_2106_and_in[1]) );
  XOR2_X1 cell_2106_U1 ( .A(signal_2364), .B(signal_2371), .Z(
        cell_2106_and_in[0]) );
  XOR2_X1 cell_2106_a_HPC2_and_U14 ( .A(Fresh[392]), .B(cell_2106_and_in[0]), 
        .Z(cell_2106_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2106_a_HPC2_and_U13 ( .A(Fresh[392]), .B(cell_2106_and_in[1]), 
        .Z(cell_2106_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2106_a_HPC2_and_U12 ( .A1(cell_2106_a_HPC2_and_a_reg[1]), .A2(
        cell_2106_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2106_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2106_a_HPC2_and_U11 ( .A1(cell_2106_a_HPC2_and_a_reg[0]), .A2(
        cell_2106_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2106_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2106_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2106_a_HPC2_and_n9), .ZN(cell_2106_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2106_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2106_a_HPC2_and_n9), .ZN(cell_2106_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2106_a_HPC2_and_U8 ( .A(Fresh[392]), .ZN(cell_2106_a_HPC2_and_n9) );
  AND2_X1 cell_2106_a_HPC2_and_U7 ( .A1(cell_2106_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2106_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2106_a_HPC2_and_U6 ( .A1(cell_2106_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2106_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2106_a_HPC2_and_U5 ( .A(cell_2106_a_HPC2_and_n8), .B(
        cell_2106_a_HPC2_and_z_1__1_), .ZN(cell_2106_and_out[1]) );
  XNOR2_X1 cell_2106_a_HPC2_and_U4 ( .A(
        cell_2106_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2106_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2106_a_HPC2_and_n8) );
  XNOR2_X1 cell_2106_a_HPC2_and_U3 ( .A(cell_2106_a_HPC2_and_n7), .B(
        cell_2106_a_HPC2_and_z_0__0_), .ZN(cell_2106_and_out[0]) );
  XNOR2_X1 cell_2106_a_HPC2_and_U2 ( .A(
        cell_2106_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2106_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2106_a_HPC2_and_n7) );
  DFF_X1 cell_2106_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2106_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2106_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2106_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2106_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2106_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2106_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2106_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2106_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2106_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2107_U4 ( .A(signal_4118), .B(cell_2107_and_out[1]), .Z(
        signal_4133) );
  XOR2_X1 cell_2107_U3 ( .A(signal_2368), .B(cell_2107_and_out[0]), .Z(
        signal_2375) );
  XOR2_X1 cell_2107_U2 ( .A(signal_4118), .B(signal_4100), .Z(
        cell_2107_and_in[1]) );
  XOR2_X1 cell_2107_U1 ( .A(signal_2368), .B(signal_2350), .Z(
        cell_2107_and_in[0]) );
  XOR2_X1 cell_2107_a_HPC2_and_U14 ( .A(Fresh[393]), .B(cell_2107_and_in[0]), 
        .Z(cell_2107_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2107_a_HPC2_and_U13 ( .A(Fresh[393]), .B(cell_2107_and_in[1]), 
        .Z(cell_2107_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2107_a_HPC2_and_U12 ( .A1(cell_2107_a_HPC2_and_a_reg[1]), .A2(
        cell_2107_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2107_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2107_a_HPC2_and_U11 ( .A1(cell_2107_a_HPC2_and_a_reg[0]), .A2(
        cell_2107_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2107_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2107_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2107_a_HPC2_and_n9), .ZN(cell_2107_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2107_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2107_a_HPC2_and_n9), .ZN(cell_2107_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2107_a_HPC2_and_U8 ( .A(Fresh[393]), .ZN(cell_2107_a_HPC2_and_n9) );
  AND2_X1 cell_2107_a_HPC2_and_U7 ( .A1(cell_2107_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2107_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2107_a_HPC2_and_U6 ( .A1(cell_2107_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2107_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2107_a_HPC2_and_U5 ( .A(cell_2107_a_HPC2_and_n8), .B(
        cell_2107_a_HPC2_and_z_1__1_), .ZN(cell_2107_and_out[1]) );
  XNOR2_X1 cell_2107_a_HPC2_and_U4 ( .A(
        cell_2107_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2107_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2107_a_HPC2_and_n8) );
  XNOR2_X1 cell_2107_a_HPC2_and_U3 ( .A(cell_2107_a_HPC2_and_n7), .B(
        cell_2107_a_HPC2_and_z_0__0_), .ZN(cell_2107_and_out[0]) );
  XNOR2_X1 cell_2107_a_HPC2_and_U2 ( .A(
        cell_2107_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2107_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2107_a_HPC2_and_n7) );
  DFF_X1 cell_2107_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2107_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2107_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2107_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2107_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2107_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2107_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2107_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2107_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2107_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2108_U4 ( .A(signal_4109), .B(cell_2108_and_out[1]), .Z(
        signal_4134) );
  XOR2_X1 cell_2108_U3 ( .A(signal_2359), .B(cell_2108_and_out[0]), .Z(
        signal_2376) );
  XOR2_X1 cell_2108_U2 ( .A(signal_4109), .B(signal_4094), .Z(
        cell_2108_and_in[1]) );
  XOR2_X1 cell_2108_U1 ( .A(signal_2359), .B(signal_2344), .Z(
        cell_2108_and_in[0]) );
  XOR2_X1 cell_2108_a_HPC2_and_U14 ( .A(Fresh[394]), .B(cell_2108_and_in[0]), 
        .Z(cell_2108_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2108_a_HPC2_and_U13 ( .A(Fresh[394]), .B(cell_2108_and_in[1]), 
        .Z(cell_2108_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2108_a_HPC2_and_U12 ( .A1(cell_2108_a_HPC2_and_a_reg[1]), .A2(
        cell_2108_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2108_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2108_a_HPC2_and_U11 ( .A1(cell_2108_a_HPC2_and_a_reg[0]), .A2(
        cell_2108_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2108_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2108_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2108_a_HPC2_and_n9), .ZN(cell_2108_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2108_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2108_a_HPC2_and_n9), .ZN(cell_2108_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2108_a_HPC2_and_U8 ( .A(Fresh[394]), .ZN(cell_2108_a_HPC2_and_n9) );
  AND2_X1 cell_2108_a_HPC2_and_U7 ( .A1(cell_2108_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2108_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2108_a_HPC2_and_U6 ( .A1(cell_2108_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2108_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2108_a_HPC2_and_U5 ( .A(cell_2108_a_HPC2_and_n8), .B(
        cell_2108_a_HPC2_and_z_1__1_), .ZN(cell_2108_and_out[1]) );
  XNOR2_X1 cell_2108_a_HPC2_and_U4 ( .A(
        cell_2108_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2108_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2108_a_HPC2_and_n8) );
  XNOR2_X1 cell_2108_a_HPC2_and_U3 ( .A(cell_2108_a_HPC2_and_n7), .B(
        cell_2108_a_HPC2_and_z_0__0_), .ZN(cell_2108_and_out[0]) );
  XNOR2_X1 cell_2108_a_HPC2_and_U2 ( .A(
        cell_2108_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2108_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2108_a_HPC2_and_n7) );
  DFF_X1 cell_2108_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2108_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2108_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2108_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2108_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2108_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2108_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2108_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2108_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2108_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2109_U4 ( .A(signal_4092), .B(cell_2109_and_out[1]), .Z(
        signal_4135) );
  XOR2_X1 cell_2109_U3 ( .A(signal_2342), .B(cell_2109_and_out[0]), .Z(
        signal_2377) );
  XOR2_X1 cell_2109_U2 ( .A(signal_4092), .B(signal_4102), .Z(
        cell_2109_and_in[1]) );
  XOR2_X1 cell_2109_U1 ( .A(signal_2342), .B(signal_2352), .Z(
        cell_2109_and_in[0]) );
  XOR2_X1 cell_2109_a_HPC2_and_U14 ( .A(Fresh[395]), .B(cell_2109_and_in[0]), 
        .Z(cell_2109_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2109_a_HPC2_and_U13 ( .A(Fresh[395]), .B(cell_2109_and_in[1]), 
        .Z(cell_2109_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2109_a_HPC2_and_U12 ( .A1(cell_2109_a_HPC2_and_a_reg[1]), .A2(
        cell_2109_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2109_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2109_a_HPC2_and_U11 ( .A1(cell_2109_a_HPC2_and_a_reg[0]), .A2(
        cell_2109_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2109_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2109_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2109_a_HPC2_and_n9), .ZN(cell_2109_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2109_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2109_a_HPC2_and_n9), .ZN(cell_2109_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2109_a_HPC2_and_U8 ( .A(Fresh[395]), .ZN(cell_2109_a_HPC2_and_n9) );
  AND2_X1 cell_2109_a_HPC2_and_U7 ( .A1(cell_2109_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2109_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2109_a_HPC2_and_U6 ( .A1(cell_2109_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2109_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2109_a_HPC2_and_U5 ( .A(cell_2109_a_HPC2_and_n8), .B(
        cell_2109_a_HPC2_and_z_1__1_), .ZN(cell_2109_and_out[1]) );
  XNOR2_X1 cell_2109_a_HPC2_and_U4 ( .A(
        cell_2109_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2109_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2109_a_HPC2_and_n8) );
  XNOR2_X1 cell_2109_a_HPC2_and_U3 ( .A(cell_2109_a_HPC2_and_n7), .B(
        cell_2109_a_HPC2_and_z_0__0_), .ZN(cell_2109_and_out[0]) );
  XNOR2_X1 cell_2109_a_HPC2_and_U2 ( .A(
        cell_2109_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2109_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2109_a_HPC2_and_n7) );
  DFF_X1 cell_2109_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2109_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2109_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2109_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2109_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2109_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2109_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2109_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2109_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2109_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2110_U4 ( .A(signal_4098), .B(cell_2110_and_out[1]), .Z(
        signal_4136) );
  XOR2_X1 cell_2110_U3 ( .A(signal_2348), .B(cell_2110_and_out[0]), .Z(
        signal_2378) );
  XOR2_X1 cell_2110_U2 ( .A(signal_4098), .B(signal_4108), .Z(
        cell_2110_and_in[1]) );
  XOR2_X1 cell_2110_U1 ( .A(signal_2348), .B(signal_2358), .Z(
        cell_2110_and_in[0]) );
  XOR2_X1 cell_2110_a_HPC2_and_U14 ( .A(Fresh[396]), .B(cell_2110_and_in[0]), 
        .Z(cell_2110_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2110_a_HPC2_and_U13 ( .A(Fresh[396]), .B(cell_2110_and_in[1]), 
        .Z(cell_2110_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2110_a_HPC2_and_U12 ( .A1(cell_2110_a_HPC2_and_a_reg[1]), .A2(
        cell_2110_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2110_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2110_a_HPC2_and_U11 ( .A1(cell_2110_a_HPC2_and_a_reg[0]), .A2(
        cell_2110_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2110_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2110_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2110_a_HPC2_and_n9), .ZN(cell_2110_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2110_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2110_a_HPC2_and_n9), .ZN(cell_2110_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2110_a_HPC2_and_U8 ( .A(Fresh[396]), .ZN(cell_2110_a_HPC2_and_n9) );
  AND2_X1 cell_2110_a_HPC2_and_U7 ( .A1(cell_2110_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2110_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2110_a_HPC2_and_U6 ( .A1(cell_2110_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2110_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2110_a_HPC2_and_U5 ( .A(cell_2110_a_HPC2_and_n8), .B(
        cell_2110_a_HPC2_and_z_1__1_), .ZN(cell_2110_and_out[1]) );
  XNOR2_X1 cell_2110_a_HPC2_and_U4 ( .A(
        cell_2110_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2110_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2110_a_HPC2_and_n8) );
  XNOR2_X1 cell_2110_a_HPC2_and_U3 ( .A(cell_2110_a_HPC2_and_n7), .B(
        cell_2110_a_HPC2_and_z_0__0_), .ZN(cell_2110_and_out[0]) );
  XNOR2_X1 cell_2110_a_HPC2_and_U2 ( .A(
        cell_2110_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2110_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2110_a_HPC2_and_n7) );
  DFF_X1 cell_2110_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2110_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2110_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2110_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2110_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2110_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2110_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2110_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2110_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2110_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2111_U4 ( .A(signal_4105), .B(cell_2111_and_out[1]), .Z(
        signal_4137) );
  XOR2_X1 cell_2111_U3 ( .A(signal_2355), .B(cell_2111_and_out[0]), .Z(
        signal_2379) );
  XOR2_X1 cell_2111_U2 ( .A(signal_4105), .B(signal_4107), .Z(
        cell_2111_and_in[1]) );
  XOR2_X1 cell_2111_U1 ( .A(signal_2355), .B(signal_2357), .Z(
        cell_2111_and_in[0]) );
  XOR2_X1 cell_2111_a_HPC2_and_U14 ( .A(Fresh[397]), .B(cell_2111_and_in[0]), 
        .Z(cell_2111_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2111_a_HPC2_and_U13 ( .A(Fresh[397]), .B(cell_2111_and_in[1]), 
        .Z(cell_2111_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2111_a_HPC2_and_U12 ( .A1(cell_2111_a_HPC2_and_a_reg[1]), .A2(
        cell_2111_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2111_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2111_a_HPC2_and_U11 ( .A1(cell_2111_a_HPC2_and_a_reg[0]), .A2(
        cell_2111_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2111_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2111_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2111_a_HPC2_and_n9), 
        .ZN(cell_2111_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2111_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2111_a_HPC2_and_n9), 
        .ZN(cell_2111_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2111_a_HPC2_and_U8 ( .A(Fresh[397]), .ZN(cell_2111_a_HPC2_and_n9) );
  AND2_X1 cell_2111_a_HPC2_and_U7 ( .A1(cell_2111_and_in[1]), .A2(n391), .ZN(
        cell_2111_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2111_a_HPC2_and_U6 ( .A1(cell_2111_and_in[0]), .A2(n390), .ZN(
        cell_2111_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2111_a_HPC2_and_U5 ( .A(cell_2111_a_HPC2_and_n8), .B(
        cell_2111_a_HPC2_and_z_1__1_), .ZN(cell_2111_and_out[1]) );
  XNOR2_X1 cell_2111_a_HPC2_and_U4 ( .A(
        cell_2111_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2111_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2111_a_HPC2_and_n8) );
  XNOR2_X1 cell_2111_a_HPC2_and_U3 ( .A(cell_2111_a_HPC2_and_n7), .B(
        cell_2111_a_HPC2_and_z_0__0_), .ZN(cell_2111_and_out[0]) );
  XNOR2_X1 cell_2111_a_HPC2_and_U2 ( .A(
        cell_2111_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2111_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2111_a_HPC2_and_n7) );
  DFF_X1 cell_2111_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2111_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2111_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2111_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2111_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2111_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2111_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2111_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2111_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2111_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2112_U4 ( .A(signal_4101), .B(cell_2112_and_out[1]), .Z(
        signal_4138) );
  XOR2_X1 cell_2112_U3 ( .A(signal_2351), .B(cell_2112_and_out[0]), .Z(
        signal_2380) );
  XOR2_X1 cell_2112_U2 ( .A(signal_4101), .B(signal_4104), .Z(
        cell_2112_and_in[1]) );
  XOR2_X1 cell_2112_U1 ( .A(signal_2351), .B(signal_2354), .Z(
        cell_2112_and_in[0]) );
  XOR2_X1 cell_2112_a_HPC2_and_U14 ( .A(Fresh[398]), .B(cell_2112_and_in[0]), 
        .Z(cell_2112_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2112_a_HPC2_and_U13 ( .A(Fresh[398]), .B(cell_2112_and_in[1]), 
        .Z(cell_2112_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2112_a_HPC2_and_U12 ( .A1(cell_2112_a_HPC2_and_a_reg[1]), .A2(
        cell_2112_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2112_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2112_a_HPC2_and_U11 ( .A1(cell_2112_a_HPC2_and_a_reg[0]), .A2(
        cell_2112_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2112_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2112_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2112_a_HPC2_and_n9), 
        .ZN(cell_2112_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2112_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2112_a_HPC2_and_n9), 
        .ZN(cell_2112_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2112_a_HPC2_and_U8 ( .A(Fresh[398]), .ZN(cell_2112_a_HPC2_and_n9) );
  AND2_X1 cell_2112_a_HPC2_and_U7 ( .A1(cell_2112_and_in[1]), .A2(n391), .ZN(
        cell_2112_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2112_a_HPC2_and_U6 ( .A1(cell_2112_and_in[0]), .A2(n390), .ZN(
        cell_2112_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2112_a_HPC2_and_U5 ( .A(cell_2112_a_HPC2_and_n8), .B(
        cell_2112_a_HPC2_and_z_1__1_), .ZN(cell_2112_and_out[1]) );
  XNOR2_X1 cell_2112_a_HPC2_and_U4 ( .A(
        cell_2112_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2112_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2112_a_HPC2_and_n8) );
  XNOR2_X1 cell_2112_a_HPC2_and_U3 ( .A(cell_2112_a_HPC2_and_n7), .B(
        cell_2112_a_HPC2_and_z_0__0_), .ZN(cell_2112_and_out[0]) );
  XNOR2_X1 cell_2112_a_HPC2_and_U2 ( .A(
        cell_2112_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2112_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2112_a_HPC2_and_n7) );
  DFF_X1 cell_2112_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2112_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2112_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2112_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2112_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2112_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2112_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2112_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2112_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2112_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2113_U4 ( .A(signal_4113), .B(cell_2113_and_out[1]), .Z(
        signal_4139) );
  XOR2_X1 cell_2113_U3 ( .A(signal_2363), .B(cell_2113_and_out[0]), .Z(
        signal_2381) );
  XOR2_X1 cell_2113_U2 ( .A(signal_4113), .B(signal_4115), .Z(
        cell_2113_and_in[1]) );
  XOR2_X1 cell_2113_U1 ( .A(signal_2363), .B(signal_2365), .Z(
        cell_2113_and_in[0]) );
  XOR2_X1 cell_2113_a_HPC2_and_U14 ( .A(Fresh[399]), .B(cell_2113_and_in[0]), 
        .Z(cell_2113_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2113_a_HPC2_and_U13 ( .A(Fresh[399]), .B(cell_2113_and_in[1]), 
        .Z(cell_2113_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2113_a_HPC2_and_U12 ( .A1(cell_2113_a_HPC2_and_a_reg[1]), .A2(
        cell_2113_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2113_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2113_a_HPC2_and_U11 ( .A1(cell_2113_a_HPC2_and_a_reg[0]), .A2(
        cell_2113_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2113_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2113_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2113_a_HPC2_and_n9), 
        .ZN(cell_2113_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2113_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2113_a_HPC2_and_n9), 
        .ZN(cell_2113_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2113_a_HPC2_and_U8 ( .A(Fresh[399]), .ZN(cell_2113_a_HPC2_and_n9) );
  AND2_X1 cell_2113_a_HPC2_and_U7 ( .A1(cell_2113_and_in[1]), .A2(n391), .ZN(
        cell_2113_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2113_a_HPC2_and_U6 ( .A1(cell_2113_and_in[0]), .A2(n390), .ZN(
        cell_2113_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2113_a_HPC2_and_U5 ( .A(cell_2113_a_HPC2_and_n8), .B(
        cell_2113_a_HPC2_and_z_1__1_), .ZN(cell_2113_and_out[1]) );
  XNOR2_X1 cell_2113_a_HPC2_and_U4 ( .A(
        cell_2113_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2113_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2113_a_HPC2_and_n8) );
  XNOR2_X1 cell_2113_a_HPC2_and_U3 ( .A(cell_2113_a_HPC2_and_n7), .B(
        cell_2113_a_HPC2_and_z_0__0_), .ZN(cell_2113_and_out[0]) );
  XNOR2_X1 cell_2113_a_HPC2_and_U2 ( .A(
        cell_2113_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2113_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2113_a_HPC2_and_n7) );
  DFF_X1 cell_2113_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2113_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2113_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2113_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2113_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2113_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2113_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2113_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2113_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2113_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2114_U4 ( .A(signal_4103), .B(cell_2114_and_out[1]), .Z(
        signal_4140) );
  XOR2_X1 cell_2114_U3 ( .A(signal_2353), .B(cell_2114_and_out[0]), .Z(
        signal_2382) );
  XOR2_X1 cell_2114_U2 ( .A(signal_4103), .B(signal_4106), .Z(
        cell_2114_and_in[1]) );
  XOR2_X1 cell_2114_U1 ( .A(signal_2353), .B(signal_2356), .Z(
        cell_2114_and_in[0]) );
  XOR2_X1 cell_2114_a_HPC2_and_U14 ( .A(Fresh[400]), .B(cell_2114_and_in[0]), 
        .Z(cell_2114_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2114_a_HPC2_and_U13 ( .A(Fresh[400]), .B(cell_2114_and_in[1]), 
        .Z(cell_2114_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2114_a_HPC2_and_U12 ( .A1(cell_2114_a_HPC2_and_a_reg[1]), .A2(
        cell_2114_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2114_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2114_a_HPC2_and_U11 ( .A1(cell_2114_a_HPC2_and_a_reg[0]), .A2(
        cell_2114_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2114_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2114_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2114_a_HPC2_and_n9), 
        .ZN(cell_2114_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2114_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2114_a_HPC2_and_n9), 
        .ZN(cell_2114_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2114_a_HPC2_and_U8 ( .A(Fresh[400]), .ZN(cell_2114_a_HPC2_and_n9) );
  AND2_X1 cell_2114_a_HPC2_and_U7 ( .A1(cell_2114_and_in[1]), .A2(n391), .ZN(
        cell_2114_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2114_a_HPC2_and_U6 ( .A1(cell_2114_and_in[0]), .A2(n390), .ZN(
        cell_2114_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2114_a_HPC2_and_U5 ( .A(cell_2114_a_HPC2_and_n8), .B(
        cell_2114_a_HPC2_and_z_1__1_), .ZN(cell_2114_and_out[1]) );
  XNOR2_X1 cell_2114_a_HPC2_and_U4 ( .A(
        cell_2114_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2114_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2114_a_HPC2_and_n8) );
  XNOR2_X1 cell_2114_a_HPC2_and_U3 ( .A(cell_2114_a_HPC2_and_n7), .B(
        cell_2114_a_HPC2_and_z_0__0_), .ZN(cell_2114_and_out[0]) );
  XNOR2_X1 cell_2114_a_HPC2_and_U2 ( .A(
        cell_2114_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2114_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2114_a_HPC2_and_n7) );
  DFF_X1 cell_2114_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2114_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2114_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2114_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2114_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2114_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2114_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2114_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2114_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2114_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2115_U4 ( .A(signal_4097), .B(cell_2115_and_out[1]), .Z(
        signal_4141) );
  XOR2_X1 cell_2115_U3 ( .A(signal_2347), .B(cell_2115_and_out[0]), .Z(
        signal_2383) );
  XOR2_X1 cell_2115_U2 ( .A(signal_4097), .B(signal_4116), .Z(
        cell_2115_and_in[1]) );
  XOR2_X1 cell_2115_U1 ( .A(signal_2347), .B(signal_2366), .Z(
        cell_2115_and_in[0]) );
  XOR2_X1 cell_2115_a_HPC2_and_U14 ( .A(Fresh[401]), .B(cell_2115_and_in[0]), 
        .Z(cell_2115_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2115_a_HPC2_and_U13 ( .A(Fresh[401]), .B(cell_2115_and_in[1]), 
        .Z(cell_2115_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2115_a_HPC2_and_U12 ( .A1(cell_2115_a_HPC2_and_a_reg[1]), .A2(
        cell_2115_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2115_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2115_a_HPC2_and_U11 ( .A1(cell_2115_a_HPC2_and_a_reg[0]), .A2(
        cell_2115_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2115_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2115_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2115_a_HPC2_and_n9), 
        .ZN(cell_2115_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2115_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2115_a_HPC2_and_n9), 
        .ZN(cell_2115_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2115_a_HPC2_and_U8 ( .A(Fresh[401]), .ZN(cell_2115_a_HPC2_and_n9) );
  AND2_X1 cell_2115_a_HPC2_and_U7 ( .A1(cell_2115_and_in[1]), .A2(n391), .ZN(
        cell_2115_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2115_a_HPC2_and_U6 ( .A1(cell_2115_and_in[0]), .A2(n390), .ZN(
        cell_2115_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2115_a_HPC2_and_U5 ( .A(cell_2115_a_HPC2_and_n8), .B(
        cell_2115_a_HPC2_and_z_1__1_), .ZN(cell_2115_and_out[1]) );
  XNOR2_X1 cell_2115_a_HPC2_and_U4 ( .A(
        cell_2115_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2115_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2115_a_HPC2_and_n8) );
  XNOR2_X1 cell_2115_a_HPC2_and_U3 ( .A(cell_2115_a_HPC2_and_n7), .B(
        cell_2115_a_HPC2_and_z_0__0_), .ZN(cell_2115_and_out[0]) );
  XNOR2_X1 cell_2115_a_HPC2_and_U2 ( .A(
        cell_2115_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2115_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2115_a_HPC2_and_n7) );
  DFF_X1 cell_2115_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2115_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2115_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2115_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2115_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2115_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2115_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2115_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2115_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2115_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2116_U4 ( .A(signal_4095), .B(cell_2116_and_out[1]), .Z(
        signal_4142) );
  XOR2_X1 cell_2116_U3 ( .A(signal_2345), .B(cell_2116_and_out[0]), .Z(
        signal_2384) );
  XOR2_X1 cell_2116_U2 ( .A(signal_4095), .B(signal_4090), .Z(
        cell_2116_and_in[1]) );
  XOR2_X1 cell_2116_U1 ( .A(signal_2345), .B(signal_2340), .Z(
        cell_2116_and_in[0]) );
  XOR2_X1 cell_2116_a_HPC2_and_U14 ( .A(Fresh[402]), .B(cell_2116_and_in[0]), 
        .Z(cell_2116_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2116_a_HPC2_and_U13 ( .A(Fresh[402]), .B(cell_2116_and_in[1]), 
        .Z(cell_2116_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2116_a_HPC2_and_U12 ( .A1(cell_2116_a_HPC2_and_a_reg[1]), .A2(
        cell_2116_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2116_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2116_a_HPC2_and_U11 ( .A1(cell_2116_a_HPC2_and_a_reg[0]), .A2(
        cell_2116_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2116_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2116_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2116_a_HPC2_and_n9), 
        .ZN(cell_2116_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2116_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2116_a_HPC2_and_n9), 
        .ZN(cell_2116_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2116_a_HPC2_and_U8 ( .A(Fresh[402]), .ZN(cell_2116_a_HPC2_and_n9) );
  AND2_X1 cell_2116_a_HPC2_and_U7 ( .A1(cell_2116_and_in[1]), .A2(n391), .ZN(
        cell_2116_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2116_a_HPC2_and_U6 ( .A1(cell_2116_and_in[0]), .A2(n390), .ZN(
        cell_2116_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2116_a_HPC2_and_U5 ( .A(cell_2116_a_HPC2_and_n8), .B(
        cell_2116_a_HPC2_and_z_1__1_), .ZN(cell_2116_and_out[1]) );
  XNOR2_X1 cell_2116_a_HPC2_and_U4 ( .A(
        cell_2116_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2116_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2116_a_HPC2_and_n8) );
  XNOR2_X1 cell_2116_a_HPC2_and_U3 ( .A(cell_2116_a_HPC2_and_n7), .B(
        cell_2116_a_HPC2_and_z_0__0_), .ZN(cell_2116_and_out[0]) );
  XNOR2_X1 cell_2116_a_HPC2_and_U2 ( .A(
        cell_2116_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2116_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2116_a_HPC2_and_n7) );
  DFF_X1 cell_2116_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2116_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2116_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2116_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2116_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2116_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2116_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2116_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2116_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2116_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2117_U4 ( .A(signal_4112), .B(cell_2117_and_out[1]), .Z(
        signal_4143) );
  XOR2_X1 cell_2117_U3 ( .A(signal_2362), .B(cell_2117_and_out[0]), .Z(
        signal_2385) );
  XOR2_X1 cell_2117_U2 ( .A(signal_4112), .B(signal_4120), .Z(
        cell_2117_and_in[1]) );
  XOR2_X1 cell_2117_U1 ( .A(signal_2362), .B(signal_2370), .Z(
        cell_2117_and_in[0]) );
  XOR2_X1 cell_2117_a_HPC2_and_U14 ( .A(Fresh[403]), .B(cell_2117_and_in[0]), 
        .Z(cell_2117_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2117_a_HPC2_and_U13 ( .A(Fresh[403]), .B(cell_2117_and_in[1]), 
        .Z(cell_2117_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2117_a_HPC2_and_U12 ( .A1(cell_2117_a_HPC2_and_a_reg[1]), .A2(
        cell_2117_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2117_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2117_a_HPC2_and_U11 ( .A1(cell_2117_a_HPC2_and_a_reg[0]), .A2(
        cell_2117_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2117_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2117_a_HPC2_and_U10 ( .A1(n391), .A2(cell_2117_a_HPC2_and_n9), 
        .ZN(cell_2117_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2117_a_HPC2_and_U9 ( .A1(n390), .A2(cell_2117_a_HPC2_and_n9), 
        .ZN(cell_2117_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2117_a_HPC2_and_U8 ( .A(Fresh[403]), .ZN(cell_2117_a_HPC2_and_n9) );
  AND2_X1 cell_2117_a_HPC2_and_U7 ( .A1(cell_2117_and_in[1]), .A2(n391), .ZN(
        cell_2117_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2117_a_HPC2_and_U6 ( .A1(cell_2117_and_in[0]), .A2(n390), .ZN(
        cell_2117_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2117_a_HPC2_and_U5 ( .A(cell_2117_a_HPC2_and_n8), .B(
        cell_2117_a_HPC2_and_z_1__1_), .ZN(cell_2117_and_out[1]) );
  XNOR2_X1 cell_2117_a_HPC2_and_U4 ( .A(
        cell_2117_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2117_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2117_a_HPC2_and_n8) );
  XNOR2_X1 cell_2117_a_HPC2_and_U3 ( .A(cell_2117_a_HPC2_and_n7), .B(
        cell_2117_a_HPC2_and_z_0__0_), .ZN(cell_2117_and_out[0]) );
  XNOR2_X1 cell_2117_a_HPC2_and_U2 ( .A(
        cell_2117_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2117_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2117_a_HPC2_and_n7) );
  DFF_X1 cell_2117_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2117_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2117_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_a_i_0_s_current_state_reg ( .D(n390), .CK(clk), 
        .Q(cell_2117_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2117_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2117_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_a_i_1_s_current_state_reg ( .D(n391), .CK(clk), 
        .Q(cell_2117_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2117_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2117_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2117_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2118_U4 ( .A(signal_4117), .B(cell_2118_and_out[1]), .Z(
        signal_4144) );
  XOR2_X1 cell_2118_U3 ( .A(signal_2367), .B(cell_2118_and_out[0]), .Z(
        signal_2386) );
  XOR2_X1 cell_2118_U2 ( .A(signal_4117), .B(signal_4110), .Z(
        cell_2118_and_in[1]) );
  XOR2_X1 cell_2118_U1 ( .A(signal_2367), .B(signal_2360), .Z(
        cell_2118_and_in[0]) );
  XOR2_X1 cell_2118_a_HPC2_and_U14 ( .A(Fresh[404]), .B(cell_2118_and_in[0]), 
        .Z(cell_2118_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2118_a_HPC2_and_U13 ( .A(Fresh[404]), .B(cell_2118_and_in[1]), 
        .Z(cell_2118_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2118_a_HPC2_and_U12 ( .A1(cell_2118_a_HPC2_and_a_reg[1]), .A2(
        cell_2118_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2118_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2118_a_HPC2_and_U11 ( .A1(cell_2118_a_HPC2_and_a_reg[0]), .A2(
        cell_2118_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2118_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2118_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2118_a_HPC2_and_n9), .ZN(cell_2118_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2118_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2118_a_HPC2_and_n9), .ZN(cell_2118_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2118_a_HPC2_and_U8 ( .A(Fresh[404]), .ZN(cell_2118_a_HPC2_and_n9) );
  AND2_X1 cell_2118_a_HPC2_and_U7 ( .A1(cell_2118_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2118_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2118_a_HPC2_and_U6 ( .A1(cell_2118_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2118_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2118_a_HPC2_and_U5 ( .A(cell_2118_a_HPC2_and_n8), .B(
        cell_2118_a_HPC2_and_z_1__1_), .ZN(cell_2118_and_out[1]) );
  XNOR2_X1 cell_2118_a_HPC2_and_U4 ( .A(
        cell_2118_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2118_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2118_a_HPC2_and_n8) );
  XNOR2_X1 cell_2118_a_HPC2_and_U3 ( .A(cell_2118_a_HPC2_and_n7), .B(
        cell_2118_a_HPC2_and_z_0__0_), .ZN(cell_2118_and_out[0]) );
  XNOR2_X1 cell_2118_a_HPC2_and_U2 ( .A(
        cell_2118_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2118_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2118_a_HPC2_and_n7) );
  DFF_X1 cell_2118_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2118_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2118_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2118_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2118_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2118_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2118_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2118_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2118_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2118_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2119_U4 ( .A(signal_4096), .B(cell_2119_and_out[1]), .Z(
        signal_4145) );
  XOR2_X1 cell_2119_U3 ( .A(signal_2346), .B(cell_2119_and_out[0]), .Z(
        signal_2387) );
  XOR2_X1 cell_2119_U2 ( .A(signal_4096), .B(signal_4093), .Z(
        cell_2119_and_in[1]) );
  XOR2_X1 cell_2119_U1 ( .A(signal_2346), .B(signal_2343), .Z(
        cell_2119_and_in[0]) );
  XOR2_X1 cell_2119_a_HPC2_and_U14 ( .A(Fresh[405]), .B(cell_2119_and_in[0]), 
        .Z(cell_2119_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2119_a_HPC2_and_U13 ( .A(Fresh[405]), .B(cell_2119_and_in[1]), 
        .Z(cell_2119_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2119_a_HPC2_and_U12 ( .A1(cell_2119_a_HPC2_and_a_reg[1]), .A2(
        cell_2119_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2119_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2119_a_HPC2_and_U11 ( .A1(cell_2119_a_HPC2_and_a_reg[0]), .A2(
        cell_2119_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2119_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2119_a_HPC2_and_U10 ( .A1(signal_3239), .A2(
        cell_2119_a_HPC2_and_n9), .ZN(cell_2119_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2119_a_HPC2_and_U9 ( .A1(signal_1510), .A2(
        cell_2119_a_HPC2_and_n9), .ZN(cell_2119_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2119_a_HPC2_and_U8 ( .A(Fresh[405]), .ZN(cell_2119_a_HPC2_and_n9) );
  AND2_X1 cell_2119_a_HPC2_and_U7 ( .A1(cell_2119_and_in[1]), .A2(signal_3239), 
        .ZN(cell_2119_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2119_a_HPC2_and_U6 ( .A1(cell_2119_and_in[0]), .A2(signal_1510), 
        .ZN(cell_2119_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2119_a_HPC2_and_U5 ( .A(cell_2119_a_HPC2_and_n8), .B(
        cell_2119_a_HPC2_and_z_1__1_), .ZN(cell_2119_and_out[1]) );
  XNOR2_X1 cell_2119_a_HPC2_and_U4 ( .A(
        cell_2119_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2119_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2119_a_HPC2_and_n8) );
  XNOR2_X1 cell_2119_a_HPC2_and_U3 ( .A(cell_2119_a_HPC2_and_n7), .B(
        cell_2119_a_HPC2_and_z_0__0_), .ZN(cell_2119_and_out[0]) );
  XNOR2_X1 cell_2119_a_HPC2_and_U2 ( .A(
        cell_2119_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2119_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2119_a_HPC2_and_n7) );
  DFF_X1 cell_2119_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2119_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2119_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1510), 
        .CK(clk), .Q(cell_2119_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2119_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2119_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3239), 
        .CK(clk), .Q(cell_2119_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2119_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2119_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2119_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  MUX2_X1 cell_56_Ins_0_U1 ( .A(signal_1405), .B(signal_1413), .S(n473), .Z(
        signal_1421) );
  MUX2_X1 cell_56_Ins_1_U1 ( .A(signal_4146), .B(signal_2390), .S(n473), .Z(
        signal_4154) );
  MUX2_X1 cell_57_Ins_0_U1 ( .A(signal_1404), .B(signal_1412), .S(n473), .Z(
        signal_1420) );
  MUX2_X1 cell_57_Ins_1_U1 ( .A(signal_4151), .B(signal_2393), .S(n473), .Z(
        signal_4155) );
  MUX2_X1 cell_58_Ins_0_U1 ( .A(signal_1403), .B(signal_1411), .S(n473), .Z(
        signal_1419) );
  MUX2_X1 cell_58_Ins_1_U1 ( .A(signal_4148), .B(signal_2396), .S(n473), .Z(
        signal_4156) );
  MUX2_X1 cell_59_Ins_0_U1 ( .A(signal_1402), .B(signal_1410), .S(signal_399), 
        .Z(signal_1418) );
  MUX2_X1 cell_59_Ins_1_U1 ( .A(signal_4150), .B(signal_2399), .S(signal_399), 
        .Z(signal_4157) );
  MUX2_X1 cell_60_Ins_0_U1 ( .A(signal_1401), .B(signal_1409), .S(signal_399), 
        .Z(signal_1417) );
  MUX2_X1 cell_60_Ins_1_U1 ( .A(signal_4152), .B(signal_2402), .S(signal_399), 
        .Z(signal_4158) );
  MUX2_X1 cell_61_Ins_0_U1 ( .A(signal_1400), .B(signal_1408), .S(signal_399), 
        .Z(signal_1416) );
  MUX2_X1 cell_61_Ins_1_U1 ( .A(signal_4153), .B(signal_2405), .S(signal_399), 
        .Z(signal_4159) );
  MUX2_X1 cell_62_Ins_0_U1 ( .A(signal_1399), .B(signal_1407), .S(signal_399), 
        .Z(signal_1415) );
  MUX2_X1 cell_62_Ins_1_U1 ( .A(signal_4147), .B(signal_2408), .S(signal_399), 
        .Z(signal_4160) );
  MUX2_X1 cell_63_Ins_0_U1 ( .A(signal_1398), .B(signal_1406), .S(signal_399), 
        .Z(signal_1414) );
  MUX2_X1 cell_63_Ins_1_U1 ( .A(signal_4149), .B(signal_2411), .S(signal_399), 
        .Z(signal_4161) );
  MUX2_X1 cell_445_Ins_0_U1 ( .A(signal_1557), .B(ciphertext_s0[8]), .S(n349), 
        .Z(signal_705) );
  MUX2_X1 cell_445_Ins_1_U1 ( .A(signal_4187), .B(ciphertext_s1[8]), .S(n349), 
        .Z(signal_4210) );
  MUX2_X1 cell_448_Ins_0_U1 ( .A(signal_1556), .B(ciphertext_s0[9]), .S(n338), 
        .Z(signal_707) );
  MUX2_X1 cell_448_Ins_1_U1 ( .A(signal_4189), .B(ciphertext_s1[9]), .S(n338), 
        .Z(signal_4211) );
  MUX2_X1 cell_451_Ins_0_U1 ( .A(signal_1555), .B(ciphertext_s0[10]), .S(n345), 
        .Z(signal_709) );
  MUX2_X1 cell_451_Ins_1_U1 ( .A(signal_4191), .B(ciphertext_s1[10]), .S(n345), 
        .Z(signal_4212) );
  MUX2_X1 cell_454_Ins_0_U1 ( .A(signal_1554), .B(ciphertext_s0[11]), .S(n339), 
        .Z(signal_711) );
  MUX2_X1 cell_454_Ins_1_U1 ( .A(signal_4193), .B(ciphertext_s1[11]), .S(n339), 
        .Z(signal_4213) );
  MUX2_X1 cell_457_Ins_0_U1 ( .A(signal_1553), .B(ciphertext_s0[12]), .S(n339), 
        .Z(signal_713) );
  MUX2_X1 cell_457_Ins_1_U1 ( .A(signal_4195), .B(ciphertext_s1[12]), .S(n339), 
        .Z(signal_4214) );
  MUX2_X1 cell_460_Ins_0_U1 ( .A(signal_1552), .B(ciphertext_s0[13]), .S(n339), 
        .Z(signal_715) );
  MUX2_X1 cell_460_Ins_1_U1 ( .A(signal_4197), .B(ciphertext_s1[13]), .S(n339), 
        .Z(signal_4215) );
  MUX2_X1 cell_463_Ins_0_U1 ( .A(signal_1551), .B(ciphertext_s0[14]), .S(n338), 
        .Z(signal_717) );
  MUX2_X1 cell_463_Ins_1_U1 ( .A(signal_4199), .B(ciphertext_s1[14]), .S(n338), 
        .Z(signal_4216) );
  MUX2_X1 cell_466_Ins_0_U1 ( .A(signal_1550), .B(ciphertext_s0[15]), .S(n338), 
        .Z(signal_719) );
  MUX2_X1 cell_466_Ins_1_U1 ( .A(signal_4201), .B(ciphertext_s1[15]), .S(n338), 
        .Z(signal_4217) );
  MUX2_X1 cell_613_Ins_0_U1 ( .A(signal_1421), .B(signal_1453), .S(n323), .Z(
        signal_1525) );
  MUX2_X1 cell_613_Ins_1_U1 ( .A(signal_4154), .B(signal_3262), .S(n323), .Z(
        signal_4170) );
  MUX2_X1 cell_614_Ins_0_U1 ( .A(signal_1420), .B(signal_1452), .S(n311), .Z(
        signal_1524) );
  MUX2_X1 cell_614_Ins_1_U1 ( .A(signal_4155), .B(signal_3263), .S(n311), .Z(
        signal_4171) );
  MUX2_X1 cell_615_Ins_0_U1 ( .A(signal_1419), .B(signal_1451), .S(n309), .Z(
        signal_1523) );
  MUX2_X1 cell_615_Ins_1_U1 ( .A(signal_4156), .B(signal_3240), .S(n309), .Z(
        signal_4172) );
  MUX2_X1 cell_616_Ins_0_U1 ( .A(signal_1418), .B(signal_1450), .S(n315), .Z(
        signal_1522) );
  MUX2_X1 cell_616_Ins_1_U1 ( .A(signal_4157), .B(signal_3264), .S(n315), .Z(
        signal_4173) );
  MUX2_X1 cell_617_Ins_0_U1 ( .A(signal_1417), .B(signal_1449), .S(n321), .Z(
        signal_1521) );
  MUX2_X1 cell_617_Ins_1_U1 ( .A(signal_4158), .B(signal_3265), .S(n321), .Z(
        signal_4174) );
  MUX2_X1 cell_618_Ins_0_U1 ( .A(signal_1416), .B(signal_1448), .S(n310), .Z(
        signal_1520) );
  MUX2_X1 cell_618_Ins_1_U1 ( .A(signal_4159), .B(signal_3241), .S(n310), .Z(
        signal_4175) );
  MUX2_X1 cell_619_Ins_0_U1 ( .A(signal_1415), .B(signal_1447), .S(n315), .Z(
        signal_1519) );
  MUX2_X1 cell_619_Ins_1_U1 ( .A(signal_4160), .B(signal_3242), .S(n315), .Z(
        signal_4176) );
  MUX2_X1 cell_620_Ins_0_U1 ( .A(signal_1414), .B(signal_1446), .S(n321), .Z(
        signal_1518) );
  MUX2_X1 cell_620_Ins_1_U1 ( .A(signal_4161), .B(signal_3243), .S(n321), .Z(
        signal_4177) );
  MUX2_X1 cell_621_Ins_0_U1 ( .A(plaintext_s0[0]), .B(signal_1525), .S(n302), 
        .Z(signal_1557) );
  MUX2_X1 cell_621_Ins_1_U1 ( .A(plaintext_s1[0]), .B(signal_4170), .S(n302), 
        .Z(signal_4187) );
  MUX2_X1 cell_622_Ins_0_U1 ( .A(plaintext_s0[1]), .B(signal_1524), .S(n306), 
        .Z(signal_1556) );
  MUX2_X1 cell_622_Ins_1_U1 ( .A(plaintext_s1[1]), .B(signal_4171), .S(n306), 
        .Z(signal_4189) );
  MUX2_X1 cell_623_Ins_0_U1 ( .A(plaintext_s0[2]), .B(signal_1523), .S(n306), 
        .Z(signal_1555) );
  MUX2_X1 cell_623_Ins_1_U1 ( .A(plaintext_s1[2]), .B(signal_4172), .S(n306), 
        .Z(signal_4191) );
  MUX2_X1 cell_624_Ins_0_U1 ( .A(plaintext_s0[3]), .B(signal_1522), .S(n295), 
        .Z(signal_1554) );
  MUX2_X1 cell_624_Ins_1_U1 ( .A(plaintext_s1[3]), .B(signal_4173), .S(n295), 
        .Z(signal_4193) );
  MUX2_X1 cell_625_Ins_0_U1 ( .A(plaintext_s0[4]), .B(signal_1521), .S(n297), 
        .Z(signal_1553) );
  MUX2_X1 cell_625_Ins_1_U1 ( .A(plaintext_s1[4]), .B(signal_4174), .S(n297), 
        .Z(signal_4195) );
  MUX2_X1 cell_626_Ins_0_U1 ( .A(plaintext_s0[5]), .B(signal_1520), .S(n296), 
        .Z(signal_1552) );
  MUX2_X1 cell_626_Ins_1_U1 ( .A(plaintext_s1[5]), .B(signal_4175), .S(n296), 
        .Z(signal_4197) );
  MUX2_X1 cell_627_Ins_0_U1 ( .A(plaintext_s0[6]), .B(signal_1519), .S(n300), 
        .Z(signal_1551) );
  MUX2_X1 cell_627_Ins_1_U1 ( .A(plaintext_s1[6]), .B(signal_4176), .S(n300), 
        .Z(signal_4199) );
  MUX2_X1 cell_628_Ins_0_U1 ( .A(plaintext_s0[7]), .B(signal_1518), .S(n289), 
        .Z(signal_1550) );
  MUX2_X1 cell_628_Ins_1_U1 ( .A(plaintext_s1[7]), .B(signal_4177), .S(n289), 
        .Z(signal_4201) );
  XNOR2_X1 cell_672_Ins0_U1 ( .A(signal_724), .B(signal_1486), .ZN(signal_1750) );
  XOR2_X1 cell_672_Ins_1_U1 ( .A(signal_4162), .B(signal_2410), .Z(signal_4178) );
  XNOR2_X1 cell_673_Ins0_U1 ( .A(signal_1494), .B(signal_1398), .ZN(signal_724) );
  XOR2_X1 cell_673_Ins_1_U1 ( .A(1'b0), .B(signal_4149), .Z(signal_4162) );
  XNOR2_X1 cell_674_Ins0_U1 ( .A(signal_725), .B(signal_1487), .ZN(signal_1751) );
  XOR2_X1 cell_674_Ins_1_U1 ( .A(signal_4163), .B(signal_2407), .Z(signal_4179) );
  XNOR2_X1 cell_675_Ins0_U1 ( .A(signal_1495), .B(signal_1399), .ZN(signal_725) );
  XOR2_X1 cell_675_Ins_1_U1 ( .A(1'b0), .B(signal_4147), .Z(signal_4163) );
  XNOR2_X1 cell_676_Ins0_U1 ( .A(signal_726), .B(signal_1488), .ZN(signal_1752) );
  XOR2_X1 cell_676_Ins_1_U1 ( .A(signal_4164), .B(signal_2404), .Z(signal_4180) );
  XNOR2_X1 cell_677_Ins0_U1 ( .A(signal_1496), .B(signal_1400), .ZN(signal_726) );
  XOR2_X1 cell_677_Ins_1_U1 ( .A(1'b0), .B(signal_4153), .Z(signal_4164) );
  XNOR2_X1 cell_678_Ins0_U1 ( .A(signal_727), .B(signal_1489), .ZN(signal_1753) );
  XOR2_X1 cell_678_Ins_1_U1 ( .A(signal_4165), .B(signal_2401), .Z(signal_4181) );
  XNOR2_X1 cell_679_Ins0_U1 ( .A(signal_1497), .B(signal_1401), .ZN(signal_727) );
  XOR2_X1 cell_679_Ins_1_U1 ( .A(1'b0), .B(signal_4152), .Z(signal_4165) );
  XNOR2_X1 cell_680_Ins0_U1 ( .A(signal_728), .B(signal_1490), .ZN(signal_1754) );
  XOR2_X1 cell_680_Ins_1_U1 ( .A(signal_4166), .B(signal_2398), .Z(signal_4182) );
  XNOR2_X1 cell_681_Ins0_U1 ( .A(signal_1498), .B(signal_1402), .ZN(signal_728) );
  XOR2_X1 cell_681_Ins_1_U1 ( .A(1'b0), .B(signal_4150), .Z(signal_4166) );
  XNOR2_X1 cell_682_Ins0_U1 ( .A(signal_729), .B(signal_1491), .ZN(signal_1755) );
  XOR2_X1 cell_682_Ins_1_U1 ( .A(signal_4167), .B(signal_2395), .Z(signal_4183) );
  XNOR2_X1 cell_683_Ins0_U1 ( .A(signal_1499), .B(signal_1403), .ZN(signal_729) );
  XOR2_X1 cell_683_Ins_1_U1 ( .A(1'b0), .B(signal_4148), .Z(signal_4167) );
  XNOR2_X1 cell_684_Ins0_U1 ( .A(signal_730), .B(signal_1492), .ZN(signal_1756) );
  XOR2_X1 cell_684_Ins_1_U1 ( .A(signal_4168), .B(signal_2392), .Z(signal_4184) );
  XNOR2_X1 cell_685_Ins0_U1 ( .A(signal_1500), .B(signal_1404), .ZN(signal_730) );
  XOR2_X1 cell_685_Ins_1_U1 ( .A(1'b0), .B(signal_4151), .Z(signal_4168) );
  XNOR2_X1 cell_686_Ins0_U1 ( .A(signal_731), .B(signal_1493), .ZN(signal_1757) );
  XOR2_X1 cell_686_Ins_1_U1 ( .A(signal_4169), .B(signal_2389), .Z(signal_4185) );
  XNOR2_X1 cell_687_Ins0_U1 ( .A(signal_1501), .B(signal_1405), .ZN(signal_731) );
  XOR2_X1 cell_687_Ins_1_U1 ( .A(1'b0), .B(signal_4146), .Z(signal_4169) );
  MUX2_X1 cell_1098_Ins_0_U1 ( .A(signal_1749), .B(signal_1055), .S(n328), .Z(
        signal_1054) );
  MUX2_X1 cell_1098_Ins_1_U1 ( .A(signal_3089), .B(signal_4202), .S(n328), .Z(
        signal_4218) );
  MUX2_X1 cell_1099_Ins_0_U1 ( .A(signal_1765), .B(signal_1757), .S(n316), .Z(
        signal_1055) );
  MUX2_X1 cell_1099_Ins_1_U1 ( .A(signal_3114), .B(signal_4185), .S(n316), .Z(
        signal_4202) );
  MUX2_X1 cell_1102_Ins_0_U1 ( .A(signal_1748), .B(signal_1058), .S(n336), .Z(
        signal_1057) );
  MUX2_X1 cell_1102_Ins_1_U1 ( .A(signal_3092), .B(signal_4203), .S(n336), .Z(
        signal_4219) );
  MUX2_X1 cell_1103_Ins_0_U1 ( .A(signal_1764), .B(signal_1756), .S(n321), .Z(
        signal_1058) );
  MUX2_X1 cell_1103_Ins_1_U1 ( .A(signal_3117), .B(signal_4184), .S(n321), .Z(
        signal_4203) );
  MUX2_X1 cell_1106_Ins_0_U1 ( .A(signal_1747), .B(signal_1061), .S(n325), .Z(
        signal_1060) );
  MUX2_X1 cell_1106_Ins_1_U1 ( .A(signal_3095), .B(signal_4204), .S(n325), .Z(
        signal_4220) );
  MUX2_X1 cell_1107_Ins_0_U1 ( .A(signal_1763), .B(signal_1755), .S(n319), .Z(
        signal_1061) );
  MUX2_X1 cell_1107_Ins_1_U1 ( .A(signal_3120), .B(signal_4183), .S(n319), .Z(
        signal_4204) );
  MUX2_X1 cell_1110_Ins_0_U1 ( .A(signal_1746), .B(signal_1064), .S(n332), .Z(
        signal_1063) );
  MUX2_X1 cell_1110_Ins_1_U1 ( .A(signal_3098), .B(signal_4205), .S(n332), .Z(
        signal_4221) );
  MUX2_X1 cell_1111_Ins_0_U1 ( .A(signal_1762), .B(signal_1754), .S(n317), .Z(
        signal_1064) );
  MUX2_X1 cell_1111_Ins_1_U1 ( .A(signal_3123), .B(signal_4182), .S(n317), .Z(
        signal_4205) );
  MUX2_X1 cell_1114_Ins_0_U1 ( .A(signal_1745), .B(signal_1067), .S(n329), .Z(
        signal_1066) );
  MUX2_X1 cell_1114_Ins_1_U1 ( .A(signal_3101), .B(signal_4206), .S(n329), .Z(
        signal_4222) );
  MUX2_X1 cell_1115_Ins_0_U1 ( .A(signal_1761), .B(signal_1753), .S(n310), .Z(
        signal_1067) );
  MUX2_X1 cell_1115_Ins_1_U1 ( .A(signal_3126), .B(signal_4181), .S(n310), .Z(
        signal_4206) );
  MUX2_X1 cell_1118_Ins_0_U1 ( .A(signal_1744), .B(signal_1070), .S(n329), .Z(
        signal_1069) );
  MUX2_X1 cell_1118_Ins_1_U1 ( .A(signal_3104), .B(signal_4207), .S(n329), .Z(
        signal_4223) );
  MUX2_X1 cell_1119_Ins_0_U1 ( .A(signal_1760), .B(signal_1752), .S(n318), .Z(
        signal_1070) );
  MUX2_X1 cell_1119_Ins_1_U1 ( .A(signal_3129), .B(signal_4180), .S(n318), .Z(
        signal_4207) );
  MUX2_X1 cell_1122_Ins_0_U1 ( .A(signal_1743), .B(signal_1073), .S(n335), .Z(
        signal_1072) );
  MUX2_X1 cell_1122_Ins_1_U1 ( .A(signal_3107), .B(signal_4208), .S(n335), .Z(
        signal_4224) );
  MUX2_X1 cell_1123_Ins_0_U1 ( .A(signal_1759), .B(signal_1751), .S(n316), .Z(
        signal_1073) );
  MUX2_X1 cell_1123_Ins_1_U1 ( .A(signal_3132), .B(signal_4179), .S(n316), .Z(
        signal_4208) );
  MUX2_X1 cell_1126_Ins_0_U1 ( .A(signal_1742), .B(signal_1076), .S(n333), .Z(
        signal_1075) );
  MUX2_X1 cell_1126_Ins_1_U1 ( .A(signal_3110), .B(signal_4209), .S(n333), .Z(
        signal_4225) );
  MUX2_X1 cell_1127_Ins_0_U1 ( .A(signal_1758), .B(signal_1750), .S(n314), .Z(
        signal_1076) );
  MUX2_X1 cell_1127_Ins_1_U1 ( .A(signal_3135), .B(signal_4178), .S(n314), .Z(
        signal_4209) );
  XOR2_X1 cell_2120_U4 ( .A(signal_4141), .B(cell_2120_and_out[1]), .Z(
        signal_4146) );
  XOR2_X1 cell_2120_U3 ( .A(signal_2383), .B(cell_2120_and_out[0]), .Z(
        signal_1405) );
  XOR2_X1 cell_2120_U2 ( .A(signal_4141), .B(signal_4135), .Z(
        cell_2120_and_in[1]) );
  XOR2_X1 cell_2120_U1 ( .A(signal_2383), .B(signal_2377), .Z(
        cell_2120_and_in[0]) );
  XOR2_X1 cell_2120_a_HPC2_and_U14 ( .A(Fresh[406]), .B(cell_2120_and_in[0]), 
        .Z(cell_2120_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2120_a_HPC2_and_U13 ( .A(Fresh[406]), .B(cell_2120_and_in[1]), 
        .Z(cell_2120_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2120_a_HPC2_and_U12 ( .A1(cell_2120_a_HPC2_and_a_reg[1]), .A2(
        cell_2120_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2120_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2120_a_HPC2_and_U11 ( .A1(cell_2120_a_HPC2_and_a_reg[0]), .A2(
        cell_2120_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2120_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2120_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2120_a_HPC2_and_n9), .ZN(cell_2120_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2120_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2120_a_HPC2_and_n9), .ZN(cell_2120_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2120_a_HPC2_and_U8 ( .A(Fresh[406]), .ZN(cell_2120_a_HPC2_and_n9) );
  AND2_X1 cell_2120_a_HPC2_and_U7 ( .A1(cell_2120_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2120_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2120_a_HPC2_and_U6 ( .A1(cell_2120_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2120_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2120_a_HPC2_and_U5 ( .A(cell_2120_a_HPC2_and_n8), .B(
        cell_2120_a_HPC2_and_z_1__1_), .ZN(cell_2120_and_out[1]) );
  XNOR2_X1 cell_2120_a_HPC2_and_U4 ( .A(
        cell_2120_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2120_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2120_a_HPC2_and_n8) );
  XNOR2_X1 cell_2120_a_HPC2_and_U3 ( .A(cell_2120_a_HPC2_and_n7), .B(
        cell_2120_a_HPC2_and_z_0__0_), .ZN(cell_2120_and_out[0]) );
  XNOR2_X1 cell_2120_a_HPC2_and_U2 ( .A(
        cell_2120_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2120_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2120_a_HPC2_and_n7) );
  DFF_X1 cell_2120_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2120_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2120_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2120_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2120_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2120_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2120_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2120_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2120_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2120_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2121_U4 ( .A(signal_4134), .B(cell_2121_and_out[1]), .Z(
        signal_4147) );
  XOR2_X1 cell_2121_U3 ( .A(signal_2376), .B(cell_2121_and_out[0]), .Z(
        signal_1399) );
  XOR2_X1 cell_2121_U2 ( .A(signal_4134), .B(signal_4145), .Z(
        cell_2121_and_in[1]) );
  XOR2_X1 cell_2121_U1 ( .A(signal_2376), .B(signal_2387), .Z(
        cell_2121_and_in[0]) );
  XOR2_X1 cell_2121_a_HPC2_and_U14 ( .A(Fresh[407]), .B(cell_2121_and_in[0]), 
        .Z(cell_2121_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2121_a_HPC2_and_U13 ( .A(Fresh[407]), .B(cell_2121_and_in[1]), 
        .Z(cell_2121_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2121_a_HPC2_and_U12 ( .A1(cell_2121_a_HPC2_and_a_reg[1]), .A2(
        cell_2121_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2121_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2121_a_HPC2_and_U11 ( .A1(cell_2121_a_HPC2_and_a_reg[0]), .A2(
        cell_2121_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2121_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2121_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2121_a_HPC2_and_n9), .ZN(cell_2121_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2121_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2121_a_HPC2_and_n9), .ZN(cell_2121_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2121_a_HPC2_and_U8 ( .A(Fresh[407]), .ZN(cell_2121_a_HPC2_and_n9) );
  AND2_X1 cell_2121_a_HPC2_and_U7 ( .A1(cell_2121_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2121_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2121_a_HPC2_and_U6 ( .A1(cell_2121_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2121_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2121_a_HPC2_and_U5 ( .A(cell_2121_a_HPC2_and_n8), .B(
        cell_2121_a_HPC2_and_z_1__1_), .ZN(cell_2121_and_out[1]) );
  XNOR2_X1 cell_2121_a_HPC2_and_U4 ( .A(
        cell_2121_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2121_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2121_a_HPC2_and_n8) );
  XNOR2_X1 cell_2121_a_HPC2_and_U3 ( .A(cell_2121_a_HPC2_and_n7), .B(
        cell_2121_a_HPC2_and_z_0__0_), .ZN(cell_2121_and_out[0]) );
  XNOR2_X1 cell_2121_a_HPC2_and_U2 ( .A(
        cell_2121_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2121_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2121_a_HPC2_and_n7) );
  DFF_X1 cell_2121_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2121_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2121_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2121_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2121_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2121_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2121_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2121_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2121_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2121_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2122_U4 ( .A(signal_4142), .B(cell_2122_and_out[1]), .Z(
        signal_4148) );
  XOR2_X1 cell_2122_U3 ( .A(signal_2384), .B(cell_2122_and_out[0]), .Z(
        signal_1403) );
  XOR2_X1 cell_2122_U2 ( .A(signal_4142), .B(signal_4133), .Z(
        cell_2122_and_in[1]) );
  XOR2_X1 cell_2122_U1 ( .A(signal_2384), .B(signal_2375), .Z(
        cell_2122_and_in[0]) );
  XOR2_X1 cell_2122_a_HPC2_and_U14 ( .A(Fresh[408]), .B(cell_2122_and_in[0]), 
        .Z(cell_2122_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2122_a_HPC2_and_U13 ( .A(Fresh[408]), .B(cell_2122_and_in[1]), 
        .Z(cell_2122_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2122_a_HPC2_and_U12 ( .A1(cell_2122_a_HPC2_and_a_reg[1]), .A2(
        cell_2122_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2122_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2122_a_HPC2_and_U11 ( .A1(cell_2122_a_HPC2_and_a_reg[0]), .A2(
        cell_2122_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2122_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2122_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2122_a_HPC2_and_n9), .ZN(cell_2122_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2122_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2122_a_HPC2_and_n9), .ZN(cell_2122_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2122_a_HPC2_and_U8 ( .A(Fresh[408]), .ZN(cell_2122_a_HPC2_and_n9) );
  AND2_X1 cell_2122_a_HPC2_and_U7 ( .A1(cell_2122_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2122_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2122_a_HPC2_and_U6 ( .A1(cell_2122_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2122_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2122_a_HPC2_and_U5 ( .A(cell_2122_a_HPC2_and_n8), .B(
        cell_2122_a_HPC2_and_z_1__1_), .ZN(cell_2122_and_out[1]) );
  XNOR2_X1 cell_2122_a_HPC2_and_U4 ( .A(
        cell_2122_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2122_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2122_a_HPC2_and_n8) );
  XNOR2_X1 cell_2122_a_HPC2_and_U3 ( .A(cell_2122_a_HPC2_and_n7), .B(
        cell_2122_a_HPC2_and_z_0__0_), .ZN(cell_2122_and_out[0]) );
  XNOR2_X1 cell_2122_a_HPC2_and_U2 ( .A(
        cell_2122_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2122_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2122_a_HPC2_and_n7) );
  DFF_X1 cell_2122_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2122_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2122_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2122_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2122_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2122_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2122_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2122_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2122_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2122_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2123_U4 ( .A(signal_4136), .B(cell_2123_and_out[1]), .Z(
        signal_4149) );
  XOR2_X1 cell_2123_U3 ( .A(signal_2378), .B(cell_2123_and_out[0]), .Z(
        signal_1398) );
  XOR2_X1 cell_2123_U2 ( .A(signal_4136), .B(signal_4143), .Z(
        cell_2123_and_in[1]) );
  XOR2_X1 cell_2123_U1 ( .A(signal_2378), .B(signal_2385), .Z(
        cell_2123_and_in[0]) );
  XOR2_X1 cell_2123_a_HPC2_and_U14 ( .A(Fresh[409]), .B(cell_2123_and_in[0]), 
        .Z(cell_2123_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2123_a_HPC2_and_U13 ( .A(Fresh[409]), .B(cell_2123_and_in[1]), 
        .Z(cell_2123_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2123_a_HPC2_and_U12 ( .A1(cell_2123_a_HPC2_and_a_reg[1]), .A2(
        cell_2123_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2123_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2123_a_HPC2_and_U11 ( .A1(cell_2123_a_HPC2_and_a_reg[0]), .A2(
        cell_2123_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2123_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2123_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2123_a_HPC2_and_n9), .ZN(cell_2123_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2123_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2123_a_HPC2_and_n9), .ZN(cell_2123_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2123_a_HPC2_and_U8 ( .A(Fresh[409]), .ZN(cell_2123_a_HPC2_and_n9) );
  AND2_X1 cell_2123_a_HPC2_and_U7 ( .A1(cell_2123_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2123_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2123_a_HPC2_and_U6 ( .A1(cell_2123_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2123_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2123_a_HPC2_and_U5 ( .A(cell_2123_a_HPC2_and_n8), .B(
        cell_2123_a_HPC2_and_z_1__1_), .ZN(cell_2123_and_out[1]) );
  XNOR2_X1 cell_2123_a_HPC2_and_U4 ( .A(
        cell_2123_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2123_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2123_a_HPC2_and_n8) );
  XNOR2_X1 cell_2123_a_HPC2_and_U3 ( .A(cell_2123_a_HPC2_and_n7), .B(
        cell_2123_a_HPC2_and_z_0__0_), .ZN(cell_2123_and_out[0]) );
  XNOR2_X1 cell_2123_a_HPC2_and_U2 ( .A(
        cell_2123_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2123_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2123_a_HPC2_and_n7) );
  DFF_X1 cell_2123_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2123_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2123_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2123_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2123_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2123_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2123_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2123_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2123_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2123_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2124_U4 ( .A(signal_4140), .B(cell_2124_and_out[1]), .Z(
        signal_4150) );
  XOR2_X1 cell_2124_U3 ( .A(signal_2382), .B(cell_2124_and_out[0]), .Z(
        signal_1402) );
  XOR2_X1 cell_2124_U2 ( .A(signal_4140), .B(signal_4130), .Z(
        cell_2124_and_in[1]) );
  XOR2_X1 cell_2124_U1 ( .A(signal_2382), .B(signal_2372), .Z(
        cell_2124_and_in[0]) );
  XOR2_X1 cell_2124_a_HPC2_and_U14 ( .A(Fresh[410]), .B(cell_2124_and_in[0]), 
        .Z(cell_2124_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2124_a_HPC2_and_U13 ( .A(Fresh[410]), .B(cell_2124_and_in[1]), 
        .Z(cell_2124_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2124_a_HPC2_and_U12 ( .A1(cell_2124_a_HPC2_and_a_reg[1]), .A2(
        cell_2124_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2124_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2124_a_HPC2_and_U11 ( .A1(cell_2124_a_HPC2_and_a_reg[0]), .A2(
        cell_2124_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2124_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2124_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2124_a_HPC2_and_n9), .ZN(cell_2124_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2124_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2124_a_HPC2_and_n9), .ZN(cell_2124_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2124_a_HPC2_and_U8 ( .A(Fresh[410]), .ZN(cell_2124_a_HPC2_and_n9) );
  AND2_X1 cell_2124_a_HPC2_and_U7 ( .A1(cell_2124_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2124_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2124_a_HPC2_and_U6 ( .A1(cell_2124_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2124_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2124_a_HPC2_and_U5 ( .A(cell_2124_a_HPC2_and_n8), .B(
        cell_2124_a_HPC2_and_z_1__1_), .ZN(cell_2124_and_out[1]) );
  XNOR2_X1 cell_2124_a_HPC2_and_U4 ( .A(
        cell_2124_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2124_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2124_a_HPC2_and_n8) );
  XNOR2_X1 cell_2124_a_HPC2_and_U3 ( .A(cell_2124_a_HPC2_and_n7), .B(
        cell_2124_a_HPC2_and_z_0__0_), .ZN(cell_2124_and_out[0]) );
  XNOR2_X1 cell_2124_a_HPC2_and_U2 ( .A(
        cell_2124_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2124_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2124_a_HPC2_and_n7) );
  DFF_X1 cell_2124_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2124_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2124_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2124_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2124_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2124_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2124_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2124_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2124_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2124_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2125_U4 ( .A(signal_4138), .B(cell_2125_and_out[1]), .Z(
        signal_4151) );
  XOR2_X1 cell_2125_U3 ( .A(signal_2380), .B(cell_2125_and_out[0]), .Z(
        signal_1404) );
  XOR2_X1 cell_2125_U2 ( .A(signal_4138), .B(signal_4137), .Z(
        cell_2125_and_in[1]) );
  XOR2_X1 cell_2125_U1 ( .A(signal_2380), .B(signal_2379), .Z(
        cell_2125_and_in[0]) );
  XOR2_X1 cell_2125_a_HPC2_and_U14 ( .A(Fresh[411]), .B(cell_2125_and_in[0]), 
        .Z(cell_2125_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2125_a_HPC2_and_U13 ( .A(Fresh[411]), .B(cell_2125_and_in[1]), 
        .Z(cell_2125_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2125_a_HPC2_and_U12 ( .A1(cell_2125_a_HPC2_and_a_reg[1]), .A2(
        cell_2125_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2125_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2125_a_HPC2_and_U11 ( .A1(cell_2125_a_HPC2_and_a_reg[0]), .A2(
        cell_2125_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2125_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2125_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2125_a_HPC2_and_n9), .ZN(cell_2125_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2125_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2125_a_HPC2_and_n9), .ZN(cell_2125_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2125_a_HPC2_and_U8 ( .A(Fresh[411]), .ZN(cell_2125_a_HPC2_and_n9) );
  AND2_X1 cell_2125_a_HPC2_and_U7 ( .A1(cell_2125_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2125_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2125_a_HPC2_and_U6 ( .A1(cell_2125_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2125_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2125_a_HPC2_and_U5 ( .A(cell_2125_a_HPC2_and_n8), .B(
        cell_2125_a_HPC2_and_z_1__1_), .ZN(cell_2125_and_out[1]) );
  XNOR2_X1 cell_2125_a_HPC2_and_U4 ( .A(
        cell_2125_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2125_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2125_a_HPC2_and_n8) );
  XNOR2_X1 cell_2125_a_HPC2_and_U3 ( .A(cell_2125_a_HPC2_and_n7), .B(
        cell_2125_a_HPC2_and_z_0__0_), .ZN(cell_2125_and_out[0]) );
  XNOR2_X1 cell_2125_a_HPC2_and_U2 ( .A(
        cell_2125_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2125_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2125_a_HPC2_and_n7) );
  DFF_X1 cell_2125_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2125_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2125_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2125_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2125_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2125_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2125_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2125_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2125_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2125_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2126_U4 ( .A(signal_4131), .B(cell_2126_and_out[1]), .Z(
        signal_4152) );
  XOR2_X1 cell_2126_U3 ( .A(signal_2373), .B(cell_2126_and_out[0]), .Z(
        signal_1401) );
  XOR2_X1 cell_2126_U2 ( .A(signal_4131), .B(signal_4139), .Z(
        cell_2126_and_in[1]) );
  XOR2_X1 cell_2126_U1 ( .A(signal_2373), .B(signal_2381), .Z(
        cell_2126_and_in[0]) );
  XOR2_X1 cell_2126_a_HPC2_and_U14 ( .A(Fresh[412]), .B(cell_2126_and_in[0]), 
        .Z(cell_2126_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2126_a_HPC2_and_U13 ( .A(Fresh[412]), .B(cell_2126_and_in[1]), 
        .Z(cell_2126_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2126_a_HPC2_and_U12 ( .A1(cell_2126_a_HPC2_and_a_reg[1]), .A2(
        cell_2126_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2126_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2126_a_HPC2_and_U11 ( .A1(cell_2126_a_HPC2_and_a_reg[0]), .A2(
        cell_2126_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2126_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2126_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2126_a_HPC2_and_n9), .ZN(cell_2126_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2126_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2126_a_HPC2_and_n9), .ZN(cell_2126_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2126_a_HPC2_and_U8 ( .A(Fresh[412]), .ZN(cell_2126_a_HPC2_and_n9) );
  AND2_X1 cell_2126_a_HPC2_and_U7 ( .A1(cell_2126_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2126_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2126_a_HPC2_and_U6 ( .A1(cell_2126_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2126_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2126_a_HPC2_and_U5 ( .A(cell_2126_a_HPC2_and_n8), .B(
        cell_2126_a_HPC2_and_z_1__1_), .ZN(cell_2126_and_out[1]) );
  XNOR2_X1 cell_2126_a_HPC2_and_U4 ( .A(
        cell_2126_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2126_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2126_a_HPC2_and_n8) );
  XNOR2_X1 cell_2126_a_HPC2_and_U3 ( .A(cell_2126_a_HPC2_and_n7), .B(
        cell_2126_a_HPC2_and_z_0__0_), .ZN(cell_2126_and_out[0]) );
  XNOR2_X1 cell_2126_a_HPC2_and_U2 ( .A(
        cell_2126_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2126_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2126_a_HPC2_and_n7) );
  DFF_X1 cell_2126_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2126_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2126_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2126_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2126_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2126_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2126_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2126_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2126_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2126_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  XOR2_X1 cell_2127_U4 ( .A(signal_4132), .B(cell_2127_and_out[1]), .Z(
        signal_4153) );
  XOR2_X1 cell_2127_U3 ( .A(signal_2374), .B(cell_2127_and_out[0]), .Z(
        signal_1400) );
  XOR2_X1 cell_2127_U2 ( .A(signal_4132), .B(signal_4144), .Z(
        cell_2127_and_in[1]) );
  XOR2_X1 cell_2127_U1 ( .A(signal_2374), .B(signal_2386), .Z(
        cell_2127_and_in[0]) );
  XOR2_X1 cell_2127_a_HPC2_and_U14 ( .A(Fresh[413]), .B(cell_2127_and_in[0]), 
        .Z(cell_2127_a_HPC2_and_s_in_1__0_) );
  XOR2_X1 cell_2127_a_HPC2_and_U13 ( .A(Fresh[413]), .B(cell_2127_and_in[1]), 
        .Z(cell_2127_a_HPC2_and_s_in_0__1_) );
  AND2_X1 cell_2127_a_HPC2_and_U12 ( .A1(cell_2127_a_HPC2_and_a_reg[1]), .A2(
        cell_2127_a_HPC2_and_s_out_1__0_), .ZN(
        cell_2127_a_HPC2_and_p_1_in_1__0_) );
  AND2_X1 cell_2127_a_HPC2_and_U11 ( .A1(cell_2127_a_HPC2_and_a_reg[0]), .A2(
        cell_2127_a_HPC2_and_s_out_0__1_), .ZN(
        cell_2127_a_HPC2_and_p_1_in_0__1_) );
  NOR2_X1 cell_2127_a_HPC2_and_U10 ( .A1(signal_3236), .A2(
        cell_2127_a_HPC2_and_n9), .ZN(cell_2127_a_HPC2_and_p_0_in_1__0_) );
  NOR2_X1 cell_2127_a_HPC2_and_U9 ( .A1(signal_1513), .A2(
        cell_2127_a_HPC2_and_n9), .ZN(cell_2127_a_HPC2_and_p_0_in_0__1_) );
  INV_X1 cell_2127_a_HPC2_and_U8 ( .A(Fresh[413]), .ZN(cell_2127_a_HPC2_and_n9) );
  AND2_X1 cell_2127_a_HPC2_and_U7 ( .A1(cell_2127_and_in[1]), .A2(signal_3236), 
        .ZN(cell_2127_a_HPC2_and_mul[1]) );
  AND2_X1 cell_2127_a_HPC2_and_U6 ( .A1(cell_2127_and_in[0]), .A2(signal_1513), 
        .ZN(cell_2127_a_HPC2_and_mul[0]) );
  XNOR2_X1 cell_2127_a_HPC2_and_U5 ( .A(cell_2127_a_HPC2_and_n8), .B(
        cell_2127_a_HPC2_and_z_1__1_), .ZN(cell_2127_and_out[1]) );
  XNOR2_X1 cell_2127_a_HPC2_and_U4 ( .A(
        cell_2127_a_HPC2_and_p_0_pipe_out_1__0_), .B(
        cell_2127_a_HPC2_and_p_1_out_1__0_), .ZN(cell_2127_a_HPC2_and_n8) );
  XNOR2_X1 cell_2127_a_HPC2_and_U3 ( .A(cell_2127_a_HPC2_and_n7), .B(
        cell_2127_a_HPC2_and_z_0__0_), .ZN(cell_2127_and_out[0]) );
  XNOR2_X1 cell_2127_a_HPC2_and_U2 ( .A(
        cell_2127_a_HPC2_and_p_0_pipe_out_0__1_), .B(
        cell_2127_a_HPC2_and_p_1_out_0__1_), .ZN(cell_2127_a_HPC2_and_n7) );
  DFF_X1 cell_2127_a_HPC2_and_mul_pipe_s1_0_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_mul[0]), .CK(clk), .Q(
        cell_2127_a_HPC2_and_mul_s1_out[0]), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_mul_pipe_s2_0_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_mul_s1_out[0]), .CK(clk), .Q(
        cell_2127_a_HPC2_and_z_0__0_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_a_i_0_s_current_state_reg ( .D(signal_1513), 
        .CK(clk), .Q(cell_2127_a_HPC2_and_a_reg[0]), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_s_reg_0_1_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_s_in_0__1_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_s_out_0__1_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_p_0_reg_0_1_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_p_0_in_0__1_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_p_0_out_0__1_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_p_1_reg_0_1_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_p_1_in_0__1_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_p_1_out_0__1_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_p_0_pipe_0_1_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_p_0_out_0__1_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_p_0_pipe_out_0__1_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_mul_pipe_s1_1_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_mul[1]), .CK(clk), .Q(
        cell_2127_a_HPC2_and_mul_s1_out[1]), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_mul_pipe_s2_1_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_mul_s1_out[1]), .CK(clk), .Q(
        cell_2127_a_HPC2_and_z_1__1_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_a_i_1_s_current_state_reg ( .D(signal_3236), 
        .CK(clk), .Q(cell_2127_a_HPC2_and_a_reg[1]), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_s_reg_1_0_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_s_in_1__0_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_s_out_1__0_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_p_0_reg_1_0_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_p_0_in_1__0_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_p_0_out_1__0_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_p_1_reg_1_0_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_p_1_in_1__0_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_p_1_out_1__0_), .QN() );
  DFF_X1 cell_2127_a_HPC2_and_p_0_pipe_1_0_s_current_state_reg ( .D(
        cell_2127_a_HPC2_and_p_0_out_1__0_), .CK(clk), .Q(
        cell_2127_a_HPC2_and_p_0_pipe_out_1__0_), .QN() );
  DFF_X1 cell_87_s_reg_0_s_current_state_reg ( .D(signal_465), .CK(signal_4640), .Q(ciphertext_s0[120]), .QN() );
  DFF_X1 cell_87_s_reg_1_s_current_state_reg ( .D(signal_3786), .CK(
        signal_4640), .Q(ciphertext_s1[120]), .QN() );
  DFF_X1 cell_90_s_reg_0_s_current_state_reg ( .D(signal_467), .CK(signal_4640), .Q(ciphertext_s0[121]), .QN() );
  DFF_X1 cell_90_s_reg_1_s_current_state_reg ( .D(signal_3787), .CK(
        signal_4640), .Q(ciphertext_s1[121]), .QN() );
  DFF_X1 cell_93_s_reg_0_s_current_state_reg ( .D(signal_469), .CK(signal_4640), .Q(ciphertext_s0[122]), .QN() );
  DFF_X1 cell_93_s_reg_1_s_current_state_reg ( .D(signal_3788), .CK(
        signal_4640), .Q(ciphertext_s1[122]), .QN() );
  DFF_X1 cell_96_s_reg_0_s_current_state_reg ( .D(signal_471), .CK(signal_4640), .Q(ciphertext_s0[123]), .QN() );
  DFF_X1 cell_96_s_reg_1_s_current_state_reg ( .D(signal_3789), .CK(
        signal_4640), .Q(ciphertext_s1[123]), .QN() );
  DFF_X1 cell_99_s_reg_0_s_current_state_reg ( .D(signal_473), .CK(signal_4640), .Q(ciphertext_s0[124]), .QN() );
  DFF_X1 cell_99_s_reg_1_s_current_state_reg ( .D(signal_3790), .CK(
        signal_4640), .Q(ciphertext_s1[124]), .QN() );
  DFF_X1 cell_102_s_reg_0_s_current_state_reg ( .D(signal_475), .CK(
        signal_4640), .Q(ciphertext_s0[125]), .QN() );
  DFF_X1 cell_102_s_reg_1_s_current_state_reg ( .D(signal_3791), .CK(
        signal_4640), .Q(ciphertext_s1[125]), .QN() );
  DFF_X1 cell_105_s_reg_0_s_current_state_reg ( .D(signal_477), .CK(
        signal_4640), .Q(ciphertext_s0[126]), .QN() );
  DFF_X1 cell_105_s_reg_1_s_current_state_reg ( .D(signal_3792), .CK(
        signal_4640), .Q(ciphertext_s1[126]), .QN() );
  DFF_X1 cell_108_s_reg_0_s_current_state_reg ( .D(signal_479), .CK(
        signal_4640), .Q(ciphertext_s0[127]), .QN() );
  DFF_X1 cell_108_s_reg_1_s_current_state_reg ( .D(signal_3793), .CK(
        signal_4640), .Q(ciphertext_s1[127]), .QN() );
  DFF_X1 cell_111_s_reg_0_s_current_state_reg ( .D(signal_481), .CK(
        signal_4640), .Q(ciphertext_s0[112]), .QN() );
  DFF_X1 cell_111_s_reg_1_s_current_state_reg ( .D(signal_3794), .CK(
        signal_4640), .Q(ciphertext_s1[112]), .QN() );
  DFF_X1 cell_114_s_reg_0_s_current_state_reg ( .D(signal_483), .CK(
        signal_4640), .Q(ciphertext_s0[113]), .QN() );
  DFF_X1 cell_114_s_reg_1_s_current_state_reg ( .D(signal_3795), .CK(
        signal_4640), .Q(ciphertext_s1[113]), .QN() );
  DFF_X1 cell_117_s_reg_0_s_current_state_reg ( .D(signal_485), .CK(
        signal_4640), .Q(ciphertext_s0[114]), .QN() );
  DFF_X1 cell_117_s_reg_1_s_current_state_reg ( .D(signal_3796), .CK(
        signal_4640), .Q(ciphertext_s1[114]), .QN() );
  DFF_X1 cell_120_s_reg_0_s_current_state_reg ( .D(signal_487), .CK(
        signal_4640), .Q(ciphertext_s0[115]), .QN() );
  DFF_X1 cell_120_s_reg_1_s_current_state_reg ( .D(signal_3797), .CK(
        signal_4640), .Q(ciphertext_s1[115]), .QN() );
  DFF_X1 cell_123_s_reg_0_s_current_state_reg ( .D(signal_489), .CK(
        signal_4640), .Q(ciphertext_s0[116]), .QN() );
  DFF_X1 cell_123_s_reg_1_s_current_state_reg ( .D(signal_3798), .CK(
        signal_4640), .Q(ciphertext_s1[116]), .QN() );
  DFF_X1 cell_126_s_reg_0_s_current_state_reg ( .D(signal_491), .CK(
        signal_4640), .Q(ciphertext_s0[117]), .QN() );
  DFF_X1 cell_126_s_reg_1_s_current_state_reg ( .D(signal_3799), .CK(
        signal_4640), .Q(ciphertext_s1[117]), .QN() );
  DFF_X1 cell_129_s_reg_0_s_current_state_reg ( .D(signal_493), .CK(
        signal_4640), .Q(ciphertext_s0[118]), .QN() );
  DFF_X1 cell_129_s_reg_1_s_current_state_reg ( .D(signal_3800), .CK(
        signal_4640), .Q(ciphertext_s1[118]), .QN() );
  DFF_X1 cell_132_s_reg_0_s_current_state_reg ( .D(signal_495), .CK(
        signal_4640), .Q(ciphertext_s0[119]), .QN() );
  DFF_X1 cell_132_s_reg_1_s_current_state_reg ( .D(signal_3801), .CK(
        signal_4640), .Q(ciphertext_s1[119]), .QN() );
  DFF_X1 cell_135_s_reg_0_s_current_state_reg ( .D(signal_497), .CK(
        signal_4640), .Q(ciphertext_s0[104]), .QN() );
  DFF_X1 cell_135_s_reg_1_s_current_state_reg ( .D(signal_3802), .CK(
        signal_4640), .Q(ciphertext_s1[104]), .QN() );
  DFF_X1 cell_138_s_reg_0_s_current_state_reg ( .D(signal_499), .CK(
        signal_4640), .Q(ciphertext_s0[105]), .QN() );
  DFF_X1 cell_138_s_reg_1_s_current_state_reg ( .D(signal_3803), .CK(
        signal_4640), .Q(ciphertext_s1[105]), .QN() );
  DFF_X1 cell_141_s_reg_0_s_current_state_reg ( .D(signal_501), .CK(
        signal_4640), .Q(ciphertext_s0[106]), .QN() );
  DFF_X1 cell_141_s_reg_1_s_current_state_reg ( .D(signal_3804), .CK(
        signal_4640), .Q(ciphertext_s1[106]), .QN() );
  DFF_X1 cell_144_s_reg_0_s_current_state_reg ( .D(signal_503), .CK(
        signal_4640), .Q(ciphertext_s0[107]), .QN() );
  DFF_X1 cell_144_s_reg_1_s_current_state_reg ( .D(signal_3805), .CK(
        signal_4640), .Q(ciphertext_s1[107]), .QN() );
  DFF_X1 cell_147_s_reg_0_s_current_state_reg ( .D(signal_505), .CK(
        signal_4640), .Q(ciphertext_s0[108]), .QN() );
  DFF_X1 cell_147_s_reg_1_s_current_state_reg ( .D(signal_3806), .CK(
        signal_4640), .Q(ciphertext_s1[108]), .QN() );
  DFF_X1 cell_150_s_reg_0_s_current_state_reg ( .D(signal_507), .CK(
        signal_4640), .Q(ciphertext_s0[109]), .QN() );
  DFF_X1 cell_150_s_reg_1_s_current_state_reg ( .D(signal_3807), .CK(
        signal_4640), .Q(ciphertext_s1[109]), .QN() );
  DFF_X1 cell_153_s_reg_0_s_current_state_reg ( .D(signal_509), .CK(
        signal_4640), .Q(ciphertext_s0[110]), .QN() );
  DFF_X1 cell_153_s_reg_1_s_current_state_reg ( .D(signal_3808), .CK(
        signal_4640), .Q(ciphertext_s1[110]), .QN() );
  DFF_X1 cell_156_s_reg_0_s_current_state_reg ( .D(signal_511), .CK(
        signal_4640), .Q(ciphertext_s0[111]), .QN() );
  DFF_X1 cell_156_s_reg_1_s_current_state_reg ( .D(signal_3809), .CK(
        signal_4640), .Q(ciphertext_s1[111]), .QN() );
  DFF_X1 cell_159_s_reg_0_s_current_state_reg ( .D(signal_513), .CK(
        signal_4640), .Q(ciphertext_s0[96]), .QN() );
  DFF_X1 cell_159_s_reg_1_s_current_state_reg ( .D(signal_3810), .CK(
        signal_4640), .Q(ciphertext_s1[96]), .QN() );
  DFF_X1 cell_162_s_reg_0_s_current_state_reg ( .D(signal_515), .CK(
        signal_4640), .Q(ciphertext_s0[97]), .QN() );
  DFF_X1 cell_162_s_reg_1_s_current_state_reg ( .D(signal_3811), .CK(
        signal_4640), .Q(ciphertext_s1[97]), .QN() );
  DFF_X1 cell_165_s_reg_0_s_current_state_reg ( .D(signal_517), .CK(
        signal_4640), .Q(ciphertext_s0[98]), .QN() );
  DFF_X1 cell_165_s_reg_1_s_current_state_reg ( .D(signal_3812), .CK(
        signal_4640), .Q(ciphertext_s1[98]), .QN() );
  DFF_X1 cell_168_s_reg_0_s_current_state_reg ( .D(signal_519), .CK(
        signal_4640), .Q(ciphertext_s0[99]), .QN() );
  DFF_X1 cell_168_s_reg_1_s_current_state_reg ( .D(signal_3813), .CK(
        signal_4640), .Q(ciphertext_s1[99]), .QN() );
  DFF_X1 cell_171_s_reg_0_s_current_state_reg ( .D(signal_521), .CK(
        signal_4640), .Q(ciphertext_s0[100]), .QN() );
  DFF_X1 cell_171_s_reg_1_s_current_state_reg ( .D(signal_3814), .CK(
        signal_4640), .Q(ciphertext_s1[100]), .QN() );
  DFF_X1 cell_174_s_reg_0_s_current_state_reg ( .D(signal_523), .CK(
        signal_4640), .Q(ciphertext_s0[101]), .QN() );
  DFF_X1 cell_174_s_reg_1_s_current_state_reg ( .D(signal_3815), .CK(
        signal_4640), .Q(ciphertext_s1[101]), .QN() );
  DFF_X1 cell_177_s_reg_0_s_current_state_reg ( .D(signal_525), .CK(
        signal_4640), .Q(ciphertext_s0[102]), .QN() );
  DFF_X1 cell_177_s_reg_1_s_current_state_reg ( .D(signal_3816), .CK(
        signal_4640), .Q(ciphertext_s1[102]), .QN() );
  DFF_X1 cell_180_s_reg_0_s_current_state_reg ( .D(signal_527), .CK(
        signal_4640), .Q(ciphertext_s0[103]), .QN() );
  DFF_X1 cell_180_s_reg_1_s_current_state_reg ( .D(signal_3817), .CK(
        signal_4640), .Q(ciphertext_s1[103]), .QN() );
  DFF_X1 cell_183_s_reg_0_s_current_state_reg ( .D(signal_529), .CK(
        signal_4640), .Q(ciphertext_s0[88]), .QN() );
  DFF_X1 cell_183_s_reg_1_s_current_state_reg ( .D(signal_3818), .CK(
        signal_4640), .Q(ciphertext_s1[88]), .QN() );
  DFF_X1 cell_186_s_reg_0_s_current_state_reg ( .D(signal_531), .CK(
        signal_4640), .Q(ciphertext_s0[89]), .QN() );
  DFF_X1 cell_186_s_reg_1_s_current_state_reg ( .D(signal_3819), .CK(
        signal_4640), .Q(ciphertext_s1[89]), .QN() );
  DFF_X1 cell_189_s_reg_0_s_current_state_reg ( .D(signal_533), .CK(
        signal_4640), .Q(ciphertext_s0[90]), .QN() );
  DFF_X1 cell_189_s_reg_1_s_current_state_reg ( .D(signal_3820), .CK(
        signal_4640), .Q(ciphertext_s1[90]), .QN() );
  DFF_X1 cell_192_s_reg_0_s_current_state_reg ( .D(signal_535), .CK(
        signal_4640), .Q(ciphertext_s0[91]), .QN() );
  DFF_X1 cell_192_s_reg_1_s_current_state_reg ( .D(signal_3821), .CK(
        signal_4640), .Q(ciphertext_s1[91]), .QN() );
  DFF_X1 cell_195_s_reg_0_s_current_state_reg ( .D(signal_537), .CK(
        signal_4640), .Q(ciphertext_s0[92]), .QN() );
  DFF_X1 cell_195_s_reg_1_s_current_state_reg ( .D(signal_3822), .CK(
        signal_4640), .Q(ciphertext_s1[92]), .QN() );
  DFF_X1 cell_198_s_reg_0_s_current_state_reg ( .D(signal_539), .CK(
        signal_4640), .Q(ciphertext_s0[93]), .QN() );
  DFF_X1 cell_198_s_reg_1_s_current_state_reg ( .D(signal_3823), .CK(
        signal_4640), .Q(ciphertext_s1[93]), .QN() );
  DFF_X1 cell_201_s_reg_0_s_current_state_reg ( .D(signal_541), .CK(
        signal_4640), .Q(ciphertext_s0[94]), .QN() );
  DFF_X1 cell_201_s_reg_1_s_current_state_reg ( .D(signal_3824), .CK(
        signal_4640), .Q(ciphertext_s1[94]), .QN() );
  DFF_X1 cell_204_s_reg_0_s_current_state_reg ( .D(signal_543), .CK(
        signal_4640), .Q(ciphertext_s0[95]), .QN() );
  DFF_X1 cell_204_s_reg_1_s_current_state_reg ( .D(signal_3825), .CK(
        signal_4640), .Q(ciphertext_s1[95]), .QN() );
  DFF_X1 cell_207_s_reg_0_s_current_state_reg ( .D(signal_545), .CK(
        signal_4640), .Q(ciphertext_s0[80]), .QN() );
  DFF_X1 cell_207_s_reg_1_s_current_state_reg ( .D(signal_3826), .CK(
        signal_4640), .Q(ciphertext_s1[80]), .QN() );
  DFF_X1 cell_210_s_reg_0_s_current_state_reg ( .D(signal_547), .CK(
        signal_4640), .Q(ciphertext_s0[81]), .QN() );
  DFF_X1 cell_210_s_reg_1_s_current_state_reg ( .D(signal_3827), .CK(
        signal_4640), .Q(ciphertext_s1[81]), .QN() );
  DFF_X1 cell_213_s_reg_0_s_current_state_reg ( .D(signal_549), .CK(
        signal_4640), .Q(ciphertext_s0[82]), .QN() );
  DFF_X1 cell_213_s_reg_1_s_current_state_reg ( .D(signal_3828), .CK(
        signal_4640), .Q(ciphertext_s1[82]), .QN() );
  DFF_X1 cell_216_s_reg_0_s_current_state_reg ( .D(signal_551), .CK(
        signal_4640), .Q(ciphertext_s0[83]), .QN() );
  DFF_X1 cell_216_s_reg_1_s_current_state_reg ( .D(signal_3829), .CK(
        signal_4640), .Q(ciphertext_s1[83]), .QN() );
  DFF_X1 cell_219_s_reg_0_s_current_state_reg ( .D(signal_553), .CK(
        signal_4640), .Q(ciphertext_s0[84]), .QN() );
  DFF_X1 cell_219_s_reg_1_s_current_state_reg ( .D(signal_3830), .CK(
        signal_4640), .Q(ciphertext_s1[84]), .QN() );
  DFF_X1 cell_222_s_reg_0_s_current_state_reg ( .D(signal_555), .CK(
        signal_4640), .Q(ciphertext_s0[85]), .QN() );
  DFF_X1 cell_222_s_reg_1_s_current_state_reg ( .D(signal_3831), .CK(
        signal_4640), .Q(ciphertext_s1[85]), .QN() );
  DFF_X1 cell_225_s_reg_0_s_current_state_reg ( .D(signal_557), .CK(
        signal_4640), .Q(ciphertext_s0[86]), .QN() );
  DFF_X1 cell_225_s_reg_1_s_current_state_reg ( .D(signal_3832), .CK(
        signal_4640), .Q(ciphertext_s1[86]), .QN() );
  DFF_X1 cell_228_s_reg_0_s_current_state_reg ( .D(signal_559), .CK(
        signal_4640), .Q(ciphertext_s0[87]), .QN() );
  DFF_X1 cell_228_s_reg_1_s_current_state_reg ( .D(signal_3833), .CK(
        signal_4640), .Q(ciphertext_s1[87]), .QN() );
  DFF_X1 cell_231_s_reg_0_s_current_state_reg ( .D(signal_561), .CK(
        signal_4640), .Q(ciphertext_s0[72]), .QN() );
  DFF_X1 cell_231_s_reg_1_s_current_state_reg ( .D(signal_3834), .CK(
        signal_4640), .Q(ciphertext_s1[72]), .QN() );
  DFF_X1 cell_234_s_reg_0_s_current_state_reg ( .D(signal_563), .CK(
        signal_4640), .Q(ciphertext_s0[73]), .QN() );
  DFF_X1 cell_234_s_reg_1_s_current_state_reg ( .D(signal_3835), .CK(
        signal_4640), .Q(ciphertext_s1[73]), .QN() );
  DFF_X1 cell_237_s_reg_0_s_current_state_reg ( .D(signal_565), .CK(
        signal_4640), .Q(ciphertext_s0[74]), .QN() );
  DFF_X1 cell_237_s_reg_1_s_current_state_reg ( .D(signal_3836), .CK(
        signal_4640), .Q(ciphertext_s1[74]), .QN() );
  DFF_X1 cell_240_s_reg_0_s_current_state_reg ( .D(signal_567), .CK(
        signal_4640), .Q(ciphertext_s0[75]), .QN() );
  DFF_X1 cell_240_s_reg_1_s_current_state_reg ( .D(signal_3837), .CK(
        signal_4640), .Q(ciphertext_s1[75]), .QN() );
  DFF_X1 cell_243_s_reg_0_s_current_state_reg ( .D(signal_569), .CK(
        signal_4640), .Q(ciphertext_s0[76]), .QN() );
  DFF_X1 cell_243_s_reg_1_s_current_state_reg ( .D(signal_3838), .CK(
        signal_4640), .Q(ciphertext_s1[76]), .QN() );
  DFF_X1 cell_246_s_reg_0_s_current_state_reg ( .D(signal_571), .CK(
        signal_4640), .Q(ciphertext_s0[77]), .QN() );
  DFF_X1 cell_246_s_reg_1_s_current_state_reg ( .D(signal_3839), .CK(
        signal_4640), .Q(ciphertext_s1[77]), .QN() );
  DFF_X1 cell_249_s_reg_0_s_current_state_reg ( .D(signal_573), .CK(
        signal_4640), .Q(ciphertext_s0[78]), .QN() );
  DFF_X1 cell_249_s_reg_1_s_current_state_reg ( .D(signal_3840), .CK(
        signal_4640), .Q(ciphertext_s1[78]), .QN() );
  DFF_X1 cell_252_s_reg_0_s_current_state_reg ( .D(signal_575), .CK(
        signal_4640), .Q(ciphertext_s0[79]), .QN() );
  DFF_X1 cell_252_s_reg_1_s_current_state_reg ( .D(signal_3841), .CK(
        signal_4640), .Q(ciphertext_s1[79]), .QN() );
  DFF_X1 cell_255_s_reg_0_s_current_state_reg ( .D(signal_577), .CK(
        signal_4640), .Q(ciphertext_s0[64]), .QN() );
  DFF_X1 cell_255_s_reg_1_s_current_state_reg ( .D(signal_3842), .CK(
        signal_4640), .Q(ciphertext_s1[64]), .QN() );
  DFF_X1 cell_258_s_reg_0_s_current_state_reg ( .D(signal_579), .CK(
        signal_4640), .Q(ciphertext_s0[65]), .QN() );
  DFF_X1 cell_258_s_reg_1_s_current_state_reg ( .D(signal_3843), .CK(
        signal_4640), .Q(ciphertext_s1[65]), .QN() );
  DFF_X1 cell_261_s_reg_0_s_current_state_reg ( .D(signal_581), .CK(
        signal_4640), .Q(ciphertext_s0[66]), .QN() );
  DFF_X1 cell_261_s_reg_1_s_current_state_reg ( .D(signal_3844), .CK(
        signal_4640), .Q(ciphertext_s1[66]), .QN() );
  DFF_X1 cell_264_s_reg_0_s_current_state_reg ( .D(signal_583), .CK(
        signal_4640), .Q(ciphertext_s0[67]), .QN() );
  DFF_X1 cell_264_s_reg_1_s_current_state_reg ( .D(signal_3845), .CK(
        signal_4640), .Q(ciphertext_s1[67]), .QN() );
  DFF_X1 cell_267_s_reg_0_s_current_state_reg ( .D(signal_585), .CK(
        signal_4640), .Q(ciphertext_s0[68]), .QN() );
  DFF_X1 cell_267_s_reg_1_s_current_state_reg ( .D(signal_3846), .CK(
        signal_4640), .Q(ciphertext_s1[68]), .QN() );
  DFF_X1 cell_270_s_reg_0_s_current_state_reg ( .D(signal_587), .CK(
        signal_4640), .Q(ciphertext_s0[69]), .QN() );
  DFF_X1 cell_270_s_reg_1_s_current_state_reg ( .D(signal_3847), .CK(
        signal_4640), .Q(ciphertext_s1[69]), .QN() );
  DFF_X1 cell_273_s_reg_0_s_current_state_reg ( .D(signal_589), .CK(
        signal_4640), .Q(ciphertext_s0[70]), .QN() );
  DFF_X1 cell_273_s_reg_1_s_current_state_reg ( .D(signal_3848), .CK(
        signal_4640), .Q(ciphertext_s1[70]), .QN() );
  DFF_X1 cell_276_s_reg_0_s_current_state_reg ( .D(signal_591), .CK(
        signal_4640), .Q(ciphertext_s0[71]), .QN() );
  DFF_X1 cell_276_s_reg_1_s_current_state_reg ( .D(signal_3849), .CK(
        signal_4640), .Q(ciphertext_s1[71]), .QN() );
  DFF_X1 cell_279_s_reg_0_s_current_state_reg ( .D(signal_593), .CK(
        signal_4640), .Q(ciphertext_s0[56]), .QN() );
  DFF_X1 cell_279_s_reg_1_s_current_state_reg ( .D(signal_3850), .CK(
        signal_4640), .Q(ciphertext_s1[56]), .QN() );
  DFF_X1 cell_282_s_reg_0_s_current_state_reg ( .D(signal_595), .CK(
        signal_4640), .Q(ciphertext_s0[57]), .QN() );
  DFF_X1 cell_282_s_reg_1_s_current_state_reg ( .D(signal_3851), .CK(
        signal_4640), .Q(ciphertext_s1[57]), .QN() );
  DFF_X1 cell_285_s_reg_0_s_current_state_reg ( .D(signal_597), .CK(
        signal_4640), .Q(ciphertext_s0[58]), .QN() );
  DFF_X1 cell_285_s_reg_1_s_current_state_reg ( .D(signal_3852), .CK(
        signal_4640), .Q(ciphertext_s1[58]), .QN() );
  DFF_X1 cell_288_s_reg_0_s_current_state_reg ( .D(signal_599), .CK(
        signal_4640), .Q(ciphertext_s0[59]), .QN() );
  DFF_X1 cell_288_s_reg_1_s_current_state_reg ( .D(signal_3853), .CK(
        signal_4640), .Q(ciphertext_s1[59]), .QN() );
  DFF_X1 cell_291_s_reg_0_s_current_state_reg ( .D(signal_601), .CK(
        signal_4640), .Q(ciphertext_s0[60]), .QN() );
  DFF_X1 cell_291_s_reg_1_s_current_state_reg ( .D(signal_3854), .CK(
        signal_4640), .Q(ciphertext_s1[60]), .QN() );
  DFF_X1 cell_294_s_reg_0_s_current_state_reg ( .D(signal_603), .CK(
        signal_4640), .Q(ciphertext_s0[61]), .QN() );
  DFF_X1 cell_294_s_reg_1_s_current_state_reg ( .D(signal_3855), .CK(
        signal_4640), .Q(ciphertext_s1[61]), .QN() );
  DFF_X1 cell_297_s_reg_0_s_current_state_reg ( .D(signal_605), .CK(
        signal_4640), .Q(ciphertext_s0[62]), .QN() );
  DFF_X1 cell_297_s_reg_1_s_current_state_reg ( .D(signal_3856), .CK(
        signal_4640), .Q(ciphertext_s1[62]), .QN() );
  DFF_X1 cell_300_s_reg_0_s_current_state_reg ( .D(signal_607), .CK(
        signal_4640), .Q(ciphertext_s0[63]), .QN() );
  DFF_X1 cell_300_s_reg_1_s_current_state_reg ( .D(signal_3857), .CK(
        signal_4640), .Q(ciphertext_s1[63]), .QN() );
  DFF_X1 cell_303_s_reg_0_s_current_state_reg ( .D(signal_609), .CK(
        signal_4640), .Q(ciphertext_s0[48]), .QN() );
  DFF_X1 cell_303_s_reg_1_s_current_state_reg ( .D(signal_3858), .CK(
        signal_4640), .Q(ciphertext_s1[48]), .QN() );
  DFF_X1 cell_306_s_reg_0_s_current_state_reg ( .D(signal_611), .CK(
        signal_4640), .Q(ciphertext_s0[49]), .QN() );
  DFF_X1 cell_306_s_reg_1_s_current_state_reg ( .D(signal_3859), .CK(
        signal_4640), .Q(ciphertext_s1[49]), .QN() );
  DFF_X1 cell_309_s_reg_0_s_current_state_reg ( .D(signal_613), .CK(
        signal_4640), .Q(ciphertext_s0[50]), .QN() );
  DFF_X1 cell_309_s_reg_1_s_current_state_reg ( .D(signal_3860), .CK(
        signal_4640), .Q(ciphertext_s1[50]), .QN() );
  DFF_X1 cell_312_s_reg_0_s_current_state_reg ( .D(signal_615), .CK(
        signal_4640), .Q(ciphertext_s0[51]), .QN() );
  DFF_X1 cell_312_s_reg_1_s_current_state_reg ( .D(signal_3861), .CK(
        signal_4640), .Q(ciphertext_s1[51]), .QN() );
  DFF_X1 cell_315_s_reg_0_s_current_state_reg ( .D(signal_617), .CK(
        signal_4640), .Q(ciphertext_s0[52]), .QN() );
  DFF_X1 cell_315_s_reg_1_s_current_state_reg ( .D(signal_3862), .CK(
        signal_4640), .Q(ciphertext_s1[52]), .QN() );
  DFF_X1 cell_318_s_reg_0_s_current_state_reg ( .D(signal_619), .CK(
        signal_4640), .Q(ciphertext_s0[53]), .QN() );
  DFF_X1 cell_318_s_reg_1_s_current_state_reg ( .D(signal_3863), .CK(
        signal_4640), .Q(ciphertext_s1[53]), .QN() );
  DFF_X1 cell_321_s_reg_0_s_current_state_reg ( .D(signal_621), .CK(
        signal_4640), .Q(ciphertext_s0[54]), .QN() );
  DFF_X1 cell_321_s_reg_1_s_current_state_reg ( .D(signal_3864), .CK(
        signal_4640), .Q(ciphertext_s1[54]), .QN() );
  DFF_X1 cell_324_s_reg_0_s_current_state_reg ( .D(signal_623), .CK(
        signal_4640), .Q(ciphertext_s0[55]), .QN() );
  DFF_X1 cell_324_s_reg_1_s_current_state_reg ( .D(signal_3865), .CK(
        signal_4640), .Q(ciphertext_s1[55]), .QN() );
  DFF_X1 cell_327_s_reg_0_s_current_state_reg ( .D(signal_625), .CK(
        signal_4640), .Q(ciphertext_s0[40]), .QN() );
  DFF_X1 cell_327_s_reg_1_s_current_state_reg ( .D(signal_3866), .CK(
        signal_4640), .Q(ciphertext_s1[40]), .QN() );
  DFF_X1 cell_330_s_reg_0_s_current_state_reg ( .D(signal_627), .CK(
        signal_4640), .Q(ciphertext_s0[41]), .QN() );
  DFF_X1 cell_330_s_reg_1_s_current_state_reg ( .D(signal_3867), .CK(
        signal_4640), .Q(ciphertext_s1[41]), .QN() );
  DFF_X1 cell_333_s_reg_0_s_current_state_reg ( .D(signal_629), .CK(
        signal_4640), .Q(ciphertext_s0[42]), .QN() );
  DFF_X1 cell_333_s_reg_1_s_current_state_reg ( .D(signal_3868), .CK(
        signal_4640), .Q(ciphertext_s1[42]), .QN() );
  DFF_X1 cell_336_s_reg_0_s_current_state_reg ( .D(signal_631), .CK(
        signal_4640), .Q(ciphertext_s0[43]), .QN() );
  DFF_X1 cell_336_s_reg_1_s_current_state_reg ( .D(signal_3869), .CK(
        signal_4640), .Q(ciphertext_s1[43]), .QN() );
  DFF_X1 cell_339_s_reg_0_s_current_state_reg ( .D(signal_633), .CK(
        signal_4640), .Q(ciphertext_s0[44]), .QN() );
  DFF_X1 cell_339_s_reg_1_s_current_state_reg ( .D(signal_3870), .CK(
        signal_4640), .Q(ciphertext_s1[44]), .QN() );
  DFF_X1 cell_342_s_reg_0_s_current_state_reg ( .D(signal_635), .CK(
        signal_4640), .Q(ciphertext_s0[45]), .QN() );
  DFF_X1 cell_342_s_reg_1_s_current_state_reg ( .D(signal_3871), .CK(
        signal_4640), .Q(ciphertext_s1[45]), .QN() );
  DFF_X1 cell_345_s_reg_0_s_current_state_reg ( .D(signal_637), .CK(
        signal_4640), .Q(ciphertext_s0[46]), .QN() );
  DFF_X1 cell_345_s_reg_1_s_current_state_reg ( .D(signal_3872), .CK(
        signal_4640), .Q(ciphertext_s1[46]), .QN() );
  DFF_X1 cell_348_s_reg_0_s_current_state_reg ( .D(signal_639), .CK(
        signal_4640), .Q(ciphertext_s0[47]), .QN() );
  DFF_X1 cell_348_s_reg_1_s_current_state_reg ( .D(signal_3873), .CK(
        signal_4640), .Q(ciphertext_s1[47]), .QN() );
  DFF_X1 cell_351_s_reg_0_s_current_state_reg ( .D(signal_641), .CK(
        signal_4640), .Q(ciphertext_s0[32]), .QN() );
  DFF_X1 cell_351_s_reg_1_s_current_state_reg ( .D(signal_3874), .CK(
        signal_4640), .Q(ciphertext_s1[32]), .QN() );
  DFF_X1 cell_354_s_reg_0_s_current_state_reg ( .D(signal_643), .CK(
        signal_4640), .Q(ciphertext_s0[33]), .QN() );
  DFF_X1 cell_354_s_reg_1_s_current_state_reg ( .D(signal_3875), .CK(
        signal_4640), .Q(ciphertext_s1[33]), .QN() );
  DFF_X1 cell_357_s_reg_0_s_current_state_reg ( .D(signal_645), .CK(
        signal_4640), .Q(ciphertext_s0[34]), .QN() );
  DFF_X1 cell_357_s_reg_1_s_current_state_reg ( .D(signal_3876), .CK(
        signal_4640), .Q(ciphertext_s1[34]), .QN() );
  DFF_X1 cell_360_s_reg_0_s_current_state_reg ( .D(signal_647), .CK(
        signal_4640), .Q(ciphertext_s0[35]), .QN() );
  DFF_X1 cell_360_s_reg_1_s_current_state_reg ( .D(signal_3877), .CK(
        signal_4640), .Q(ciphertext_s1[35]), .QN() );
  DFF_X1 cell_363_s_reg_0_s_current_state_reg ( .D(signal_649), .CK(
        signal_4640), .Q(ciphertext_s0[36]), .QN() );
  DFF_X1 cell_363_s_reg_1_s_current_state_reg ( .D(signal_3878), .CK(
        signal_4640), .Q(ciphertext_s1[36]), .QN() );
  DFF_X1 cell_366_s_reg_0_s_current_state_reg ( .D(signal_651), .CK(
        signal_4640), .Q(ciphertext_s0[37]), .QN() );
  DFF_X1 cell_366_s_reg_1_s_current_state_reg ( .D(signal_3879), .CK(
        signal_4640), .Q(ciphertext_s1[37]), .QN() );
  DFF_X1 cell_369_s_reg_0_s_current_state_reg ( .D(signal_653), .CK(
        signal_4640), .Q(ciphertext_s0[38]), .QN() );
  DFF_X1 cell_369_s_reg_1_s_current_state_reg ( .D(signal_3880), .CK(
        signal_4640), .Q(ciphertext_s1[38]), .QN() );
  DFF_X1 cell_372_s_reg_0_s_current_state_reg ( .D(signal_655), .CK(
        signal_4640), .Q(ciphertext_s0[39]), .QN() );
  DFF_X1 cell_372_s_reg_1_s_current_state_reg ( .D(signal_3881), .CK(
        signal_4640), .Q(ciphertext_s1[39]), .QN() );
  DFF_X1 cell_375_s_reg_0_s_current_state_reg ( .D(signal_657), .CK(
        signal_4640), .Q(ciphertext_s0[24]), .QN() );
  DFF_X1 cell_375_s_reg_1_s_current_state_reg ( .D(signal_3882), .CK(
        signal_4640), .Q(ciphertext_s1[24]), .QN() );
  DFF_X1 cell_378_s_reg_0_s_current_state_reg ( .D(signal_659), .CK(
        signal_4640), .Q(ciphertext_s0[25]), .QN() );
  DFF_X1 cell_378_s_reg_1_s_current_state_reg ( .D(signal_3883), .CK(
        signal_4640), .Q(ciphertext_s1[25]), .QN() );
  DFF_X1 cell_381_s_reg_0_s_current_state_reg ( .D(signal_661), .CK(
        signal_4640), .Q(ciphertext_s0[26]), .QN() );
  DFF_X1 cell_381_s_reg_1_s_current_state_reg ( .D(signal_3884), .CK(
        signal_4640), .Q(ciphertext_s1[26]), .QN() );
  DFF_X1 cell_384_s_reg_0_s_current_state_reg ( .D(signal_663), .CK(
        signal_4640), .Q(ciphertext_s0[27]), .QN() );
  DFF_X1 cell_384_s_reg_1_s_current_state_reg ( .D(signal_3885), .CK(
        signal_4640), .Q(ciphertext_s1[27]), .QN() );
  DFF_X1 cell_387_s_reg_0_s_current_state_reg ( .D(signal_665), .CK(
        signal_4640), .Q(ciphertext_s0[28]), .QN() );
  DFF_X1 cell_387_s_reg_1_s_current_state_reg ( .D(signal_3886), .CK(
        signal_4640), .Q(ciphertext_s1[28]), .QN() );
  DFF_X1 cell_390_s_reg_0_s_current_state_reg ( .D(signal_667), .CK(
        signal_4640), .Q(ciphertext_s0[29]), .QN() );
  DFF_X1 cell_390_s_reg_1_s_current_state_reg ( .D(signal_3887), .CK(
        signal_4640), .Q(ciphertext_s1[29]), .QN() );
  DFF_X1 cell_393_s_reg_0_s_current_state_reg ( .D(signal_669), .CK(
        signal_4640), .Q(ciphertext_s0[30]), .QN() );
  DFF_X1 cell_393_s_reg_1_s_current_state_reg ( .D(signal_3888), .CK(
        signal_4640), .Q(ciphertext_s1[30]), .QN() );
  DFF_X1 cell_396_s_reg_0_s_current_state_reg ( .D(signal_671), .CK(
        signal_4640), .Q(ciphertext_s0[31]), .QN() );
  DFF_X1 cell_396_s_reg_1_s_current_state_reg ( .D(signal_3889), .CK(
        signal_4640), .Q(ciphertext_s1[31]), .QN() );
  DFF_X1 cell_399_s_reg_0_s_current_state_reg ( .D(signal_673), .CK(
        signal_4640), .Q(ciphertext_s0[16]), .QN() );
  DFF_X1 cell_399_s_reg_1_s_current_state_reg ( .D(signal_3890), .CK(
        signal_4640), .Q(ciphertext_s1[16]), .QN() );
  DFF_X1 cell_402_s_reg_0_s_current_state_reg ( .D(signal_675), .CK(
        signal_4640), .Q(ciphertext_s0[17]), .QN() );
  DFF_X1 cell_402_s_reg_1_s_current_state_reg ( .D(signal_3891), .CK(
        signal_4640), .Q(ciphertext_s1[17]), .QN() );
  DFF_X1 cell_405_s_reg_0_s_current_state_reg ( .D(signal_677), .CK(
        signal_4640), .Q(ciphertext_s0[18]), .QN() );
  DFF_X1 cell_405_s_reg_1_s_current_state_reg ( .D(signal_3892), .CK(
        signal_4640), .Q(ciphertext_s1[18]), .QN() );
  DFF_X1 cell_408_s_reg_0_s_current_state_reg ( .D(signal_679), .CK(
        signal_4640), .Q(ciphertext_s0[19]), .QN() );
  DFF_X1 cell_408_s_reg_1_s_current_state_reg ( .D(signal_3893), .CK(
        signal_4640), .Q(ciphertext_s1[19]), .QN() );
  DFF_X1 cell_411_s_reg_0_s_current_state_reg ( .D(signal_681), .CK(
        signal_4640), .Q(ciphertext_s0[20]), .QN() );
  DFF_X1 cell_411_s_reg_1_s_current_state_reg ( .D(signal_3894), .CK(
        signal_4640), .Q(ciphertext_s1[20]), .QN() );
  DFF_X1 cell_414_s_reg_0_s_current_state_reg ( .D(signal_683), .CK(
        signal_4640), .Q(ciphertext_s0[21]), .QN() );
  DFF_X1 cell_414_s_reg_1_s_current_state_reg ( .D(signal_3895), .CK(
        signal_4640), .Q(ciphertext_s1[21]), .QN() );
  DFF_X1 cell_417_s_reg_0_s_current_state_reg ( .D(signal_685), .CK(
        signal_4640), .Q(ciphertext_s0[22]), .QN() );
  DFF_X1 cell_417_s_reg_1_s_current_state_reg ( .D(signal_3896), .CK(
        signal_4640), .Q(ciphertext_s1[22]), .QN() );
  DFF_X1 cell_420_s_reg_0_s_current_state_reg ( .D(signal_687), .CK(
        signal_4640), .Q(ciphertext_s0[23]), .QN() );
  DFF_X1 cell_420_s_reg_1_s_current_state_reg ( .D(signal_3897), .CK(
        signal_4640), .Q(ciphertext_s1[23]), .QN() );
  DFF_X1 cell_423_s_reg_0_s_current_state_reg ( .D(signal_689), .CK(
        signal_4640), .Q(ciphertext_s0[8]), .QN() );
  DFF_X1 cell_423_s_reg_1_s_current_state_reg ( .D(signal_3898), .CK(
        signal_4640), .Q(ciphertext_s1[8]), .QN() );
  DFF_X1 cell_426_s_reg_0_s_current_state_reg ( .D(signal_691), .CK(
        signal_4640), .Q(ciphertext_s0[9]), .QN() );
  DFF_X1 cell_426_s_reg_1_s_current_state_reg ( .D(signal_3899), .CK(
        signal_4640), .Q(ciphertext_s1[9]), .QN() );
  DFF_X1 cell_429_s_reg_0_s_current_state_reg ( .D(signal_693), .CK(
        signal_4640), .Q(ciphertext_s0[10]), .QN() );
  DFF_X1 cell_429_s_reg_1_s_current_state_reg ( .D(signal_3900), .CK(
        signal_4640), .Q(ciphertext_s1[10]), .QN() );
  DFF_X1 cell_432_s_reg_0_s_current_state_reg ( .D(signal_695), .CK(
        signal_4640), .Q(ciphertext_s0[11]), .QN() );
  DFF_X1 cell_432_s_reg_1_s_current_state_reg ( .D(signal_3901), .CK(
        signal_4640), .Q(ciphertext_s1[11]), .QN() );
  DFF_X1 cell_435_s_reg_0_s_current_state_reg ( .D(signal_697), .CK(
        signal_4640), .Q(ciphertext_s0[12]), .QN() );
  DFF_X1 cell_435_s_reg_1_s_current_state_reg ( .D(signal_3902), .CK(
        signal_4640), .Q(ciphertext_s1[12]), .QN() );
  DFF_X1 cell_438_s_reg_0_s_current_state_reg ( .D(signal_699), .CK(
        signal_4640), .Q(ciphertext_s0[13]), .QN() );
  DFF_X1 cell_438_s_reg_1_s_current_state_reg ( .D(signal_3903), .CK(
        signal_4640), .Q(ciphertext_s1[13]), .QN() );
  DFF_X1 cell_441_s_reg_0_s_current_state_reg ( .D(signal_701), .CK(
        signal_4640), .Q(ciphertext_s0[14]), .QN() );
  DFF_X1 cell_441_s_reg_1_s_current_state_reg ( .D(signal_3904), .CK(
        signal_4640), .Q(ciphertext_s1[14]), .QN() );
  DFF_X1 cell_444_s_reg_0_s_current_state_reg ( .D(signal_703), .CK(
        signal_4640), .Q(ciphertext_s0[15]), .QN() );
  DFF_X1 cell_444_s_reg_1_s_current_state_reg ( .D(signal_3905), .CK(
        signal_4640), .Q(ciphertext_s1[15]), .QN() );
  DFF_X1 cell_447_s_reg_0_s_current_state_reg ( .D(signal_705), .CK(
        signal_4640), .Q(ciphertext_s0[0]), .QN() );
  DFF_X1 cell_447_s_reg_1_s_current_state_reg ( .D(signal_4210), .CK(
        signal_4640), .Q(ciphertext_s1[0]), .QN() );
  DFF_X1 cell_450_s_reg_0_s_current_state_reg ( .D(signal_707), .CK(
        signal_4640), .Q(ciphertext_s0[1]), .QN() );
  DFF_X1 cell_450_s_reg_1_s_current_state_reg ( .D(signal_4211), .CK(
        signal_4640), .Q(ciphertext_s1[1]), .QN() );
  DFF_X1 cell_453_s_reg_0_s_current_state_reg ( .D(signal_709), .CK(
        signal_4640), .Q(ciphertext_s0[2]), .QN() );
  DFF_X1 cell_453_s_reg_1_s_current_state_reg ( .D(signal_4212), .CK(
        signal_4640), .Q(ciphertext_s1[2]), .QN() );
  DFF_X1 cell_456_s_reg_0_s_current_state_reg ( .D(signal_711), .CK(
        signal_4640), .Q(ciphertext_s0[3]), .QN() );
  DFF_X1 cell_456_s_reg_1_s_current_state_reg ( .D(signal_4213), .CK(
        signal_4640), .Q(ciphertext_s1[3]), .QN() );
  DFF_X1 cell_459_s_reg_0_s_current_state_reg ( .D(signal_713), .CK(
        signal_4640), .Q(ciphertext_s0[4]), .QN() );
  DFF_X1 cell_459_s_reg_1_s_current_state_reg ( .D(signal_4214), .CK(
        signal_4640), .Q(ciphertext_s1[4]), .QN() );
  DFF_X1 cell_462_s_reg_0_s_current_state_reg ( .D(signal_715), .CK(
        signal_4640), .Q(ciphertext_s0[5]), .QN() );
  DFF_X1 cell_462_s_reg_1_s_current_state_reg ( .D(signal_4215), .CK(
        signal_4640), .Q(ciphertext_s1[5]), .QN() );
  DFF_X1 cell_465_s_reg_0_s_current_state_reg ( .D(signal_717), .CK(
        signal_4640), .Q(ciphertext_s0[6]), .QN() );
  DFF_X1 cell_465_s_reg_1_s_current_state_reg ( .D(signal_4216), .CK(
        signal_4640), .Q(ciphertext_s1[6]), .QN() );
  DFF_X1 cell_468_s_reg_0_s_current_state_reg ( .D(signal_719), .CK(
        signal_4640), .Q(ciphertext_s0[7]), .QN() );
  DFF_X1 cell_468_s_reg_1_s_current_state_reg ( .D(signal_4217), .CK(
        signal_4640), .Q(ciphertext_s1[7]), .QN() );
  DFF_X1 cell_717_s_reg_0_s_current_state_reg ( .D(signal_766), .CK(
        signal_4640), .Q(signal_1493), .QN() );
  DFF_X1 cell_717_s_reg_1_s_current_state_reg ( .D(signal_4122), .CK(
        signal_4640), .Q(signal_2389), .QN() );
  DFF_X1 cell_721_s_reg_0_s_current_state_reg ( .D(signal_769), .CK(
        signal_4640), .Q(signal_1492), .QN() );
  DFF_X1 cell_721_s_reg_1_s_current_state_reg ( .D(signal_4123), .CK(
        signal_4640), .Q(signal_2392), .QN() );
  DFF_X1 cell_725_s_reg_0_s_current_state_reg ( .D(signal_772), .CK(
        signal_4640), .Q(signal_1491), .QN() );
  DFF_X1 cell_725_s_reg_1_s_current_state_reg ( .D(signal_4124), .CK(
        signal_4640), .Q(signal_2395), .QN() );
  DFF_X1 cell_729_s_reg_0_s_current_state_reg ( .D(signal_775), .CK(
        signal_4640), .Q(signal_1490), .QN() );
  DFF_X1 cell_729_s_reg_1_s_current_state_reg ( .D(signal_4125), .CK(
        signal_4640), .Q(signal_2398), .QN() );
  DFF_X1 cell_733_s_reg_0_s_current_state_reg ( .D(signal_778), .CK(
        signal_4640), .Q(signal_1489), .QN() );
  DFF_X1 cell_733_s_reg_1_s_current_state_reg ( .D(signal_4126), .CK(
        signal_4640), .Q(signal_2401), .QN() );
  DFF_X1 cell_737_s_reg_0_s_current_state_reg ( .D(signal_781), .CK(
        signal_4640), .Q(signal_1488), .QN() );
  DFF_X1 cell_737_s_reg_1_s_current_state_reg ( .D(signal_4127), .CK(
        signal_4640), .Q(signal_2404), .QN() );
  DFF_X1 cell_741_s_reg_0_s_current_state_reg ( .D(signal_784), .CK(
        signal_4640), .Q(signal_1487), .QN() );
  DFF_X1 cell_741_s_reg_1_s_current_state_reg ( .D(signal_4128), .CK(
        signal_4640), .Q(signal_2407), .QN() );
  DFF_X1 cell_745_s_reg_0_s_current_state_reg ( .D(signal_787), .CK(
        signal_4640), .Q(signal_1486), .QN() );
  DFF_X1 cell_745_s_reg_1_s_current_state_reg ( .D(signal_4129), .CK(
        signal_4640), .Q(signal_2410), .QN() );
  DFF_X1 cell_749_s_reg_0_s_current_state_reg ( .D(signal_790), .CK(
        signal_4640), .Q(signal_758), .QN() );
  DFF_X1 cell_749_s_reg_1_s_current_state_reg ( .D(signal_3994), .CK(
        signal_4640), .Q(signal_2426), .QN() );
  DFF_X1 cell_753_s_reg_0_s_current_state_reg ( .D(signal_793), .CK(
        signal_4640), .Q(signal_759), .QN() );
  DFF_X1 cell_753_s_reg_1_s_current_state_reg ( .D(signal_3995), .CK(
        signal_4640), .Q(signal_2424), .QN() );
  DFF_X1 cell_757_s_reg_0_s_current_state_reg ( .D(signal_796), .CK(
        signal_4640), .Q(signal_760), .QN() );
  DFF_X1 cell_757_s_reg_1_s_current_state_reg ( .D(signal_3996), .CK(
        signal_4640), .Q(signal_2422), .QN() );
  DFF_X1 cell_761_s_reg_0_s_current_state_reg ( .D(signal_799), .CK(
        signal_4640), .Q(signal_761), .QN() );
  DFF_X1 cell_761_s_reg_1_s_current_state_reg ( .D(signal_3997), .CK(
        signal_4640), .Q(signal_2420), .QN() );
  DFF_X1 cell_765_s_reg_0_s_current_state_reg ( .D(signal_802), .CK(
        signal_4640), .Q(signal_762), .QN() );
  DFF_X1 cell_765_s_reg_1_s_current_state_reg ( .D(signal_3998), .CK(
        signal_4640), .Q(signal_2418), .QN() );
  DFF_X1 cell_769_s_reg_0_s_current_state_reg ( .D(signal_805), .CK(
        signal_4640), .Q(signal_763), .QN() );
  DFF_X1 cell_769_s_reg_1_s_current_state_reg ( .D(signal_3999), .CK(
        signal_4640), .Q(signal_2416), .QN() );
  DFF_X1 cell_773_s_reg_0_s_current_state_reg ( .D(signal_808), .CK(
        signal_4640), .Q(signal_764), .QN() );
  DFF_X1 cell_773_s_reg_1_s_current_state_reg ( .D(signal_4000), .CK(
        signal_4640), .Q(signal_2414), .QN() );
  DFF_X1 cell_777_s_reg_0_s_current_state_reg ( .D(signal_811), .CK(
        signal_4640), .Q(signal_765), .QN() );
  DFF_X1 cell_777_s_reg_1_s_current_state_reg ( .D(signal_4001), .CK(
        signal_4640), .Q(signal_2412), .QN() );
  DFF_X1 cell_781_s_reg_0_s_current_state_reg ( .D(signal_814), .CK(
        signal_4640), .Q(signal_1909), .QN() );
  DFF_X1 cell_781_s_reg_1_s_current_state_reg ( .D(signal_4002), .CK(
        signal_4640), .Q(signal_2849), .QN() );
  DFF_X1 cell_785_s_reg_0_s_current_state_reg ( .D(signal_817), .CK(
        signal_4640), .Q(signal_1908), .QN() );
  DFF_X1 cell_785_s_reg_1_s_current_state_reg ( .D(signal_4003), .CK(
        signal_4640), .Q(signal_2852), .QN() );
  DFF_X1 cell_789_s_reg_0_s_current_state_reg ( .D(signal_820), .CK(
        signal_4640), .Q(signal_1907), .QN() );
  DFF_X1 cell_789_s_reg_1_s_current_state_reg ( .D(signal_4004), .CK(
        signal_4640), .Q(signal_2855), .QN() );
  DFF_X1 cell_793_s_reg_0_s_current_state_reg ( .D(signal_823), .CK(
        signal_4640), .Q(signal_1906), .QN() );
  DFF_X1 cell_793_s_reg_1_s_current_state_reg ( .D(signal_4005), .CK(
        signal_4640), .Q(signal_2858), .QN() );
  DFF_X1 cell_797_s_reg_0_s_current_state_reg ( .D(signal_826), .CK(
        signal_4640), .Q(signal_1905), .QN() );
  DFF_X1 cell_797_s_reg_1_s_current_state_reg ( .D(signal_4006), .CK(
        signal_4640), .Q(signal_2861), .QN() );
  DFF_X1 cell_801_s_reg_0_s_current_state_reg ( .D(signal_829), .CK(
        signal_4640), .Q(signal_1904), .QN() );
  DFF_X1 cell_801_s_reg_1_s_current_state_reg ( .D(signal_4007), .CK(
        signal_4640), .Q(signal_2864), .QN() );
  DFF_X1 cell_805_s_reg_0_s_current_state_reg ( .D(signal_832), .CK(
        signal_4640), .Q(signal_1903), .QN() );
  DFF_X1 cell_805_s_reg_1_s_current_state_reg ( .D(signal_4008), .CK(
        signal_4640), .Q(signal_2867), .QN() );
  DFF_X1 cell_809_s_reg_0_s_current_state_reg ( .D(signal_835), .CK(
        signal_4640), .Q(signal_1902), .QN() );
  DFF_X1 cell_809_s_reg_1_s_current_state_reg ( .D(signal_4009), .CK(
        signal_4640), .Q(signal_2870), .QN() );
  DFF_X1 cell_813_s_reg_0_s_current_state_reg ( .D(signal_838), .CK(
        signal_4640), .Q(signal_1893), .QN() );
  DFF_X1 cell_813_s_reg_1_s_current_state_reg ( .D(signal_4010), .CK(
        signal_4640), .Q(signal_2873), .QN() );
  DFF_X1 cell_817_s_reg_0_s_current_state_reg ( .D(signal_841), .CK(
        signal_4640), .Q(signal_1892), .QN() );
  DFF_X1 cell_817_s_reg_1_s_current_state_reg ( .D(signal_4011), .CK(
        signal_4640), .Q(signal_2876), .QN() );
  DFF_X1 cell_821_s_reg_0_s_current_state_reg ( .D(signal_844), .CK(
        signal_4640), .Q(signal_1891), .QN() );
  DFF_X1 cell_821_s_reg_1_s_current_state_reg ( .D(signal_4012), .CK(
        signal_4640), .Q(signal_2879), .QN() );
  DFF_X1 cell_825_s_reg_0_s_current_state_reg ( .D(signal_847), .CK(
        signal_4640), .Q(signal_1890), .QN() );
  DFF_X1 cell_825_s_reg_1_s_current_state_reg ( .D(signal_4013), .CK(
        signal_4640), .Q(signal_2882), .QN() );
  DFF_X1 cell_829_s_reg_0_s_current_state_reg ( .D(signal_850), .CK(
        signal_4640), .Q(signal_1889), .QN() );
  DFF_X1 cell_829_s_reg_1_s_current_state_reg ( .D(signal_4014), .CK(
        signal_4640), .Q(signal_2885), .QN() );
  DFF_X1 cell_833_s_reg_0_s_current_state_reg ( .D(signal_853), .CK(
        signal_4640), .Q(signal_1888), .QN() );
  DFF_X1 cell_833_s_reg_1_s_current_state_reg ( .D(signal_4015), .CK(
        signal_4640), .Q(signal_2888), .QN() );
  DFF_X1 cell_837_s_reg_0_s_current_state_reg ( .D(signal_856), .CK(
        signal_4640), .Q(signal_1887), .QN() );
  DFF_X1 cell_837_s_reg_1_s_current_state_reg ( .D(signal_4016), .CK(
        signal_4640), .Q(signal_2891), .QN() );
  DFF_X1 cell_841_s_reg_0_s_current_state_reg ( .D(signal_859), .CK(
        signal_4640), .Q(signal_1886), .QN() );
  DFF_X1 cell_841_s_reg_1_s_current_state_reg ( .D(signal_4017), .CK(
        signal_4640), .Q(signal_2894), .QN() );
  DFF_X1 cell_845_s_reg_0_s_current_state_reg ( .D(signal_862), .CK(
        signal_4640), .Q(signal_1877), .QN() );
  DFF_X1 cell_845_s_reg_1_s_current_state_reg ( .D(signal_4018), .CK(
        signal_4640), .Q(signal_2897), .QN() );
  DFF_X1 cell_849_s_reg_0_s_current_state_reg ( .D(signal_865), .CK(
        signal_4640), .Q(signal_1876), .QN() );
  DFF_X1 cell_849_s_reg_1_s_current_state_reg ( .D(signal_4019), .CK(
        signal_4640), .Q(signal_2900), .QN() );
  DFF_X1 cell_853_s_reg_0_s_current_state_reg ( .D(signal_868), .CK(
        signal_4640), .Q(signal_1875), .QN() );
  DFF_X1 cell_853_s_reg_1_s_current_state_reg ( .D(signal_4020), .CK(
        signal_4640), .Q(signal_2903), .QN() );
  DFF_X1 cell_857_s_reg_0_s_current_state_reg ( .D(signal_871), .CK(
        signal_4640), .Q(signal_1874), .QN() );
  DFF_X1 cell_857_s_reg_1_s_current_state_reg ( .D(signal_4021), .CK(
        signal_4640), .Q(signal_2906), .QN() );
  DFF_X1 cell_861_s_reg_0_s_current_state_reg ( .D(signal_874), .CK(
        signal_4640), .Q(signal_1873), .QN() );
  DFF_X1 cell_861_s_reg_1_s_current_state_reg ( .D(signal_4022), .CK(
        signal_4640), .Q(signal_2909), .QN() );
  DFF_X1 cell_865_s_reg_0_s_current_state_reg ( .D(signal_877), .CK(
        signal_4640), .Q(signal_1872), .QN() );
  DFF_X1 cell_865_s_reg_1_s_current_state_reg ( .D(signal_4023), .CK(
        signal_4640), .Q(signal_2912), .QN() );
  DFF_X1 cell_869_s_reg_0_s_current_state_reg ( .D(signal_880), .CK(
        signal_4640), .Q(signal_1871), .QN() );
  DFF_X1 cell_869_s_reg_1_s_current_state_reg ( .D(signal_4024), .CK(
        signal_4640), .Q(signal_2915), .QN() );
  DFF_X1 cell_873_s_reg_0_s_current_state_reg ( .D(signal_883), .CK(
        signal_4640), .Q(signal_1870), .QN() );
  DFF_X1 cell_873_s_reg_1_s_current_state_reg ( .D(signal_4025), .CK(
        signal_4640), .Q(signal_2918), .QN() );
  DFF_X1 cell_877_s_reg_0_s_current_state_reg ( .D(signal_886), .CK(
        signal_4640), .Q(signal_1861), .QN() );
  DFF_X1 cell_877_s_reg_1_s_current_state_reg ( .D(signal_4026), .CK(
        signal_4640), .Q(signal_2921), .QN() );
  DFF_X1 cell_881_s_reg_0_s_current_state_reg ( .D(signal_889), .CK(
        signal_4640), .Q(signal_1860), .QN() );
  DFF_X1 cell_881_s_reg_1_s_current_state_reg ( .D(signal_4027), .CK(
        signal_4640), .Q(signal_2924), .QN() );
  DFF_X1 cell_885_s_reg_0_s_current_state_reg ( .D(signal_892), .CK(
        signal_4640), .Q(signal_1859), .QN() );
  DFF_X1 cell_885_s_reg_1_s_current_state_reg ( .D(signal_4028), .CK(
        signal_4640), .Q(signal_2927), .QN() );
  DFF_X1 cell_889_s_reg_0_s_current_state_reg ( .D(signal_895), .CK(
        signal_4640), .Q(signal_1858), .QN() );
  DFF_X1 cell_889_s_reg_1_s_current_state_reg ( .D(signal_4029), .CK(
        signal_4640), .Q(signal_2930), .QN() );
  DFF_X1 cell_893_s_reg_0_s_current_state_reg ( .D(signal_898), .CK(
        signal_4640), .Q(signal_1857), .QN() );
  DFF_X1 cell_893_s_reg_1_s_current_state_reg ( .D(signal_4030), .CK(
        signal_4640), .Q(signal_2933), .QN() );
  DFF_X1 cell_897_s_reg_0_s_current_state_reg ( .D(signal_901), .CK(
        signal_4640), .Q(signal_1856), .QN() );
  DFF_X1 cell_897_s_reg_1_s_current_state_reg ( .D(signal_4031), .CK(
        signal_4640), .Q(signal_2936), .QN() );
  DFF_X1 cell_901_s_reg_0_s_current_state_reg ( .D(signal_904), .CK(
        signal_4640), .Q(signal_1855), .QN() );
  DFF_X1 cell_901_s_reg_1_s_current_state_reg ( .D(signal_4032), .CK(
        signal_4640), .Q(signal_2939), .QN() );
  DFF_X1 cell_905_s_reg_0_s_current_state_reg ( .D(signal_907), .CK(
        signal_4640), .Q(signal_1854), .QN() );
  DFF_X1 cell_905_s_reg_1_s_current_state_reg ( .D(signal_4033), .CK(
        signal_4640), .Q(signal_2942), .QN() );
  DFF_X1 cell_909_s_reg_0_s_current_state_reg ( .D(signal_910), .CK(
        signal_4640), .Q(signal_1845), .QN() );
  DFF_X1 cell_909_s_reg_1_s_current_state_reg ( .D(signal_3639), .CK(
        signal_4640), .Q(signal_2945), .QN() );
  DFF_X1 cell_913_s_reg_0_s_current_state_reg ( .D(signal_913), .CK(
        signal_4640), .Q(signal_1844), .QN() );
  DFF_X1 cell_913_s_reg_1_s_current_state_reg ( .D(signal_3640), .CK(
        signal_4640), .Q(signal_2948), .QN() );
  DFF_X1 cell_917_s_reg_0_s_current_state_reg ( .D(signal_916), .CK(
        signal_4640), .Q(signal_1843), .QN() );
  DFF_X1 cell_917_s_reg_1_s_current_state_reg ( .D(signal_3641), .CK(
        signal_4640), .Q(signal_2951), .QN() );
  DFF_X1 cell_921_s_reg_0_s_current_state_reg ( .D(signal_919), .CK(
        signal_4640), .Q(signal_1842), .QN() );
  DFF_X1 cell_921_s_reg_1_s_current_state_reg ( .D(signal_3642), .CK(
        signal_4640), .Q(signal_2954), .QN() );
  DFF_X1 cell_925_s_reg_0_s_current_state_reg ( .D(signal_922), .CK(
        signal_4640), .Q(signal_1841), .QN() );
  DFF_X1 cell_925_s_reg_1_s_current_state_reg ( .D(signal_3643), .CK(
        signal_4640), .Q(signal_2957), .QN() );
  DFF_X1 cell_929_s_reg_0_s_current_state_reg ( .D(signal_925), .CK(
        signal_4640), .Q(signal_1840), .QN() );
  DFF_X1 cell_929_s_reg_1_s_current_state_reg ( .D(signal_3644), .CK(
        signal_4640), .Q(signal_2960), .QN() );
  DFF_X1 cell_933_s_reg_0_s_current_state_reg ( .D(signal_928), .CK(
        signal_4640), .Q(signal_1839), .QN() );
  DFF_X1 cell_933_s_reg_1_s_current_state_reg ( .D(signal_3645), .CK(
        signal_4640), .Q(signal_2963), .QN() );
  DFF_X1 cell_937_s_reg_0_s_current_state_reg ( .D(signal_931), .CK(
        signal_4640), .Q(signal_1838), .QN() );
  DFF_X1 cell_937_s_reg_1_s_current_state_reg ( .D(signal_3646), .CK(
        signal_4640), .Q(signal_2966), .QN() );
  DFF_X1 cell_941_s_reg_0_s_current_state_reg ( .D(signal_934), .CK(
        signal_4640), .Q(signal_1509), .QN() );
  DFF_X1 cell_941_s_reg_1_s_current_state_reg ( .D(signal_3647), .CK(
        signal_4640), .Q(signal_2969), .QN() );
  DFF_X1 cell_945_s_reg_0_s_current_state_reg ( .D(signal_937), .CK(
        signal_4640), .Q(signal_1508), .QN() );
  DFF_X1 cell_945_s_reg_1_s_current_state_reg ( .D(signal_3648), .CK(
        signal_4640), .Q(signal_2972), .QN() );
  DFF_X1 cell_949_s_reg_0_s_current_state_reg ( .D(signal_940), .CK(
        signal_4640), .Q(signal_1507), .QN() );
  DFF_X1 cell_949_s_reg_1_s_current_state_reg ( .D(signal_3649), .CK(
        signal_4640), .Q(signal_2975), .QN() );
  DFF_X1 cell_953_s_reg_0_s_current_state_reg ( .D(signal_943), .CK(
        signal_4640), .Q(signal_1506), .QN() );
  DFF_X1 cell_953_s_reg_1_s_current_state_reg ( .D(signal_3650), .CK(
        signal_4640), .Q(signal_2978), .QN() );
  DFF_X1 cell_957_s_reg_0_s_current_state_reg ( .D(signal_946), .CK(
        signal_4640), .Q(signal_1505), .QN() );
  DFF_X1 cell_957_s_reg_1_s_current_state_reg ( .D(signal_3651), .CK(
        signal_4640), .Q(signal_2981), .QN() );
  DFF_X1 cell_961_s_reg_0_s_current_state_reg ( .D(signal_949), .CK(
        signal_4640), .Q(signal_1504), .QN() );
  DFF_X1 cell_961_s_reg_1_s_current_state_reg ( .D(signal_3652), .CK(
        signal_4640), .Q(signal_2984), .QN() );
  DFF_X1 cell_965_s_reg_0_s_current_state_reg ( .D(signal_952), .CK(
        signal_4640), .Q(signal_1503), .QN() );
  DFF_X1 cell_965_s_reg_1_s_current_state_reg ( .D(signal_3653), .CK(
        signal_4640), .Q(signal_2987), .QN() );
  DFF_X1 cell_969_s_reg_0_s_current_state_reg ( .D(signal_955), .CK(
        signal_4640), .Q(signal_1502), .QN() );
  DFF_X1 cell_969_s_reg_1_s_current_state_reg ( .D(signal_3654), .CK(
        signal_4640), .Q(signal_2990), .QN() );
  DFF_X1 cell_973_s_reg_0_s_current_state_reg ( .D(signal_958), .CK(
        signal_4640), .Q(signal_1821), .QN() );
  DFF_X1 cell_973_s_reg_1_s_current_state_reg ( .D(signal_4034), .CK(
        signal_4640), .Q(signal_2993), .QN() );
  DFF_X1 cell_977_s_reg_0_s_current_state_reg ( .D(signal_961), .CK(
        signal_4640), .Q(signal_1820), .QN() );
  DFF_X1 cell_977_s_reg_1_s_current_state_reg ( .D(signal_4035), .CK(
        signal_4640), .Q(signal_2996), .QN() );
  DFF_X1 cell_981_s_reg_0_s_current_state_reg ( .D(signal_964), .CK(
        signal_4640), .Q(signal_1819), .QN() );
  DFF_X1 cell_981_s_reg_1_s_current_state_reg ( .D(signal_4036), .CK(
        signal_4640), .Q(signal_2999), .QN() );
  DFF_X1 cell_985_s_reg_0_s_current_state_reg ( .D(signal_967), .CK(
        signal_4640), .Q(signal_1818), .QN() );
  DFF_X1 cell_985_s_reg_1_s_current_state_reg ( .D(signal_4037), .CK(
        signal_4640), .Q(signal_3002), .QN() );
  DFF_X1 cell_989_s_reg_0_s_current_state_reg ( .D(signal_970), .CK(
        signal_4640), .Q(signal_1817), .QN() );
  DFF_X1 cell_989_s_reg_1_s_current_state_reg ( .D(signal_4038), .CK(
        signal_4640), .Q(signal_3005), .QN() );
  DFF_X1 cell_993_s_reg_0_s_current_state_reg ( .D(signal_973), .CK(
        signal_4640), .Q(signal_1816), .QN() );
  DFF_X1 cell_993_s_reg_1_s_current_state_reg ( .D(signal_4039), .CK(
        signal_4640), .Q(signal_3008), .QN() );
  DFF_X1 cell_997_s_reg_0_s_current_state_reg ( .D(signal_976), .CK(
        signal_4640), .Q(signal_1815), .QN() );
  DFF_X1 cell_997_s_reg_1_s_current_state_reg ( .D(signal_4040), .CK(
        signal_4640), .Q(signal_3011), .QN() );
  DFF_X1 cell_1001_s_reg_0_s_current_state_reg ( .D(signal_979), .CK(
        signal_4640), .Q(signal_1814), .QN() );
  DFF_X1 cell_1001_s_reg_1_s_current_state_reg ( .D(signal_4041), .CK(
        signal_4640), .Q(signal_3014), .QN() );
  DFF_X1 cell_1005_s_reg_0_s_current_state_reg ( .D(signal_982), .CK(
        signal_4640), .Q(signal_1805), .QN() );
  DFF_X1 cell_1005_s_reg_1_s_current_state_reg ( .D(signal_4042), .CK(
        signal_4640), .Q(signal_3017), .QN() );
  DFF_X1 cell_1009_s_reg_0_s_current_state_reg ( .D(signal_985), .CK(
        signal_4640), .Q(signal_1804), .QN() );
  DFF_X1 cell_1009_s_reg_1_s_current_state_reg ( .D(signal_4043), .CK(
        signal_4640), .Q(signal_3020), .QN() );
  DFF_X1 cell_1013_s_reg_0_s_current_state_reg ( .D(signal_988), .CK(
        signal_4640), .Q(signal_1803), .QN() );
  DFF_X1 cell_1013_s_reg_1_s_current_state_reg ( .D(signal_4044), .CK(
        signal_4640), .Q(signal_3023), .QN() );
  DFF_X1 cell_1017_s_reg_0_s_current_state_reg ( .D(signal_991), .CK(
        signal_4640), .Q(signal_1802), .QN() );
  DFF_X1 cell_1017_s_reg_1_s_current_state_reg ( .D(signal_4045), .CK(
        signal_4640), .Q(signal_3026), .QN() );
  DFF_X1 cell_1021_s_reg_0_s_current_state_reg ( .D(signal_994), .CK(
        signal_4640), .Q(signal_1801), .QN() );
  DFF_X1 cell_1021_s_reg_1_s_current_state_reg ( .D(signal_4046), .CK(
        signal_4640), .Q(signal_3029), .QN() );
  DFF_X1 cell_1025_s_reg_0_s_current_state_reg ( .D(signal_997), .CK(
        signal_4640), .Q(signal_1800), .QN() );
  DFF_X1 cell_1025_s_reg_1_s_current_state_reg ( .D(signal_4047), .CK(
        signal_4640), .Q(signal_3032), .QN() );
  DFF_X1 cell_1029_s_reg_0_s_current_state_reg ( .D(signal_1000), .CK(
        signal_4640), .Q(signal_1799), .QN() );
  DFF_X1 cell_1029_s_reg_1_s_current_state_reg ( .D(signal_4048), .CK(
        signal_4640), .Q(signal_3035), .QN() );
  DFF_X1 cell_1033_s_reg_0_s_current_state_reg ( .D(signal_1003), .CK(
        signal_4640), .Q(signal_1798), .QN() );
  DFF_X1 cell_1033_s_reg_1_s_current_state_reg ( .D(signal_4049), .CK(
        signal_4640), .Q(signal_3038), .QN() );
  DFF_X1 cell_1037_s_reg_0_s_current_state_reg ( .D(signal_1006), .CK(
        signal_4640), .Q(signal_1789), .QN() );
  DFF_X1 cell_1037_s_reg_1_s_current_state_reg ( .D(signal_4050), .CK(
        signal_4640), .Q(signal_3041), .QN() );
  DFF_X1 cell_1041_s_reg_0_s_current_state_reg ( .D(signal_1009), .CK(
        signal_4640), .Q(signal_1788), .QN() );
  DFF_X1 cell_1041_s_reg_1_s_current_state_reg ( .D(signal_4051), .CK(
        signal_4640), .Q(signal_3044), .QN() );
  DFF_X1 cell_1045_s_reg_0_s_current_state_reg ( .D(signal_1012), .CK(
        signal_4640), .Q(signal_1787), .QN() );
  DFF_X1 cell_1045_s_reg_1_s_current_state_reg ( .D(signal_4052), .CK(
        signal_4640), .Q(signal_3047), .QN() );
  DFF_X1 cell_1049_s_reg_0_s_current_state_reg ( .D(signal_1015), .CK(
        signal_4640), .Q(signal_1786), .QN() );
  DFF_X1 cell_1049_s_reg_1_s_current_state_reg ( .D(signal_4053), .CK(
        signal_4640), .Q(signal_3050), .QN() );
  DFF_X1 cell_1053_s_reg_0_s_current_state_reg ( .D(signal_1018), .CK(
        signal_4640), .Q(signal_1785), .QN() );
  DFF_X1 cell_1053_s_reg_1_s_current_state_reg ( .D(signal_4054), .CK(
        signal_4640), .Q(signal_3053), .QN() );
  DFF_X1 cell_1057_s_reg_0_s_current_state_reg ( .D(signal_1021), .CK(
        signal_4640), .Q(signal_1784), .QN() );
  DFF_X1 cell_1057_s_reg_1_s_current_state_reg ( .D(signal_4055), .CK(
        signal_4640), .Q(signal_3056), .QN() );
  DFF_X1 cell_1061_s_reg_0_s_current_state_reg ( .D(signal_1024), .CK(
        signal_4640), .Q(signal_1783), .QN() );
  DFF_X1 cell_1061_s_reg_1_s_current_state_reg ( .D(signal_4056), .CK(
        signal_4640), .Q(signal_3059), .QN() );
  DFF_X1 cell_1065_s_reg_0_s_current_state_reg ( .D(signal_1027), .CK(
        signal_4640), .Q(signal_1782), .QN() );
  DFF_X1 cell_1065_s_reg_1_s_current_state_reg ( .D(signal_4057), .CK(
        signal_4640), .Q(signal_3062), .QN() );
  DFF_X1 cell_1069_s_reg_0_s_current_state_reg ( .D(signal_1030), .CK(
        signal_4640), .Q(signal_1773), .QN() );
  DFF_X1 cell_1069_s_reg_1_s_current_state_reg ( .D(signal_4058), .CK(
        signal_4640), .Q(signal_3065), .QN() );
  DFF_X1 cell_1073_s_reg_0_s_current_state_reg ( .D(signal_1033), .CK(
        signal_4640), .Q(signal_1772), .QN() );
  DFF_X1 cell_1073_s_reg_1_s_current_state_reg ( .D(signal_4059), .CK(
        signal_4640), .Q(signal_3068), .QN() );
  DFF_X1 cell_1077_s_reg_0_s_current_state_reg ( .D(signal_1036), .CK(
        signal_4640), .Q(signal_1771), .QN() );
  DFF_X1 cell_1077_s_reg_1_s_current_state_reg ( .D(signal_4060), .CK(
        signal_4640), .Q(signal_3071), .QN() );
  DFF_X1 cell_1081_s_reg_0_s_current_state_reg ( .D(signal_1039), .CK(
        signal_4640), .Q(signal_1770), .QN() );
  DFF_X1 cell_1081_s_reg_1_s_current_state_reg ( .D(signal_4061), .CK(
        signal_4640), .Q(signal_3074), .QN() );
  DFF_X1 cell_1085_s_reg_0_s_current_state_reg ( .D(signal_1042), .CK(
        signal_4640), .Q(signal_1769), .QN() );
  DFF_X1 cell_1085_s_reg_1_s_current_state_reg ( .D(signal_4062), .CK(
        signal_4640), .Q(signal_3077), .QN() );
  DFF_X1 cell_1089_s_reg_0_s_current_state_reg ( .D(signal_1045), .CK(
        signal_4640), .Q(signal_1768), .QN() );
  DFF_X1 cell_1089_s_reg_1_s_current_state_reg ( .D(signal_4063), .CK(
        signal_4640), .Q(signal_3080), .QN() );
  DFF_X1 cell_1093_s_reg_0_s_current_state_reg ( .D(signal_1048), .CK(
        signal_4640), .Q(signal_1767), .QN() );
  DFF_X1 cell_1093_s_reg_1_s_current_state_reg ( .D(signal_4064), .CK(
        signal_4640), .Q(signal_3083), .QN() );
  DFF_X1 cell_1097_s_reg_0_s_current_state_reg ( .D(signal_1051), .CK(
        signal_4640), .Q(signal_1766), .QN() );
  DFF_X1 cell_1097_s_reg_1_s_current_state_reg ( .D(signal_4065), .CK(
        signal_4640), .Q(signal_3086), .QN() );
  DFF_X1 cell_1101_s_reg_0_s_current_state_reg ( .D(signal_1054), .CK(
        signal_4640), .Q(signal_1749), .QN() );
  DFF_X1 cell_1101_s_reg_1_s_current_state_reg ( .D(signal_4218), .CK(
        signal_4640), .Q(signal_3089), .QN() );
  DFF_X1 cell_1105_s_reg_0_s_current_state_reg ( .D(signal_1057), .CK(
        signal_4640), .Q(signal_1748), .QN() );
  DFF_X1 cell_1105_s_reg_1_s_current_state_reg ( .D(signal_4219), .CK(
        signal_4640), .Q(signal_3092), .QN() );
  DFF_X1 cell_1109_s_reg_0_s_current_state_reg ( .D(signal_1060), .CK(
        signal_4640), .Q(signal_1747), .QN() );
  DFF_X1 cell_1109_s_reg_1_s_current_state_reg ( .D(signal_4220), .CK(
        signal_4640), .Q(signal_3095), .QN() );
  DFF_X1 cell_1113_s_reg_0_s_current_state_reg ( .D(signal_1063), .CK(
        signal_4640), .Q(signal_1746), .QN() );
  DFF_X1 cell_1113_s_reg_1_s_current_state_reg ( .D(signal_4221), .CK(
        signal_4640), .Q(signal_3098), .QN() );
  DFF_X1 cell_1117_s_reg_0_s_current_state_reg ( .D(signal_1066), .CK(
        signal_4640), .Q(signal_1745), .QN() );
  DFF_X1 cell_1117_s_reg_1_s_current_state_reg ( .D(signal_4222), .CK(
        signal_4640), .Q(signal_3101), .QN() );
  DFF_X1 cell_1121_s_reg_0_s_current_state_reg ( .D(signal_1069), .CK(
        signal_4640), .Q(signal_1744), .QN() );
  DFF_X1 cell_1121_s_reg_1_s_current_state_reg ( .D(signal_4223), .CK(
        signal_4640), .Q(signal_3104), .QN() );
  DFF_X1 cell_1125_s_reg_0_s_current_state_reg ( .D(signal_1072), .CK(
        signal_4640), .Q(signal_1743), .QN() );
  DFF_X1 cell_1125_s_reg_1_s_current_state_reg ( .D(signal_4224), .CK(
        signal_4640), .Q(signal_3107), .QN() );
  DFF_X1 cell_1129_s_reg_0_s_current_state_reg ( .D(signal_1075), .CK(
        signal_4640), .Q(signal_1742), .QN() );
  DFF_X1 cell_1129_s_reg_1_s_current_state_reg ( .D(signal_4225), .CK(
        signal_4640), .Q(signal_3110), .QN() );
  DFF_X1 cell_1133_s_reg_0_s_current_state_reg ( .D(signal_1078), .CK(
        signal_4640), .Q(signal_1733), .QN() );
  DFF_X1 cell_1133_s_reg_1_s_current_state_reg ( .D(signal_4066), .CK(
        signal_4640), .Q(signal_3113), .QN() );
  DFF_X1 cell_1137_s_reg_0_s_current_state_reg ( .D(signal_1081), .CK(
        signal_4640), .Q(signal_1732), .QN() );
  DFF_X1 cell_1137_s_reg_1_s_current_state_reg ( .D(signal_4067), .CK(
        signal_4640), .Q(signal_3116), .QN() );
  DFF_X1 cell_1141_s_reg_0_s_current_state_reg ( .D(signal_1084), .CK(
        signal_4640), .Q(signal_1731), .QN() );
  DFF_X1 cell_1141_s_reg_1_s_current_state_reg ( .D(signal_4068), .CK(
        signal_4640), .Q(signal_3119), .QN() );
  DFF_X1 cell_1145_s_reg_0_s_current_state_reg ( .D(signal_1087), .CK(
        signal_4640), .Q(signal_1730), .QN() );
  DFF_X1 cell_1145_s_reg_1_s_current_state_reg ( .D(signal_4069), .CK(
        signal_4640), .Q(signal_3122), .QN() );
  DFF_X1 cell_1149_s_reg_0_s_current_state_reg ( .D(signal_1090), .CK(
        signal_4640), .Q(signal_1729), .QN() );
  DFF_X1 cell_1149_s_reg_1_s_current_state_reg ( .D(signal_4070), .CK(
        signal_4640), .Q(signal_3125), .QN() );
  DFF_X1 cell_1153_s_reg_0_s_current_state_reg ( .D(signal_1093), .CK(
        signal_4640), .Q(signal_1728), .QN() );
  DFF_X1 cell_1153_s_reg_1_s_current_state_reg ( .D(signal_4071), .CK(
        signal_4640), .Q(signal_3128), .QN() );
  DFF_X1 cell_1157_s_reg_0_s_current_state_reg ( .D(signal_1096), .CK(
        signal_4640), .Q(signal_1727), .QN() );
  DFF_X1 cell_1157_s_reg_1_s_current_state_reg ( .D(signal_4072), .CK(
        signal_4640), .Q(signal_3131), .QN() );
  DFF_X1 cell_1161_s_reg_0_s_current_state_reg ( .D(signal_1099), .CK(
        signal_4640), .Q(signal_1726), .QN() );
  DFF_X1 cell_1161_s_reg_1_s_current_state_reg ( .D(signal_4073), .CK(
        signal_4640), .Q(signal_3134), .QN() );
  DFF_X1 cell_1165_s_reg_0_s_current_state_reg ( .D(signal_1102), .CK(
        signal_4640), .Q(signal_1717), .QN() );
  DFF_X1 cell_1165_s_reg_1_s_current_state_reg ( .D(signal_4074), .CK(
        signal_4640), .Q(signal_3137), .QN() );
  DFF_X1 cell_1169_s_reg_0_s_current_state_reg ( .D(signal_1105), .CK(
        signal_4640), .Q(signal_1716), .QN() );
  DFF_X1 cell_1169_s_reg_1_s_current_state_reg ( .D(signal_4075), .CK(
        signal_4640), .Q(signal_3140), .QN() );
  DFF_X1 cell_1173_s_reg_0_s_current_state_reg ( .D(signal_1108), .CK(
        signal_4640), .Q(signal_1715), .QN() );
  DFF_X1 cell_1173_s_reg_1_s_current_state_reg ( .D(signal_4076), .CK(
        signal_4640), .Q(signal_3143), .QN() );
  DFF_X1 cell_1177_s_reg_0_s_current_state_reg ( .D(signal_1111), .CK(
        signal_4640), .Q(signal_1714), .QN() );
  DFF_X1 cell_1177_s_reg_1_s_current_state_reg ( .D(signal_4077), .CK(
        signal_4640), .Q(signal_3146), .QN() );
  DFF_X1 cell_1181_s_reg_0_s_current_state_reg ( .D(signal_1114), .CK(
        signal_4640), .Q(signal_1713), .QN() );
  DFF_X1 cell_1181_s_reg_1_s_current_state_reg ( .D(signal_4078), .CK(
        signal_4640), .Q(signal_3149), .QN() );
  DFF_X1 cell_1185_s_reg_0_s_current_state_reg ( .D(signal_1117), .CK(
        signal_4640), .Q(signal_1712), .QN() );
  DFF_X1 cell_1185_s_reg_1_s_current_state_reg ( .D(signal_4079), .CK(
        signal_4640), .Q(signal_3152), .QN() );
  DFF_X1 cell_1189_s_reg_0_s_current_state_reg ( .D(signal_1120), .CK(
        signal_4640), .Q(signal_1711), .QN() );
  DFF_X1 cell_1189_s_reg_1_s_current_state_reg ( .D(signal_4080), .CK(
        signal_4640), .Q(signal_3155), .QN() );
  DFF_X1 cell_1193_s_reg_0_s_current_state_reg ( .D(signal_1123), .CK(
        signal_4640), .Q(signal_1710), .QN() );
  DFF_X1 cell_1193_s_reg_1_s_current_state_reg ( .D(signal_4081), .CK(
        signal_4640), .Q(signal_3158), .QN() );
  DFF_X1 cell_1197_s_reg_0_s_current_state_reg ( .D(signal_1126), .CK(
        signal_4640), .Q(signal_1701), .QN() );
  DFF_X1 cell_1197_s_reg_1_s_current_state_reg ( .D(signal_4082), .CK(
        signal_4640), .Q(signal_3161), .QN() );
  DFF_X1 cell_1201_s_reg_0_s_current_state_reg ( .D(signal_1129), .CK(
        signal_4640), .Q(signal_1700), .QN() );
  DFF_X1 cell_1201_s_reg_1_s_current_state_reg ( .D(signal_4083), .CK(
        signal_4640), .Q(signal_3164), .QN() );
  DFF_X1 cell_1205_s_reg_0_s_current_state_reg ( .D(signal_1132), .CK(
        signal_4640), .Q(signal_1699), .QN() );
  DFF_X1 cell_1205_s_reg_1_s_current_state_reg ( .D(signal_4084), .CK(
        signal_4640), .Q(signal_3167), .QN() );
  DFF_X1 cell_1209_s_reg_0_s_current_state_reg ( .D(signal_1135), .CK(
        signal_4640), .Q(signal_1698), .QN() );
  DFF_X1 cell_1209_s_reg_1_s_current_state_reg ( .D(signal_4085), .CK(
        signal_4640), .Q(signal_3170), .QN() );
  DFF_X1 cell_1213_s_reg_0_s_current_state_reg ( .D(signal_1138), .CK(
        signal_4640), .Q(signal_1697), .QN() );
  DFF_X1 cell_1213_s_reg_1_s_current_state_reg ( .D(signal_4086), .CK(
        signal_4640), .Q(signal_3173), .QN() );
  DFF_X1 cell_1217_s_reg_0_s_current_state_reg ( .D(signal_1141), .CK(
        signal_4640), .Q(signal_1696), .QN() );
  DFF_X1 cell_1217_s_reg_1_s_current_state_reg ( .D(signal_4087), .CK(
        signal_4640), .Q(signal_3176), .QN() );
  DFF_X1 cell_1221_s_reg_0_s_current_state_reg ( .D(signal_1144), .CK(
        signal_4640), .Q(signal_1695), .QN() );
  DFF_X1 cell_1221_s_reg_1_s_current_state_reg ( .D(signal_4088), .CK(
        signal_4640), .Q(signal_3179), .QN() );
  DFF_X1 cell_1225_s_reg_0_s_current_state_reg ( .D(signal_1147), .CK(
        signal_4640), .Q(signal_1694), .QN() );
  DFF_X1 cell_1225_s_reg_1_s_current_state_reg ( .D(signal_4089), .CK(
        signal_4640), .Q(signal_3182), .QN() );
endmodule

