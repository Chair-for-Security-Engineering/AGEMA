/* modified netlist. Source: module AES in file AES.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module AES_HPC3_Pipeline_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [271:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire AKSRnotDone ;
    wire LastRoundorDone ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire n55 ;
    wire n56 ;
    wire n57 ;
    wire n58 ;
    wire n59 ;
    wire n60 ;
    wire n61 ;
    wire n62 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire MuxSboxIn_n7 ;
    wire MuxSboxIn_n6 ;
    wire MuxSboxIn_n5 ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire MixColumnsIns_n64 ;
    wire MixColumnsIns_n63 ;
    wire MixColumnsIns_n62 ;
    wire MixColumnsIns_n61 ;
    wire MixColumnsIns_n60 ;
    wire MixColumnsIns_n59 ;
    wire MixColumnsIns_n58 ;
    wire MixColumnsIns_n57 ;
    wire MixColumnsIns_n56 ;
    wire MixColumnsIns_n55 ;
    wire MixColumnsIns_n54 ;
    wire MixColumnsIns_n53 ;
    wire MixColumnsIns_n52 ;
    wire MixColumnsIns_n51 ;
    wire MixColumnsIns_n50 ;
    wire MixColumnsIns_n49 ;
    wire MixColumnsIns_n48 ;
    wire MixColumnsIns_n47 ;
    wire MixColumnsIns_n46 ;
    wire MixColumnsIns_n45 ;
    wire MixColumnsIns_n44 ;
    wire MixColumnsIns_n43 ;
    wire MixColumnsIns_n42 ;
    wire MixColumnsIns_n41 ;
    wire MixColumnsIns_n40 ;
    wire MixColumnsIns_n39 ;
    wire MixColumnsIns_n38 ;
    wire MixColumnsIns_n37 ;
    wire MixColumnsIns_n36 ;
    wire MixColumnsIns_n35 ;
    wire MixColumnsIns_n34 ;
    wire MixColumnsIns_n33 ;
    wire MixColumnsIns_n32 ;
    wire MixColumnsIns_n31 ;
    wire MixColumnsIns_n30 ;
    wire MixColumnsIns_n29 ;
    wire MixColumnsIns_n28 ;
    wire MixColumnsIns_n27 ;
    wire MixColumnsIns_n26 ;
    wire MixColumnsIns_n25 ;
    wire MixColumnsIns_n24 ;
    wire MixColumnsIns_n23 ;
    wire MixColumnsIns_n22 ;
    wire MixColumnsIns_n21 ;
    wire MixColumnsIns_n20 ;
    wire MixColumnsIns_n19 ;
    wire MixColumnsIns_n18 ;
    wire MixColumnsIns_n17 ;
    wire MixColumnsIns_n16 ;
    wire MixColumnsIns_n15 ;
    wire MixColumnsIns_n14 ;
    wire MixColumnsIns_n13 ;
    wire MixColumnsIns_n12 ;
    wire MixColumnsIns_n11 ;
    wire MixColumnsIns_n10 ;
    wire MixColumnsIns_n9 ;
    wire MixColumnsIns_n8 ;
    wire MixColumnsIns_n7 ;
    wire MixColumnsIns_n6 ;
    wire MixColumnsIns_n5 ;
    wire MixColumnsIns_n4 ;
    wire MixColumnsIns_n3 ;
    wire MixColumnsIns_n2 ;
    wire MixColumnsIns_n1 ;
    wire MuxMCOut_n6 ;
    wire MuxMCOut_n5 ;
    wire MuxMCOut_n4 ;
    wire MuxRound_n19 ;
    wire MuxRound_n18 ;
    wire MuxRound_n17 ;
    wire MuxRound_n16 ;
    wire MuxRound_n15 ;
    wire MuxRound_n14 ;
    wire MuxRound_n13 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire MuxKeyExpansion_n21 ;
    wire MuxKeyExpansion_n20 ;
    wire MuxKeyExpansion_n19 ;
    wire MuxKeyExpansion_n18 ;
    wire MuxKeyExpansion_n17 ;
    wire MuxKeyExpansion_n16 ;
    wire MuxKeyExpansion_n15 ;
    wire MuxKeyExpansion_n14 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n42 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n44 ;
    wire RoundCounterIns_n45 ;
    wire InRoundCounterIns_n12 ;
    wire InRoundCounterIns_n11 ;
    wire InRoundCounterIns_n10 ;
    wire InRoundCounterIns_n9 ;
    wire InRoundCounterIns_n8 ;
    wire InRoundCounterIns_n7 ;
    wire InRoundCounterIns_n5 ;
    wire InRoundCounterIns_n4 ;
    wire InRoundCounterIns_n3 ;
    wire InRoundCounterIns_n2 ;
    wire InRoundCounterIns_n1 ;
    wire InRoundCounterIns_n6 ;
    wire InRoundCounterIns_n39 ;
    wire InRoundCounterIns_n40 ;
    wire InRoundCounterIns_n41 ;
    wire [127:0] RoundOutput ;
    wire [127:0] ShiftRowsOutput ;
    wire [31:0] KSSubBytesInput ;
    wire [31:0] SubBytesInput ;
    wire [3:0] SubBytesOutput ;
    wire [31:0] MixColumnsOutput ;
    wire [31:0] ColumnOutput ;
    wire [127:0] RoundKeyOutput ;
    wire [127:32] RoundKey ;
    wire [7:0] Rcon ;
    wire [127:0] KeyExpansionOutput ;
    wire [3:0] RoundCounter ;
    wire [2:0] InRoundCounter ;
    wire [28:0] MixColumnsIns_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2340 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2346 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2352 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2358 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2364 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2370 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2376 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2382 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2388 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2394 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2400 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2406 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2412 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2418 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2424 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2432 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2438 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2444 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2450 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2456 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2462 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2468 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2474 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2580 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2586 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2592 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2598 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2604 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2610 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2616 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2622 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2630 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2636 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2642 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2648 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2654 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2660 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2666 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2672 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2678 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2684 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2690 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2696 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2702 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2708 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2714 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2720 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2728 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2734 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2740 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2746 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2752 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2758 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2764 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2770 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2778 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2784 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2790 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2796 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2802 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2808 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2814 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2820 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2826 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2832 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2838 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2844 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5185 ;
    wire new_AGEMA_signal_5186 ;
    wire new_AGEMA_signal_5187 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5194 ;
    wire new_AGEMA_signal_5195 ;
    wire new_AGEMA_signal_5196 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5203 ;
    wire new_AGEMA_signal_5204 ;
    wire new_AGEMA_signal_5205 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5212 ;
    wire new_AGEMA_signal_5213 ;
    wire new_AGEMA_signal_5214 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5221 ;
    wire new_AGEMA_signal_5222 ;
    wire new_AGEMA_signal_5223 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5230 ;
    wire new_AGEMA_signal_5231 ;
    wire new_AGEMA_signal_5232 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5239 ;
    wire new_AGEMA_signal_5240 ;
    wire new_AGEMA_signal_5241 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5248 ;
    wire new_AGEMA_signal_5249 ;
    wire new_AGEMA_signal_5250 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5257 ;
    wire new_AGEMA_signal_5258 ;
    wire new_AGEMA_signal_5259 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5266 ;
    wire new_AGEMA_signal_5267 ;
    wire new_AGEMA_signal_5268 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5275 ;
    wire new_AGEMA_signal_5276 ;
    wire new_AGEMA_signal_5277 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5284 ;
    wire new_AGEMA_signal_5285 ;
    wire new_AGEMA_signal_5286 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5293 ;
    wire new_AGEMA_signal_5294 ;
    wire new_AGEMA_signal_5295 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5302 ;
    wire new_AGEMA_signal_5303 ;
    wire new_AGEMA_signal_5304 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5311 ;
    wire new_AGEMA_signal_5312 ;
    wire new_AGEMA_signal_5313 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5320 ;
    wire new_AGEMA_signal_5321 ;
    wire new_AGEMA_signal_5322 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5329 ;
    wire new_AGEMA_signal_5330 ;
    wire new_AGEMA_signal_5331 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5338 ;
    wire new_AGEMA_signal_5339 ;
    wire new_AGEMA_signal_5340 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5347 ;
    wire new_AGEMA_signal_5348 ;
    wire new_AGEMA_signal_5349 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5356 ;
    wire new_AGEMA_signal_5357 ;
    wire new_AGEMA_signal_5358 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5365 ;
    wire new_AGEMA_signal_5366 ;
    wire new_AGEMA_signal_5367 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5374 ;
    wire new_AGEMA_signal_5375 ;
    wire new_AGEMA_signal_5376 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5383 ;
    wire new_AGEMA_signal_5384 ;
    wire new_AGEMA_signal_5385 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5392 ;
    wire new_AGEMA_signal_5393 ;
    wire new_AGEMA_signal_5394 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5401 ;
    wire new_AGEMA_signal_5402 ;
    wire new_AGEMA_signal_5403 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5410 ;
    wire new_AGEMA_signal_5411 ;
    wire new_AGEMA_signal_5412 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5419 ;
    wire new_AGEMA_signal_5420 ;
    wire new_AGEMA_signal_5421 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5428 ;
    wire new_AGEMA_signal_5429 ;
    wire new_AGEMA_signal_5430 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5437 ;
    wire new_AGEMA_signal_5438 ;
    wire new_AGEMA_signal_5439 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5446 ;
    wire new_AGEMA_signal_5447 ;
    wire new_AGEMA_signal_5448 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5455 ;
    wire new_AGEMA_signal_5456 ;
    wire new_AGEMA_signal_5457 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5464 ;
    wire new_AGEMA_signal_5465 ;
    wire new_AGEMA_signal_5466 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5473 ;
    wire new_AGEMA_signal_5474 ;
    wire new_AGEMA_signal_5475 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5482 ;
    wire new_AGEMA_signal_5483 ;
    wire new_AGEMA_signal_5484 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5491 ;
    wire new_AGEMA_signal_5492 ;
    wire new_AGEMA_signal_5493 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5500 ;
    wire new_AGEMA_signal_5501 ;
    wire new_AGEMA_signal_5502 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5509 ;
    wire new_AGEMA_signal_5510 ;
    wire new_AGEMA_signal_5511 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5518 ;
    wire new_AGEMA_signal_5519 ;
    wire new_AGEMA_signal_5520 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5527 ;
    wire new_AGEMA_signal_5528 ;
    wire new_AGEMA_signal_5529 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5536 ;
    wire new_AGEMA_signal_5537 ;
    wire new_AGEMA_signal_5538 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5545 ;
    wire new_AGEMA_signal_5546 ;
    wire new_AGEMA_signal_5547 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5554 ;
    wire new_AGEMA_signal_5555 ;
    wire new_AGEMA_signal_5556 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5563 ;
    wire new_AGEMA_signal_5564 ;
    wire new_AGEMA_signal_5565 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5572 ;
    wire new_AGEMA_signal_5573 ;
    wire new_AGEMA_signal_5574 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5581 ;
    wire new_AGEMA_signal_5582 ;
    wire new_AGEMA_signal_5583 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5590 ;
    wire new_AGEMA_signal_5591 ;
    wire new_AGEMA_signal_5592 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5599 ;
    wire new_AGEMA_signal_5600 ;
    wire new_AGEMA_signal_5601 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5608 ;
    wire new_AGEMA_signal_5609 ;
    wire new_AGEMA_signal_5610 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5617 ;
    wire new_AGEMA_signal_5618 ;
    wire new_AGEMA_signal_5619 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5626 ;
    wire new_AGEMA_signal_5627 ;
    wire new_AGEMA_signal_5628 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5635 ;
    wire new_AGEMA_signal_5636 ;
    wire new_AGEMA_signal_5637 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5644 ;
    wire new_AGEMA_signal_5645 ;
    wire new_AGEMA_signal_5646 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5653 ;
    wire new_AGEMA_signal_5654 ;
    wire new_AGEMA_signal_5655 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5662 ;
    wire new_AGEMA_signal_5663 ;
    wire new_AGEMA_signal_5664 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5671 ;
    wire new_AGEMA_signal_5672 ;
    wire new_AGEMA_signal_5673 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5680 ;
    wire new_AGEMA_signal_5681 ;
    wire new_AGEMA_signal_5682 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5689 ;
    wire new_AGEMA_signal_5690 ;
    wire new_AGEMA_signal_5691 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5698 ;
    wire new_AGEMA_signal_5699 ;
    wire new_AGEMA_signal_5700 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;

    /* cells in depth 0 */
    AND2_X1 U323 ( .A1 (n45), .A2 (n44), .ZN (AKSRnotDone) ) ;
    NOR2_X1 U324 ( .A1 (n60), .A2 (n49), .ZN (LastRoundorDone) ) ;
    AND2_X1 U325 ( .A1 (RoundCounter[0]), .A2 (LastRoundorDone), .ZN (done) ) ;
    INV_X1 U326 ( .A (RoundCounter[3]), .ZN (n60) ) ;
    NOR2_X1 U327 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (n45) ) ;
    INV_X1 U328 ( .A (RoundCounter[2]), .ZN (n46) ) ;
    NAND2_X1 U329 ( .A1 (RoundCounter[1]), .A2 (n46), .ZN (n49) ) ;
    NOR2_X1 U330 ( .A1 (done), .A2 (InRoundCounter[2]), .ZN (n44) ) ;
    INV_X1 U331 ( .A (RoundCounter[1]), .ZN (n55) ) ;
    NAND2_X1 U332 ( .A1 (n55), .A2 (n46), .ZN (n47) ) ;
    NOR2_X1 U333 ( .A1 (RoundCounter[0]), .A2 (n47), .ZN (Rcon[0]) ) ;
    NOR2_X1 U334 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n58) ) ;
    NOR2_X1 U335 ( .A1 (n58), .A2 (n47), .ZN (Rcon[1]) ) ;
    NOR2_X1 U336 ( .A1 (RoundCounter[3]), .A2 (n49), .ZN (n48) ) ;
    NOR2_X1 U337 ( .A1 (n60), .A2 (n47), .ZN (n54) ) ;
    MUX2_X1 U338 ( .S (RoundCounter[0]), .A (n48), .B (n54), .Z (Rcon[2]) ) ;
    INV_X1 U339 ( .A (RoundCounter[0]), .ZN (n50) ) ;
    NOR2_X1 U340 ( .A1 (n50), .A2 (n49), .ZN (n51) ) ;
    MUX2_X1 U341 ( .S (RoundCounter[3]), .A (n51), .B (Rcon[0]), .Z (Rcon[3]) ) ;
    NAND2_X1 U342 ( .A1 (RoundCounter[2]), .A2 (n58), .ZN (n52) ) ;
    NOR2_X1 U343 ( .A1 (RoundCounter[1]), .A2 (n52), .ZN (n53) ) ;
    OR2_X1 U344 ( .A1 (n54), .A2 (n53), .ZN (Rcon[4]) ) ;
    XNOR2_X1 U345 ( .A (RoundCounter[2]), .B (RoundCounter[3]), .ZN (n57) ) ;
    NAND2_X1 U346 ( .A1 (RoundCounter[0]), .A2 (n55), .ZN (n56) ) ;
    NOR2_X1 U347 ( .A1 (n57), .A2 (n56), .ZN (Rcon[5]) ) ;
    INV_X1 U348 ( .A (n58), .ZN (n59) ) ;
    NAND2_X1 U349 ( .A1 (RoundCounter[1]), .A2 (RoundCounter[2]), .ZN (n61) ) ;
    NOR2_X1 U350 ( .A1 (n59), .A2 (n61), .ZN (Rcon[6]) ) ;
    NAND2_X1 U351 ( .A1 (RoundCounter[0]), .A2 (n60), .ZN (n62) ) ;
    NOR2_X1 U352 ( .A1 (n62), .A2 (n61), .ZN (Rcon[7]) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U353 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_2339, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2340, ShiftRowsOutput[96]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U354 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({new_AGEMA_signal_2342, RoundKey[100]}), .c ({new_AGEMA_signal_2343, ShiftRowsOutput[68]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U355 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({new_AGEMA_signal_2345, RoundKey[101]}), .c ({new_AGEMA_signal_2346, ShiftRowsOutput[69]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U356 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({new_AGEMA_signal_2348, RoundKey[102]}), .c ({new_AGEMA_signal_2349, ShiftRowsOutput[70]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U357 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({new_AGEMA_signal_2351, RoundKey[103]}), .c ({new_AGEMA_signal_2352, ShiftRowsOutput[71]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U358 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_2354, RoundKey[104]}), .c ({new_AGEMA_signal_2355, ShiftRowsOutput[40]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U359 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({new_AGEMA_signal_2357, RoundKey[105]}), .c ({new_AGEMA_signal_2358, ShiftRowsOutput[41]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U360 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({new_AGEMA_signal_2360, RoundKey[106]}), .c ({new_AGEMA_signal_2361, ShiftRowsOutput[42]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U361 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({new_AGEMA_signal_2363, RoundKey[107]}), .c ({new_AGEMA_signal_2364, ShiftRowsOutput[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U362 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({new_AGEMA_signal_2366, RoundKey[108]}), .c ({new_AGEMA_signal_2367, ShiftRowsOutput[44]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U363 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({new_AGEMA_signal_2369, RoundKey[109]}), .c ({new_AGEMA_signal_2370, ShiftRowsOutput[45]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U364 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({new_AGEMA_signal_2372, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2373, ShiftRowsOutput[74]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U365 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({new_AGEMA_signal_2375, RoundKey[110]}), .c ({new_AGEMA_signal_2376, ShiftRowsOutput[46]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U366 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({new_AGEMA_signal_2378, RoundKey[111]}), .c ({new_AGEMA_signal_2379, ShiftRowsOutput[47]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U367 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_2381, RoundKey[112]}), .c ({new_AGEMA_signal_2382, ShiftRowsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U368 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({new_AGEMA_signal_2384, RoundKey[113]}), .c ({new_AGEMA_signal_2385, ShiftRowsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U369 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({new_AGEMA_signal_2387, RoundKey[114]}), .c ({new_AGEMA_signal_2388, ShiftRowsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U370 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({new_AGEMA_signal_2390, RoundKey[115]}), .c ({new_AGEMA_signal_2391, ShiftRowsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U371 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({new_AGEMA_signal_2393, RoundKey[116]}), .c ({new_AGEMA_signal_2394, ShiftRowsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U372 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({new_AGEMA_signal_2396, RoundKey[117]}), .c ({new_AGEMA_signal_2397, ShiftRowsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U373 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({new_AGEMA_signal_2399, RoundKey[118]}), .c ({new_AGEMA_signal_2400, ShiftRowsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U374 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({new_AGEMA_signal_2402, RoundKey[119]}), .c ({new_AGEMA_signal_2403, ShiftRowsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U375 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({new_AGEMA_signal_2405, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2406, ShiftRowsOutput[75]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U376 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2408, RoundKey[120]}), .c ({new_AGEMA_signal_2409, ShiftRowsOutput[120]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U377 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2411, RoundKey[121]}), .c ({new_AGEMA_signal_2412, ShiftRowsOutput[121]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U378 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2414, RoundKey[122]}), .c ({new_AGEMA_signal_2415, ShiftRowsOutput[122]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U379 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2417, RoundKey[123]}), .c ({new_AGEMA_signal_2418, ShiftRowsOutput[123]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U380 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2420, RoundKey[124]}), .c ({new_AGEMA_signal_2421, ShiftRowsOutput[124]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U381 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2423, RoundKey[125]}), .c ({new_AGEMA_signal_2424, ShiftRowsOutput[125]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U382 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2426, RoundKey[126]}), .c ({new_AGEMA_signal_2427, ShiftRowsOutput[126]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U383 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2429, RoundKey[127]}), .c ({new_AGEMA_signal_2430, ShiftRowsOutput[127]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U384 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({new_AGEMA_signal_2432, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2433, ShiftRowsOutput[76]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U385 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({new_AGEMA_signal_2435, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2436, ShiftRowsOutput[77]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U386 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({new_AGEMA_signal_2438, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2439, ShiftRowsOutput[78]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U387 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({new_AGEMA_signal_2441, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2442, ShiftRowsOutput[79]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U388 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_2444, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2445, ShiftRowsOutput[48]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U389 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({new_AGEMA_signal_2447, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2448, ShiftRowsOutput[49]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U390 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({new_AGEMA_signal_2450, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2451, ShiftRowsOutput[50]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U391 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({new_AGEMA_signal_2453, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2454, ShiftRowsOutput[51]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U392 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({new_AGEMA_signal_2456, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2457, ShiftRowsOutput[97]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U393 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({new_AGEMA_signal_2459, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2460, ShiftRowsOutput[52]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U394 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({new_AGEMA_signal_2462, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2463, ShiftRowsOutput[53]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U395 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({new_AGEMA_signal_2465, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2466, ShiftRowsOutput[54]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U396 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({new_AGEMA_signal_2468, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2469, ShiftRowsOutput[55]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U397 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2471, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2472, ShiftRowsOutput[24]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U398 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2474, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2475, ShiftRowsOutput[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U399 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_2477, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2478, ShiftRowsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U400 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2480, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2481, ShiftRowsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U401 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2483, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2484, ShiftRowsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U402 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2486, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2487, ShiftRowsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U403 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({new_AGEMA_signal_2489, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2490, ShiftRowsOutput[98]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U404 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2492, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2493, ShiftRowsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U405 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2495, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2496, ShiftRowsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U406 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_2498, RoundKey[32]}), .c ({new_AGEMA_signal_2499, ShiftRowsOutput[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U407 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({new_AGEMA_signal_2501, RoundKey[33]}), .c ({new_AGEMA_signal_2502, ShiftRowsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U408 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({new_AGEMA_signal_2504, RoundKey[34]}), .c ({new_AGEMA_signal_2505, ShiftRowsOutput[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U409 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({new_AGEMA_signal_2507, RoundKey[35]}), .c ({new_AGEMA_signal_2508, ShiftRowsOutput[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U410 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({new_AGEMA_signal_2510, RoundKey[36]}), .c ({new_AGEMA_signal_2511, ShiftRowsOutput[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U411 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({new_AGEMA_signal_2513, RoundKey[37]}), .c ({new_AGEMA_signal_2514, ShiftRowsOutput[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U412 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({new_AGEMA_signal_2516, RoundKey[38]}), .c ({new_AGEMA_signal_2517, ShiftRowsOutput[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U413 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({new_AGEMA_signal_2519, RoundKey[39]}), .c ({new_AGEMA_signal_2520, ShiftRowsOutput[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U414 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({new_AGEMA_signal_2522, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2523, ShiftRowsOutput[99]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U415 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_2525, RoundKey[40]}), .c ({new_AGEMA_signal_2526, ShiftRowsOutput[104]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U416 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({new_AGEMA_signal_2528, RoundKey[41]}), .c ({new_AGEMA_signal_2529, ShiftRowsOutput[105]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U417 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({new_AGEMA_signal_2531, RoundKey[42]}), .c ({new_AGEMA_signal_2532, ShiftRowsOutput[106]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U418 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({new_AGEMA_signal_2534, RoundKey[43]}), .c ({new_AGEMA_signal_2535, ShiftRowsOutput[107]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U419 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({new_AGEMA_signal_2537, RoundKey[44]}), .c ({new_AGEMA_signal_2538, ShiftRowsOutput[108]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U420 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({new_AGEMA_signal_2540, RoundKey[45]}), .c ({new_AGEMA_signal_2541, ShiftRowsOutput[109]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U421 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({new_AGEMA_signal_2543, RoundKey[46]}), .c ({new_AGEMA_signal_2544, ShiftRowsOutput[110]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U422 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({new_AGEMA_signal_2546, RoundKey[47]}), .c ({new_AGEMA_signal_2547, ShiftRowsOutput[111]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U423 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_2549, RoundKey[48]}), .c ({new_AGEMA_signal_2550, ShiftRowsOutput[80]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U424 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({new_AGEMA_signal_2552, RoundKey[49]}), .c ({new_AGEMA_signal_2553, ShiftRowsOutput[81]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U425 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({new_AGEMA_signal_2555, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2556, ShiftRowsOutput[100]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U426 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({new_AGEMA_signal_2558, RoundKey[50]}), .c ({new_AGEMA_signal_2559, ShiftRowsOutput[82]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U427 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({new_AGEMA_signal_2561, RoundKey[51]}), .c ({new_AGEMA_signal_2562, ShiftRowsOutput[83]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U428 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({new_AGEMA_signal_2564, RoundKey[52]}), .c ({new_AGEMA_signal_2565, ShiftRowsOutput[84]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U429 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({new_AGEMA_signal_2567, RoundKey[53]}), .c ({new_AGEMA_signal_2568, ShiftRowsOutput[85]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U430 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({new_AGEMA_signal_2570, RoundKey[54]}), .c ({new_AGEMA_signal_2571, ShiftRowsOutput[86]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U431 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({new_AGEMA_signal_2573, RoundKey[55]}), .c ({new_AGEMA_signal_2574, ShiftRowsOutput[87]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U432 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_2576, RoundKey[56]}), .c ({new_AGEMA_signal_2577, ShiftRowsOutput[56]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U433 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2579, RoundKey[57]}), .c ({new_AGEMA_signal_2580, ShiftRowsOutput[57]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U434 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_2582, RoundKey[58]}), .c ({new_AGEMA_signal_2583, ShiftRowsOutput[58]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U435 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2585, RoundKey[59]}), .c ({new_AGEMA_signal_2586, ShiftRowsOutput[59]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U436 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({new_AGEMA_signal_2588, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_2589, ShiftRowsOutput[101]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U437 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2591, RoundKey[60]}), .c ({new_AGEMA_signal_2592, ShiftRowsOutput[60]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U438 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2594, RoundKey[61]}), .c ({new_AGEMA_signal_2595, ShiftRowsOutput[61]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U439 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2597, RoundKey[62]}), .c ({new_AGEMA_signal_2598, ShiftRowsOutput[62]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U440 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2600, RoundKey[63]}), .c ({new_AGEMA_signal_2601, ShiftRowsOutput[63]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U441 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_2603, RoundKey[64]}), .c ({new_AGEMA_signal_2604, ShiftRowsOutput[32]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U442 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({new_AGEMA_signal_2606, RoundKey[65]}), .c ({new_AGEMA_signal_2607, ShiftRowsOutput[33]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U443 ( .a ({ciphertext_s1[98], ciphertext_s0[98]}), .b ({new_AGEMA_signal_2609, RoundKey[66]}), .c ({new_AGEMA_signal_2610, ShiftRowsOutput[34]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U444 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({new_AGEMA_signal_2612, RoundKey[67]}), .c ({new_AGEMA_signal_2613, ShiftRowsOutput[35]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U445 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({new_AGEMA_signal_2615, RoundKey[68]}), .c ({new_AGEMA_signal_2616, ShiftRowsOutput[36]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U446 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({new_AGEMA_signal_2618, RoundKey[69]}), .c ({new_AGEMA_signal_2619, ShiftRowsOutput[37]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U447 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({new_AGEMA_signal_2621, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_2622, ShiftRowsOutput[102]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U448 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({new_AGEMA_signal_2624, RoundKey[70]}), .c ({new_AGEMA_signal_2625, ShiftRowsOutput[38]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U449 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({new_AGEMA_signal_2627, RoundKey[71]}), .c ({new_AGEMA_signal_2628, ShiftRowsOutput[39]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U450 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_2630, RoundKey[72]}), .c ({new_AGEMA_signal_2631, ShiftRowsOutput[8]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U451 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({new_AGEMA_signal_2633, RoundKey[73]}), .c ({new_AGEMA_signal_2634, ShiftRowsOutput[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U452 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({new_AGEMA_signal_2636, RoundKey[74]}), .c ({new_AGEMA_signal_2637, ShiftRowsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U453 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({new_AGEMA_signal_2639, RoundKey[75]}), .c ({new_AGEMA_signal_2640, ShiftRowsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U454 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({new_AGEMA_signal_2642, RoundKey[76]}), .c ({new_AGEMA_signal_2643, ShiftRowsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U455 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({new_AGEMA_signal_2645, RoundKey[77]}), .c ({new_AGEMA_signal_2646, ShiftRowsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U456 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({new_AGEMA_signal_2648, RoundKey[78]}), .c ({new_AGEMA_signal_2649, ShiftRowsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U457 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({new_AGEMA_signal_2651, RoundKey[79]}), .c ({new_AGEMA_signal_2652, ShiftRowsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U458 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({new_AGEMA_signal_2654, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_2655, ShiftRowsOutput[103]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U459 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_2657, RoundKey[80]}), .c ({new_AGEMA_signal_2658, ShiftRowsOutput[112]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U460 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({new_AGEMA_signal_2660, RoundKey[81]}), .c ({new_AGEMA_signal_2661, ShiftRowsOutput[113]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U461 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({new_AGEMA_signal_2663, RoundKey[82]}), .c ({new_AGEMA_signal_2664, ShiftRowsOutput[114]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U462 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({new_AGEMA_signal_2666, RoundKey[83]}), .c ({new_AGEMA_signal_2667, ShiftRowsOutput[115]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U463 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({new_AGEMA_signal_2669, RoundKey[84]}), .c ({new_AGEMA_signal_2670, ShiftRowsOutput[116]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U464 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({new_AGEMA_signal_2672, RoundKey[85]}), .c ({new_AGEMA_signal_2673, ShiftRowsOutput[117]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U465 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({new_AGEMA_signal_2675, RoundKey[86]}), .c ({new_AGEMA_signal_2676, ShiftRowsOutput[118]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U466 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({new_AGEMA_signal_2678, RoundKey[87]}), .c ({new_AGEMA_signal_2679, ShiftRowsOutput[119]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U467 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_2681, RoundKey[88]}), .c ({new_AGEMA_signal_2682, ShiftRowsOutput[88]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U468 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2684, RoundKey[89]}), .c ({new_AGEMA_signal_2685, ShiftRowsOutput[89]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U469 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_2687, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_2688, ShiftRowsOutput[72]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U470 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_2690, RoundKey[90]}), .c ({new_AGEMA_signal_2691, ShiftRowsOutput[90]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U471 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2693, RoundKey[91]}), .c ({new_AGEMA_signal_2694, ShiftRowsOutput[91]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U472 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2696, RoundKey[92]}), .c ({new_AGEMA_signal_2697, ShiftRowsOutput[92]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U473 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2699, RoundKey[93]}), .c ({new_AGEMA_signal_2700, ShiftRowsOutput[93]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U474 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2702, RoundKey[94]}), .c ({new_AGEMA_signal_2703, ShiftRowsOutput[94]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U475 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2705, RoundKey[95]}), .c ({new_AGEMA_signal_2706, ShiftRowsOutput[95]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U476 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_2708, RoundKey[96]}), .c ({new_AGEMA_signal_2709, ShiftRowsOutput[64]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U477 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({new_AGEMA_signal_2711, RoundKey[97]}), .c ({new_AGEMA_signal_2712, ShiftRowsOutput[65]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U478 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({new_AGEMA_signal_2714, RoundKey[98]}), .c ({new_AGEMA_signal_2715, ShiftRowsOutput[66]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U479 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({new_AGEMA_signal_2717, RoundKey[99]}), .c ({new_AGEMA_signal_2718, ShiftRowsOutput[67]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U480 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({new_AGEMA_signal_2720, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_2721, ShiftRowsOutput[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2754, RoundOutput[32]}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_2851, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2755, RoundOutput[33]}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_2853, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2756, RoundOutput[34]}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_2855, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2757, RoundOutput[35]}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_2857, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2758, RoundOutput[36]}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_2859, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2759, RoundOutput[37]}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_2861, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2760, RoundOutput[38]}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_2863, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2761, RoundOutput[39]}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_2865, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2762, RoundOutput[40]}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_2867, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2763, RoundOutput[41]}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_2869, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2764, RoundOutput[42]}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_2871, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2765, RoundOutput[43]}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_2873, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2766, RoundOutput[44]}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_2875, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2767, RoundOutput[45]}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_2877, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2768, RoundOutput[46]}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_2879, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2769, RoundOutput[47]}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_2881, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2770, RoundOutput[48]}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_2883, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2771, RoundOutput[49]}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_2885, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2772, RoundOutput[50]}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_2887, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2773, RoundOutput[51]}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_2889, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2774, RoundOutput[52]}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_2891, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2775, RoundOutput[53]}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_2893, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2776, RoundOutput[54]}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_2895, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2777, RoundOutput[55]}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_2897, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2778, RoundOutput[56]}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_2899, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2779, RoundOutput[57]}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_2901, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2780, RoundOutput[58]}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_2903, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2781, RoundOutput[59]}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_2905, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2782, RoundOutput[60]}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_2907, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2783, RoundOutput[61]}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_2909, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2784, RoundOutput[62]}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_2911, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2785, RoundOutput[63]}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_2913, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2786, RoundOutput[64]}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_2915, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2787, RoundOutput[65]}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_2917, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2788, RoundOutput[66]}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_2919, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2789, RoundOutput[67]}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_2921, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2790, RoundOutput[68]}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_2923, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2791, RoundOutput[69]}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_2925, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2792, RoundOutput[70]}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_2927, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2793, RoundOutput[71]}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_2929, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2794, RoundOutput[72]}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_2931, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2795, RoundOutput[73]}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_2933, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2796, RoundOutput[74]}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_2935, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2797, RoundOutput[75]}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_2937, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2798, RoundOutput[76]}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_2939, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2799, RoundOutput[77]}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_2941, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2800, RoundOutput[78]}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_2943, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2801, RoundOutput[79]}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_2945, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2802, RoundOutput[80]}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_2947, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2803, RoundOutput[81]}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_2949, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2804, RoundOutput[82]}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_2951, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2805, RoundOutput[83]}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_2953, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2806, RoundOutput[84]}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_2955, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2807, RoundOutput[85]}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_2957, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2808, RoundOutput[86]}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_2959, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2809, RoundOutput[87]}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_2961, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2810, RoundOutput[88]}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_2963, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2811, RoundOutput[89]}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_2965, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2812, RoundOutput[90]}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_2967, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2813, RoundOutput[91]}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_2969, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2814, RoundOutput[92]}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_2971, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2815, RoundOutput[93]}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_2973, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2816, RoundOutput[94]}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_2975, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2817, RoundOutput[95]}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_2977, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2818, RoundOutput[96]}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_2979, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2819, RoundOutput[97]}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_2981, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2820, RoundOutput[98]}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_2983, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2821, RoundOutput[99]}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_2985, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2822, RoundOutput[100]}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_2987, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2823, RoundOutput[101]}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_2989, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2824, RoundOutput[102]}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_2991, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2825, RoundOutput[103]}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_2993, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2826, RoundOutput[104]}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_2995, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2827, RoundOutput[105]}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_2997, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2828, RoundOutput[106]}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_2999, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2829, RoundOutput[107]}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_3001, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2830, RoundOutput[108]}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_3003, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2831, RoundOutput[109]}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_3005, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2832, RoundOutput[110]}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_3007, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2833, RoundOutput[111]}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_3009, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2834, RoundOutput[112]}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_3011, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2835, RoundOutput[113]}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_3013, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2836, RoundOutput[114]}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_3015, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2837, RoundOutput[115]}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_3017, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2838, RoundOutput[116]}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_3019, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2839, RoundOutput[117]}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_3021, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2840, RoundOutput[118]}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_3023, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2841, RoundOutput[119]}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_3025, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2842, RoundOutput[120]}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_3027, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2843, RoundOutput[121]}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_3029, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2844, RoundOutput[122]}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_3031, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2845, RoundOutput[123]}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_3033, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2846, RoundOutput[124]}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_3035, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2847, RoundOutput[125]}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_3037, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2848, RoundOutput[126]}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_3039, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_2849, RoundOutput[127]}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_3041, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    INV_X1 MuxSboxIn_U3 ( .A (AKSRnotDone), .ZN (MuxSboxIn_n7) ) ;
    INV_X1 MuxSboxIn_U2 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n5) ) ;
    INV_X1 MuxSboxIn_U1 ( .A (MuxSboxIn_n7), .ZN (MuxSboxIn_n6) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_0_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .a ({new_AGEMA_signal_2444, KSSubBytesInput[0]}), .c ({new_AGEMA_signal_2723, SubBytesInput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_1_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .a ({new_AGEMA_signal_2447, KSSubBytesInput[1]}), .c ({new_AGEMA_signal_2724, SubBytesInput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_2_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .a ({new_AGEMA_signal_2450, KSSubBytesInput[2]}), .c ({new_AGEMA_signal_2725, SubBytesInput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_3_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .a ({new_AGEMA_signal_2453, KSSubBytesInput[3]}), .c ({new_AGEMA_signal_2726, SubBytesInput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_4_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .a ({new_AGEMA_signal_2459, KSSubBytesInput[4]}), .c ({new_AGEMA_signal_2727, SubBytesInput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_5_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .a ({new_AGEMA_signal_2462, KSSubBytesInput[5]}), .c ({new_AGEMA_signal_2728, SubBytesInput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_6_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .a ({new_AGEMA_signal_2465, KSSubBytesInput[6]}), .c ({new_AGEMA_signal_2729, SubBytesInput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_7_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .a ({new_AGEMA_signal_2468, KSSubBytesInput[7]}), .c ({new_AGEMA_signal_2730, SubBytesInput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_8_U1 ( .s (AKSRnotDone), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .a ({new_AGEMA_signal_2687, KSSubBytesInput[8]}), .c ({new_AGEMA_signal_2722, SubBytesInput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_9_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .a ({new_AGEMA_signal_2720, KSSubBytesInput[9]}), .c ({new_AGEMA_signal_2731, SubBytesInput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_10_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .a ({new_AGEMA_signal_2372, KSSubBytesInput[10]}), .c ({new_AGEMA_signal_2732, SubBytesInput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_11_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .a ({new_AGEMA_signal_2405, KSSubBytesInput[11]}), .c ({new_AGEMA_signal_2733, SubBytesInput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_12_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .a ({new_AGEMA_signal_2432, KSSubBytesInput[12]}), .c ({new_AGEMA_signal_2734, SubBytesInput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_13_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .a ({new_AGEMA_signal_2435, KSSubBytesInput[13]}), .c ({new_AGEMA_signal_2735, SubBytesInput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_14_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .a ({new_AGEMA_signal_2438, KSSubBytesInput[14]}), .c ({new_AGEMA_signal_2736, SubBytesInput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_15_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .a ({new_AGEMA_signal_2441, KSSubBytesInput[15]}), .c ({new_AGEMA_signal_2737, SubBytesInput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_16_U1 ( .s (MuxSboxIn_n6), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .a ({new_AGEMA_signal_2339, KSSubBytesInput[16]}), .c ({new_AGEMA_signal_2738, SubBytesInput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_17_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .a ({new_AGEMA_signal_2456, KSSubBytesInput[17]}), .c ({new_AGEMA_signal_2739, SubBytesInput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_18_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .a ({new_AGEMA_signal_2489, KSSubBytesInput[18]}), .c ({new_AGEMA_signal_2740, SubBytesInput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_19_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .a ({new_AGEMA_signal_2522, KSSubBytesInput[19]}), .c ({new_AGEMA_signal_2741, SubBytesInput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_20_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .a ({new_AGEMA_signal_2555, KSSubBytesInput[20]}), .c ({new_AGEMA_signal_2742, SubBytesInput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_21_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .a ({new_AGEMA_signal_2588, KSSubBytesInput[21]}), .c ({new_AGEMA_signal_2743, SubBytesInput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_22_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .a ({new_AGEMA_signal_2621, KSSubBytesInput[22]}), .c ({new_AGEMA_signal_2744, SubBytesInput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_23_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .a ({new_AGEMA_signal_2654, KSSubBytesInput[23]}), .c ({new_AGEMA_signal_2745, SubBytesInput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_24_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .a ({new_AGEMA_signal_2471, KSSubBytesInput[24]}), .c ({new_AGEMA_signal_2746, SubBytesInput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_25_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .a ({new_AGEMA_signal_2474, KSSubBytesInput[25]}), .c ({new_AGEMA_signal_2747, SubBytesInput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_26_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .a ({new_AGEMA_signal_2477, KSSubBytesInput[26]}), .c ({new_AGEMA_signal_2748, SubBytesInput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_27_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .a ({new_AGEMA_signal_2480, KSSubBytesInput[27]}), .c ({new_AGEMA_signal_2749, SubBytesInput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_28_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .a ({new_AGEMA_signal_2483, KSSubBytesInput[28]}), .c ({new_AGEMA_signal_2750, SubBytesInput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_29_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .a ({new_AGEMA_signal_2486, KSSubBytesInput[29]}), .c ({new_AGEMA_signal_2751, SubBytesInput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_30_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .a ({new_AGEMA_signal_2492, KSSubBytesInput[30]}), .c ({new_AGEMA_signal_2752, SubBytesInput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxSboxIn_mux_inst_31_U1 ( .s (MuxSboxIn_n5), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .a ({new_AGEMA_signal_2495, KSSubBytesInput[31]}), .c ({new_AGEMA_signal_2753, SubBytesInput[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_2730, SubBytesInput[7]}), .b ({new_AGEMA_signal_2727, SubBytesInput[4]}), .c ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_2730, SubBytesInput[7]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_2730, SubBytesInput[7]}), .b ({new_AGEMA_signal_2724, SubBytesInput[1]}), .c ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_2727, SubBytesInput[4]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_2726, SubBytesInput[3]}), .b ({new_AGEMA_signal_2724, SubBytesInput[1]}), .c ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_2729, SubBytesInput[6]}), .b ({new_AGEMA_signal_2728, SubBytesInput[5]}), .c ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_2723, SubBytesInput[0]}), .b ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_3114, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_2723, SubBytesInput[0]}), .b ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_2729, SubBytesInput[6]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3048, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_2728, SubBytesInput[5]}), .b ({new_AGEMA_signal_2725, SubBytesInput[2]}), .c ({new_AGEMA_signal_3049, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_3084, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_3048, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3116, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3048, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_3085, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_3046, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_3049, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_2727, SubBytesInput[4]}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .c ({new_AGEMA_signal_3050, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3050, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_2724, SubBytesInput[1]}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .c ({new_AGEMA_signal_3051, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_3047, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_3051, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_3119, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_3166, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_3167, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_3120, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3049, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_3089, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_2737, SubBytesInput[15]}), .b ({new_AGEMA_signal_2734, SubBytesInput[12]}), .c ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_2737, SubBytesInput[15]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_2737, SubBytesInput[15]}), .b ({new_AGEMA_signal_2731, SubBytesInput[9]}), .c ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_2734, SubBytesInput[12]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_2733, SubBytesInput[11]}), .b ({new_AGEMA_signal_2731, SubBytesInput[9]}), .c ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_2736, SubBytesInput[14]}), .b ({new_AGEMA_signal_2735, SubBytesInput[13]}), .c ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_2722, SubBytesInput[8]}), .b ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_3127, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_2722, SubBytesInput[8]}), .b ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_2736, SubBytesInput[14]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3058, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_2735, SubBytesInput[13]}), .b ({new_AGEMA_signal_2732, SubBytesInput[10]}), .c ({new_AGEMA_signal_3059, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_3092, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_3058, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3129, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3058, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_3093, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_3056, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_3059, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_2734, SubBytesInput[12]}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .c ({new_AGEMA_signal_3060, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3060, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_2731, SubBytesInput[9]}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .c ({new_AGEMA_signal_3061, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_3057, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_3061, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_3132, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_3175, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_3176, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_3133, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3059, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_3097, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_2745, SubBytesInput[23]}), .b ({new_AGEMA_signal_2742, SubBytesInput[20]}), .c ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_2745, SubBytesInput[23]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_2745, SubBytesInput[23]}), .b ({new_AGEMA_signal_2739, SubBytesInput[17]}), .c ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_2742, SubBytesInput[20]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_2741, SubBytesInput[19]}), .b ({new_AGEMA_signal_2739, SubBytesInput[17]}), .c ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_2744, SubBytesInput[22]}), .b ({new_AGEMA_signal_2743, SubBytesInput[21]}), .c ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_2738, SubBytesInput[16]}), .b ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_3140, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_2738, SubBytesInput[16]}), .b ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_2744, SubBytesInput[22]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3068, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_2743, SubBytesInput[21]}), .b ({new_AGEMA_signal_2740, SubBytesInput[18]}), .c ({new_AGEMA_signal_3069, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_3100, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_3068, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3142, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3068, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_3101, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_3066, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_3069, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_2742, SubBytesInput[20]}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .c ({new_AGEMA_signal_3070, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3070, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_2739, SubBytesInput[17]}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .c ({new_AGEMA_signal_3071, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_3067, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_3071, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_3145, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_3184, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_3185, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_3146, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3069, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_3105, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_2753, SubBytesInput[31]}), .b ({new_AGEMA_signal_2750, SubBytesInput[28]}), .c ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_2753, SubBytesInput[31]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_2753, SubBytesInput[31]}), .b ({new_AGEMA_signal_2747, SubBytesInput[25]}), .c ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_2750, SubBytesInput[28]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_2749, SubBytesInput[27]}), .b ({new_AGEMA_signal_2747, SubBytesInput[25]}), .c ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_2752, SubBytesInput[30]}), .b ({new_AGEMA_signal_2751, SubBytesInput[29]}), .c ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_2746, SubBytesInput[24]}), .b ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_3153, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_2746, SubBytesInput[24]}), .b ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_2752, SubBytesInput[30]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3078, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_2751, SubBytesInput[29]}), .b ({new_AGEMA_signal_2748, SubBytesInput[26]}), .c ({new_AGEMA_signal_3079, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_3108, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_3078, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3155, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3078, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_3109, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_3076, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_3079, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_2750, SubBytesInput[28]}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .c ({new_AGEMA_signal_3080, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3080, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_2747, SubBytesInput[25]}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .c ({new_AGEMA_signal_3081, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_3077, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_3081, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_3158, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_3193, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_3194, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_3159, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3079, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_3113, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    INV_X1 MuxMCOut_U3 ( .A (LastRoundorDone), .ZN (MuxMCOut_n6) ) ;
    INV_X1 MuxMCOut_U2 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n5) ) ;
    INV_X1 MuxMCOut_U1 ( .A (MuxMCOut_n6), .ZN (MuxMCOut_n4) ) ;
    INV_X1 MuxRound_U7 ( .A (AKSRnotDone), .ZN (MuxRound_n19) ) ;
    INV_X1 MuxRound_U6 ( .A (MuxRound_n19), .ZN (MuxRound_n16) ) ;
    INV_X1 MuxRound_U5 ( .A (MuxRound_n19), .ZN (MuxRound_n14) ) ;
    INV_X1 MuxRound_U4 ( .A (MuxRound_n19), .ZN (MuxRound_n13) ) ;
    INV_X1 MuxRound_U3 ( .A (MuxRound_n19), .ZN (MuxRound_n15) ) ;
    INV_X1 MuxRound_U2 ( .A (MuxRound_n19), .ZN (MuxRound_n18) ) ;
    INV_X1 MuxRound_U1 ( .A (MuxRound_n19), .ZN (MuxRound_n17) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_32_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .a ({new_AGEMA_signal_2604, ShiftRowsOutput[32]}), .c ({new_AGEMA_signal_2754, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_33_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .a ({new_AGEMA_signal_2607, ShiftRowsOutput[33]}), .c ({new_AGEMA_signal_2755, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_34_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .a ({new_AGEMA_signal_2610, ShiftRowsOutput[34]}), .c ({new_AGEMA_signal_2756, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_35_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .a ({new_AGEMA_signal_2613, ShiftRowsOutput[35]}), .c ({new_AGEMA_signal_2757, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_36_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .a ({new_AGEMA_signal_2616, ShiftRowsOutput[36]}), .c ({new_AGEMA_signal_2758, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_37_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .a ({new_AGEMA_signal_2619, ShiftRowsOutput[37]}), .c ({new_AGEMA_signal_2759, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_38_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .a ({new_AGEMA_signal_2625, ShiftRowsOutput[38]}), .c ({new_AGEMA_signal_2760, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_39_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .a ({new_AGEMA_signal_2628, ShiftRowsOutput[39]}), .c ({new_AGEMA_signal_2761, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_40_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .a ({new_AGEMA_signal_2355, ShiftRowsOutput[40]}), .c ({new_AGEMA_signal_2762, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_41_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .a ({new_AGEMA_signal_2358, ShiftRowsOutput[41]}), .c ({new_AGEMA_signal_2763, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_42_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .a ({new_AGEMA_signal_2361, ShiftRowsOutput[42]}), .c ({new_AGEMA_signal_2764, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_43_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .a ({new_AGEMA_signal_2364, ShiftRowsOutput[43]}), .c ({new_AGEMA_signal_2765, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_44_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .a ({new_AGEMA_signal_2367, ShiftRowsOutput[44]}), .c ({new_AGEMA_signal_2766, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_45_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .a ({new_AGEMA_signal_2370, ShiftRowsOutput[45]}), .c ({new_AGEMA_signal_2767, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_46_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .a ({new_AGEMA_signal_2376, ShiftRowsOutput[46]}), .c ({new_AGEMA_signal_2768, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_47_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .a ({new_AGEMA_signal_2379, ShiftRowsOutput[47]}), .c ({new_AGEMA_signal_2769, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_48_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .a ({new_AGEMA_signal_2445, ShiftRowsOutput[48]}), .c ({new_AGEMA_signal_2770, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_49_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .a ({new_AGEMA_signal_2448, ShiftRowsOutput[49]}), .c ({new_AGEMA_signal_2771, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_50_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .a ({new_AGEMA_signal_2451, ShiftRowsOutput[50]}), .c ({new_AGEMA_signal_2772, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_51_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .a ({new_AGEMA_signal_2454, ShiftRowsOutput[51]}), .c ({new_AGEMA_signal_2773, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_52_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .a ({new_AGEMA_signal_2460, ShiftRowsOutput[52]}), .c ({new_AGEMA_signal_2774, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_53_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .a ({new_AGEMA_signal_2463, ShiftRowsOutput[53]}), .c ({new_AGEMA_signal_2775, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_54_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .a ({new_AGEMA_signal_2466, ShiftRowsOutput[54]}), .c ({new_AGEMA_signal_2776, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_55_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .a ({new_AGEMA_signal_2469, ShiftRowsOutput[55]}), .c ({new_AGEMA_signal_2777, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_56_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_2577, ShiftRowsOutput[56]}), .c ({new_AGEMA_signal_2778, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_57_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_2580, ShiftRowsOutput[57]}), .c ({new_AGEMA_signal_2779, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_58_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_2583, ShiftRowsOutput[58]}), .c ({new_AGEMA_signal_2780, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_59_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_2586, ShiftRowsOutput[59]}), .c ({new_AGEMA_signal_2781, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_60_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_2592, ShiftRowsOutput[60]}), .c ({new_AGEMA_signal_2782, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_61_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_2595, ShiftRowsOutput[61]}), .c ({new_AGEMA_signal_2783, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_62_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_2598, ShiftRowsOutput[62]}), .c ({new_AGEMA_signal_2784, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_63_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_2601, ShiftRowsOutput[63]}), .c ({new_AGEMA_signal_2785, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_64_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .a ({new_AGEMA_signal_2709, ShiftRowsOutput[64]}), .c ({new_AGEMA_signal_2786, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_65_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .a ({new_AGEMA_signal_2712, ShiftRowsOutput[65]}), .c ({new_AGEMA_signal_2787, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_66_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .a ({new_AGEMA_signal_2715, ShiftRowsOutput[66]}), .c ({new_AGEMA_signal_2788, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_67_U1 ( .s (MuxRound_n18), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .a ({new_AGEMA_signal_2718, ShiftRowsOutput[67]}), .c ({new_AGEMA_signal_2789, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_68_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .a ({new_AGEMA_signal_2343, ShiftRowsOutput[68]}), .c ({new_AGEMA_signal_2790, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_69_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .a ({new_AGEMA_signal_2346, ShiftRowsOutput[69]}), .c ({new_AGEMA_signal_2791, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_70_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .a ({new_AGEMA_signal_2349, ShiftRowsOutput[70]}), .c ({new_AGEMA_signal_2792, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_71_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .a ({new_AGEMA_signal_2352, ShiftRowsOutput[71]}), .c ({new_AGEMA_signal_2793, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_72_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .a ({new_AGEMA_signal_2688, ShiftRowsOutput[72]}), .c ({new_AGEMA_signal_2794, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_73_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .a ({new_AGEMA_signal_2721, ShiftRowsOutput[73]}), .c ({new_AGEMA_signal_2795, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_74_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .a ({new_AGEMA_signal_2373, ShiftRowsOutput[74]}), .c ({new_AGEMA_signal_2796, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_75_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .a ({new_AGEMA_signal_2406, ShiftRowsOutput[75]}), .c ({new_AGEMA_signal_2797, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_76_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .a ({new_AGEMA_signal_2433, ShiftRowsOutput[76]}), .c ({new_AGEMA_signal_2798, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_77_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .a ({new_AGEMA_signal_2436, ShiftRowsOutput[77]}), .c ({new_AGEMA_signal_2799, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_78_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .a ({new_AGEMA_signal_2439, ShiftRowsOutput[78]}), .c ({new_AGEMA_signal_2800, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_79_U1 ( .s (MuxRound_n17), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .a ({new_AGEMA_signal_2442, ShiftRowsOutput[79]}), .c ({new_AGEMA_signal_2801, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_80_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .a ({new_AGEMA_signal_2550, ShiftRowsOutput[80]}), .c ({new_AGEMA_signal_2802, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_81_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .a ({new_AGEMA_signal_2553, ShiftRowsOutput[81]}), .c ({new_AGEMA_signal_2803, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_82_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .a ({new_AGEMA_signal_2559, ShiftRowsOutput[82]}), .c ({new_AGEMA_signal_2804, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_83_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .a ({new_AGEMA_signal_2562, ShiftRowsOutput[83]}), .c ({new_AGEMA_signal_2805, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_84_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .a ({new_AGEMA_signal_2565, ShiftRowsOutput[84]}), .c ({new_AGEMA_signal_2806, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_85_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .a ({new_AGEMA_signal_2568, ShiftRowsOutput[85]}), .c ({new_AGEMA_signal_2807, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_86_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .a ({new_AGEMA_signal_2571, ShiftRowsOutput[86]}), .c ({new_AGEMA_signal_2808, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_87_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .a ({new_AGEMA_signal_2574, ShiftRowsOutput[87]}), .c ({new_AGEMA_signal_2809, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_88_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_2682, ShiftRowsOutput[88]}), .c ({new_AGEMA_signal_2810, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_89_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_2685, ShiftRowsOutput[89]}), .c ({new_AGEMA_signal_2811, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_90_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_2691, ShiftRowsOutput[90]}), .c ({new_AGEMA_signal_2812, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_91_U1 ( .s (MuxRound_n16), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_2694, ShiftRowsOutput[91]}), .c ({new_AGEMA_signal_2813, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_92_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_2697, ShiftRowsOutput[92]}), .c ({new_AGEMA_signal_2814, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_93_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_2700, ShiftRowsOutput[93]}), .c ({new_AGEMA_signal_2815, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_94_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_2703, ShiftRowsOutput[94]}), .c ({new_AGEMA_signal_2816, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_95_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_2706, ShiftRowsOutput[95]}), .c ({new_AGEMA_signal_2817, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_96_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .a ({new_AGEMA_signal_2340, ShiftRowsOutput[96]}), .c ({new_AGEMA_signal_2818, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_97_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .a ({new_AGEMA_signal_2457, ShiftRowsOutput[97]}), .c ({new_AGEMA_signal_2819, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_98_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .a ({new_AGEMA_signal_2490, ShiftRowsOutput[98]}), .c ({new_AGEMA_signal_2820, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_99_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .a ({new_AGEMA_signal_2523, ShiftRowsOutput[99]}), .c ({new_AGEMA_signal_2821, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_100_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .a ({new_AGEMA_signal_2556, ShiftRowsOutput[100]}), .c ({new_AGEMA_signal_2822, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_101_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .a ({new_AGEMA_signal_2589, ShiftRowsOutput[101]}), .c ({new_AGEMA_signal_2823, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_102_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .a ({new_AGEMA_signal_2622, ShiftRowsOutput[102]}), .c ({new_AGEMA_signal_2824, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_103_U1 ( .s (MuxRound_n15), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .a ({new_AGEMA_signal_2655, ShiftRowsOutput[103]}), .c ({new_AGEMA_signal_2825, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_104_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .a ({new_AGEMA_signal_2526, ShiftRowsOutput[104]}), .c ({new_AGEMA_signal_2826, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_105_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .a ({new_AGEMA_signal_2529, ShiftRowsOutput[105]}), .c ({new_AGEMA_signal_2827, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_106_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .a ({new_AGEMA_signal_2532, ShiftRowsOutput[106]}), .c ({new_AGEMA_signal_2828, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_107_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .a ({new_AGEMA_signal_2535, ShiftRowsOutput[107]}), .c ({new_AGEMA_signal_2829, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_108_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .a ({new_AGEMA_signal_2538, ShiftRowsOutput[108]}), .c ({new_AGEMA_signal_2830, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_109_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .a ({new_AGEMA_signal_2541, ShiftRowsOutput[109]}), .c ({new_AGEMA_signal_2831, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_110_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .a ({new_AGEMA_signal_2544, ShiftRowsOutput[110]}), .c ({new_AGEMA_signal_2832, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_111_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .a ({new_AGEMA_signal_2547, ShiftRowsOutput[111]}), .c ({new_AGEMA_signal_2833, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_112_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .a ({new_AGEMA_signal_2658, ShiftRowsOutput[112]}), .c ({new_AGEMA_signal_2834, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_113_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .a ({new_AGEMA_signal_2661, ShiftRowsOutput[113]}), .c ({new_AGEMA_signal_2835, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_114_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .a ({new_AGEMA_signal_2664, ShiftRowsOutput[114]}), .c ({new_AGEMA_signal_2836, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_115_U1 ( .s (MuxRound_n14), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .a ({new_AGEMA_signal_2667, ShiftRowsOutput[115]}), .c ({new_AGEMA_signal_2837, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_116_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .a ({new_AGEMA_signal_2670, ShiftRowsOutput[116]}), .c ({new_AGEMA_signal_2838, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_117_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .a ({new_AGEMA_signal_2673, ShiftRowsOutput[117]}), .c ({new_AGEMA_signal_2839, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_118_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .a ({new_AGEMA_signal_2676, ShiftRowsOutput[118]}), .c ({new_AGEMA_signal_2840, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_119_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .a ({new_AGEMA_signal_2679, ShiftRowsOutput[119]}), .c ({new_AGEMA_signal_2841, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_120_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_2409, ShiftRowsOutput[120]}), .c ({new_AGEMA_signal_2842, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_121_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_2412, ShiftRowsOutput[121]}), .c ({new_AGEMA_signal_2843, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_122_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_2415, ShiftRowsOutput[122]}), .c ({new_AGEMA_signal_2844, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_123_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_2418, ShiftRowsOutput[123]}), .c ({new_AGEMA_signal_2845, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_124_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_2421, ShiftRowsOutput[124]}), .c ({new_AGEMA_signal_2846, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_125_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_2424, ShiftRowsOutput[125]}), .c ({new_AGEMA_signal_2847, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_126_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_2427, ShiftRowsOutput[126]}), .c ({new_AGEMA_signal_2848, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_127_U1 ( .s (MuxRound_n13), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_2430, ShiftRowsOutput[127]}), .c ({new_AGEMA_signal_2849, RoundOutput[127]}) ) ;
    INV_X1 MuxKeyExpansion_U8 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n14) ) ;
    INV_X1 MuxKeyExpansion_U7 ( .A (AKSRnotDone), .ZN (MuxKeyExpansion_n21) ) ;
    INV_X1 MuxKeyExpansion_U6 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n16) ) ;
    INV_X1 MuxKeyExpansion_U5 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n17) ) ;
    INV_X1 MuxKeyExpansion_U4 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n18) ) ;
    INV_X1 MuxKeyExpansion_U3 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n19) ) ;
    INV_X1 MuxKeyExpansion_U2 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n20) ) ;
    INV_X1 MuxKeyExpansion_U1 ( .A (MuxKeyExpansion_n21), .ZN (MuxKeyExpansion_n15) ) ;
    NOR2_X1 RoundCounterIns_U11 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_n45) ) ;
    XNOR2_X1 RoundCounterIns_U10 ( .A (RoundCounter[0]), .B (AKSRnotDone), .ZN (RoundCounterIns_n10) ) ;
    NOR2_X1 RoundCounterIns_U9 ( .A1 (reset), .A2 (RoundCounterIns_n9), .ZN (RoundCounterIns_n44) ) ;
    XOR2_X1 RoundCounterIns_U8 ( .A (RoundCounter[1]), .B (RoundCounterIns_n8), .Z (RoundCounterIns_n9) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (reset), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n42) ) ;
    XOR2_X1 RoundCounterIns_U6 ( .A (RoundCounter[3]), .B (RoundCounterIns_n6), .Z (RoundCounterIns_n7) ) ;
    NAND2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounter[2]), .ZN (RoundCounterIns_n6) ) ;
    NOR2_X1 RoundCounterIns_U4 ( .A1 (reset), .A2 (RoundCounterIns_n4), .ZN (RoundCounterIns_n1) ) ;
    XNOR2_X1 RoundCounterIns_U3 ( .A (RoundCounter[2]), .B (RoundCounterIns_n5), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (RoundCounterIns_n2), .A2 (RoundCounterIns_n8), .ZN (RoundCounterIns_n5) ) ;
    NAND2_X1 RoundCounterIns_U1 ( .A1 (AKSRnotDone), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_n8) ) ;
    INV_X1 RoundCounterIns_count_reg_1__U1 ( .A (RoundCounter[1]), .ZN (RoundCounterIns_n2) ) ;
    NOR2_X1 InRoundCounterIns_U13 ( .A1 (reset), .A2 (InRoundCounterIns_n12), .ZN (InRoundCounterIns_n41) ) ;
    XOR2_X1 InRoundCounterIns_U12 ( .A (InRoundCounter[0]), .B (InRoundCounterIns_n11), .Z (InRoundCounterIns_n12) ) ;
    NAND2_X1 InRoundCounterIns_U11 ( .A1 (InRoundCounterIns_n10), .A2 (1'b1), .ZN (InRoundCounterIns_n11) ) ;
    NAND2_X1 InRoundCounterIns_U10 ( .A1 (InRoundCounterIns_n9), .A2 (InRoundCounter[2]), .ZN (InRoundCounterIns_n10) ) ;
    NAND2_X1 InRoundCounterIns_U9 ( .A1 (InRoundCounter[0]), .A2 (InRoundCounter[1]), .ZN (InRoundCounterIns_n9) ) ;
    NOR2_X1 InRoundCounterIns_U8 ( .A1 (reset), .A2 (InRoundCounterIns_n8), .ZN (InRoundCounterIns_n40) ) ;
    MUX2_X1 InRoundCounterIns_U7 ( .S (InRoundCounter[1]), .A (InRoundCounterIns_n7), .B (InRoundCounterIns_n5), .Z (InRoundCounterIns_n8) ) ;
    NOR2_X1 InRoundCounterIns_U6 ( .A1 (reset), .A2 (InRoundCounterIns_n4), .ZN (InRoundCounterIns_n39) ) ;
    NOR2_X1 InRoundCounterIns_U5 ( .A1 (InRoundCounterIns_n3), .A2 (InRoundCounterIns_n2), .ZN (InRoundCounterIns_n4) ) ;
    NOR2_X1 InRoundCounterIns_U4 ( .A1 (InRoundCounterIns_n1), .A2 (InRoundCounterIns_n7), .ZN (InRoundCounterIns_n2) ) ;
    NAND2_X1 InRoundCounterIns_U3 ( .A1 (InRoundCounterIns_n5), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n7) ) ;
    AND2_X1 InRoundCounterIns_U2 ( .A1 (InRoundCounter[0]), .A2 (1'b1), .ZN (InRoundCounterIns_n5) ) ;
    NOR2_X1 InRoundCounterIns_U1 ( .A1 (1'b1), .A2 (InRoundCounterIns_n6), .ZN (InRoundCounterIns_n3) ) ;
    INV_X1 InRoundCounterIns_count_reg_1__U1 ( .A (InRoundCounter[1]), .ZN (InRoundCounterIns_n1) ) ;
    INV_X1 InRoundCounterIns_count_reg_2__U1 ( .A (InRoundCounter[2]), .ZN (InRoundCounterIns_n6) ) ;

    /* cells in depth 1 */
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_3084, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_3082, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_3121, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_3119, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_3114, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[3], Fresh[2]}), .c ({new_AGEMA_signal_3168, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_4583, new_AGEMA_signal_4582}), .b ({new_AGEMA_signal_3121, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_3169, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_3087, SubBytesIns_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_2723, SubBytesInput[0]}), .clk (clk), .r ({Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_3122, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_3122, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_3121, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_3170, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_3044, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_3086, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_3123, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_3088, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_3083, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[9], Fresh[8]}), .c ({new_AGEMA_signal_3124, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_4585, new_AGEMA_signal_4584}), .b ({new_AGEMA_signal_3123, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_3171, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_3118, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_3117, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_3172, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_3172, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_3123, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_3202, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_3042, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_3085, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_3125, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_3045, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_3089, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[15], Fresh[14]}), .c ({new_AGEMA_signal_3126, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_3126, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_3125, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_3173, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_3043, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_3115, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[17], Fresh[16]}), .c ({new_AGEMA_signal_3174, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_3174, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_3125, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_3203, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_3169, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_3168, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_3204, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_3170, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_4587, new_AGEMA_signal_4586}), .c ({new_AGEMA_signal_3205, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_3171, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_3124, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_3206, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_3202, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_3203, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_3222, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_3204, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_3173, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_3205, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_3203, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_3206, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_3173, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_3222, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_4589, new_AGEMA_signal_4588}), .c ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_3254, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_3240, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_3092, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_3090, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_3134, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_3132, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_3127, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_3177, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_4591, new_AGEMA_signal_4590}), .b ({new_AGEMA_signal_3134, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_3178, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_3095, SubBytesIns_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_2722, SubBytesInput[8]}), .clk (clk), .r ({Fresh[23], Fresh[22]}), .c ({new_AGEMA_signal_3135, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_3135, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_3134, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_3179, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_3054, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_3094, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_3136, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_3096, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_3091, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[27], Fresh[26]}), .c ({new_AGEMA_signal_3137, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_4593, new_AGEMA_signal_4592}), .b ({new_AGEMA_signal_3136, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_3180, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_3131, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_3130, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[29], Fresh[28]}), .c ({new_AGEMA_signal_3181, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_3181, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_3136, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_3207, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_3052, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_3093, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_3138, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_3055, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_3097, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[33], Fresh[32]}), .c ({new_AGEMA_signal_3139, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_3139, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_3138, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_3182, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_3053, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_3128, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[35], Fresh[34]}), .c ({new_AGEMA_signal_3183, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_3183, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_3138, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_3208, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_3178, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_3177, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_3209, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_3179, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_4595, new_AGEMA_signal_4594}), .c ({new_AGEMA_signal_3210, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_3180, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_3137, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_3211, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_3207, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_3208, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_3226, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_3209, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_3182, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_3210, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_3208, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_3211, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_3182, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_3226, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596}), .c ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_3259, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_3244, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_3100, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_3098, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_3147, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_3145, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_3140, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[39], Fresh[38]}), .c ({new_AGEMA_signal_3186, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_4599, new_AGEMA_signal_4598}), .b ({new_AGEMA_signal_3147, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_3187, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_3103, SubBytesIns_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_2738, SubBytesInput[16]}), .clk (clk), .r ({Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_3148, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_3148, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_3147, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_3188, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_3064, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_3102, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_3149, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_3104, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_3099, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[45], Fresh[44]}), .c ({new_AGEMA_signal_3150, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_4601, new_AGEMA_signal_4600}), .b ({new_AGEMA_signal_3149, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_3189, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_3144, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_3143, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[47], Fresh[46]}), .c ({new_AGEMA_signal_3190, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_3190, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_3149, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_3212, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_3062, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_3101, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_3151, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_3065, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_3105, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_3152, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_3152, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_3151, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_3191, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_3063, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_3141, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[53], Fresh[52]}), .c ({new_AGEMA_signal_3192, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_3192, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_3151, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_3213, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_3187, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_3186, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_3214, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_3188, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_4603, new_AGEMA_signal_4602}), .c ({new_AGEMA_signal_3215, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_3189, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_3150, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_3216, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_3212, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_3213, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_3230, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_3214, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_3191, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_3215, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_3213, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_3216, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_3191, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_3230, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604}), .c ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_3264, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_3248, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_3108, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_3106, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_3160, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_3158, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_3153, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[57], Fresh[56]}), .c ({new_AGEMA_signal_3195, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_4607, new_AGEMA_signal_4606}), .b ({new_AGEMA_signal_3160, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_3196, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_3111, SubBytesIns_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_2746, SubBytesInput[24]}), .clk (clk), .r ({Fresh[59], Fresh[58]}), .c ({new_AGEMA_signal_3161, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_3161, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_3160, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_3197, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_3074, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_3110, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_3162, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_3112, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_3107, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[63], Fresh[62]}), .c ({new_AGEMA_signal_3163, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_4609, new_AGEMA_signal_4608}), .b ({new_AGEMA_signal_3162, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_3198, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_3157, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_3156, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[65], Fresh[64]}), .c ({new_AGEMA_signal_3199, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_3199, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_3162, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_3217, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_3072, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_3109, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_3164, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_3075, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_3113, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[69], Fresh[68]}), .c ({new_AGEMA_signal_3165, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_3165, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_3164, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_3200, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_3073, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_3154, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[71], Fresh[70]}), .c ({new_AGEMA_signal_3201, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_3201, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_3164, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_3218, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_3196, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_3195, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_3219, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_3197, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_4611, new_AGEMA_signal_4610}), .c ({new_AGEMA_signal_3220, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_3198, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_3163, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_3221, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_3217, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_3218, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_3234, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_3219, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_3200, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_3220, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_3218, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_3221, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_3200, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_3234, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_4613, new_AGEMA_signal_4612}), .c ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_3269, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_3252, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2061 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T14), .Q (new_AGEMA_signal_4582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2062 ( .C (clk), .D (new_AGEMA_signal_3116), .Q (new_AGEMA_signal_4583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2063 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T26), .Q (new_AGEMA_signal_4584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2064 ( .C (clk), .D (new_AGEMA_signal_3120), .Q (new_AGEMA_signal_4585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2065 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T24), .Q (new_AGEMA_signal_4586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2066 ( .C (clk), .D (new_AGEMA_signal_3166), .Q (new_AGEMA_signal_4587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2067 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T25), .Q (new_AGEMA_signal_4588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2068 ( .C (clk), .D (new_AGEMA_signal_3167), .Q (new_AGEMA_signal_4589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2069 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T14), .Q (new_AGEMA_signal_4590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2070 ( .C (clk), .D (new_AGEMA_signal_3129), .Q (new_AGEMA_signal_4591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2071 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T26), .Q (new_AGEMA_signal_4592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2072 ( .C (clk), .D (new_AGEMA_signal_3133), .Q (new_AGEMA_signal_4593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2073 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T24), .Q (new_AGEMA_signal_4594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2074 ( .C (clk), .D (new_AGEMA_signal_3175), .Q (new_AGEMA_signal_4595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2075 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T25), .Q (new_AGEMA_signal_4596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2076 ( .C (clk), .D (new_AGEMA_signal_3176), .Q (new_AGEMA_signal_4597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2077 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T14), .Q (new_AGEMA_signal_4598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2078 ( .C (clk), .D (new_AGEMA_signal_3142), .Q (new_AGEMA_signal_4599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2079 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T26), .Q (new_AGEMA_signal_4600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2080 ( .C (clk), .D (new_AGEMA_signal_3146), .Q (new_AGEMA_signal_4601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2081 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T24), .Q (new_AGEMA_signal_4602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2082 ( .C (clk), .D (new_AGEMA_signal_3184), .Q (new_AGEMA_signal_4603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2083 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T25), .Q (new_AGEMA_signal_4604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2084 ( .C (clk), .D (new_AGEMA_signal_3185), .Q (new_AGEMA_signal_4605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2085 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T14), .Q (new_AGEMA_signal_4606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2086 ( .C (clk), .D (new_AGEMA_signal_3155), .Q (new_AGEMA_signal_4607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2087 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T26), .Q (new_AGEMA_signal_4608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2088 ( .C (clk), .D (new_AGEMA_signal_3159), .Q (new_AGEMA_signal_4609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2089 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T24), .Q (new_AGEMA_signal_4610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2090 ( .C (clk), .D (new_AGEMA_signal_3193), .Q (new_AGEMA_signal_4611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2091 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T25), .Q (new_AGEMA_signal_4612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2092 ( .C (clk), .D (new_AGEMA_signal_3194), .Q (new_AGEMA_signal_4613) ) ;
    buf_clk new_AGEMA_reg_buffer_2157 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_4678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2161 ( .C (clk), .D (plaintext_s0[0]), .Q (new_AGEMA_signal_4682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2165 ( .C (clk), .D (plaintext_s1[0]), .Q (new_AGEMA_signal_4686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2169 ( .C (clk), .D (plaintext_s0[1]), .Q (new_AGEMA_signal_4690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2173 ( .C (clk), .D (plaintext_s1[1]), .Q (new_AGEMA_signal_4694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2177 ( .C (clk), .D (plaintext_s0[2]), .Q (new_AGEMA_signal_4698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2181 ( .C (clk), .D (plaintext_s1[2]), .Q (new_AGEMA_signal_4702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2185 ( .C (clk), .D (plaintext_s0[3]), .Q (new_AGEMA_signal_4706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2189 ( .C (clk), .D (plaintext_s1[3]), .Q (new_AGEMA_signal_4710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2193 ( .C (clk), .D (plaintext_s0[4]), .Q (new_AGEMA_signal_4714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2197 ( .C (clk), .D (plaintext_s1[4]), .Q (new_AGEMA_signal_4718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2201 ( .C (clk), .D (plaintext_s0[5]), .Q (new_AGEMA_signal_4722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2205 ( .C (clk), .D (plaintext_s1[5]), .Q (new_AGEMA_signal_4726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2209 ( .C (clk), .D (plaintext_s0[6]), .Q (new_AGEMA_signal_4730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2213 ( .C (clk), .D (plaintext_s1[6]), .Q (new_AGEMA_signal_4734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2217 ( .C (clk), .D (plaintext_s0[7]), .Q (new_AGEMA_signal_4738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2221 ( .C (clk), .D (plaintext_s1[7]), .Q (new_AGEMA_signal_4742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2225 ( .C (clk), .D (plaintext_s0[8]), .Q (new_AGEMA_signal_4746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2229 ( .C (clk), .D (plaintext_s1[8]), .Q (new_AGEMA_signal_4750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2233 ( .C (clk), .D (plaintext_s0[9]), .Q (new_AGEMA_signal_4754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2237 ( .C (clk), .D (plaintext_s1[9]), .Q (new_AGEMA_signal_4758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2241 ( .C (clk), .D (plaintext_s0[10]), .Q (new_AGEMA_signal_4762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2245 ( .C (clk), .D (plaintext_s1[10]), .Q (new_AGEMA_signal_4766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2249 ( .C (clk), .D (plaintext_s0[11]), .Q (new_AGEMA_signal_4770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2253 ( .C (clk), .D (plaintext_s1[11]), .Q (new_AGEMA_signal_4774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2257 ( .C (clk), .D (plaintext_s0[12]), .Q (new_AGEMA_signal_4778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2261 ( .C (clk), .D (plaintext_s1[12]), .Q (new_AGEMA_signal_4782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2265 ( .C (clk), .D (plaintext_s0[13]), .Q (new_AGEMA_signal_4786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2269 ( .C (clk), .D (plaintext_s1[13]), .Q (new_AGEMA_signal_4790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2273 ( .C (clk), .D (plaintext_s0[14]), .Q (new_AGEMA_signal_4794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2277 ( .C (clk), .D (plaintext_s1[14]), .Q (new_AGEMA_signal_4798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2281 ( .C (clk), .D (plaintext_s0[15]), .Q (new_AGEMA_signal_4802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2285 ( .C (clk), .D (plaintext_s1[15]), .Q (new_AGEMA_signal_4806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2289 ( .C (clk), .D (plaintext_s0[16]), .Q (new_AGEMA_signal_4810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2293 ( .C (clk), .D (plaintext_s1[16]), .Q (new_AGEMA_signal_4814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2297 ( .C (clk), .D (plaintext_s0[17]), .Q (new_AGEMA_signal_4818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2301 ( .C (clk), .D (plaintext_s1[17]), .Q (new_AGEMA_signal_4822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2305 ( .C (clk), .D (plaintext_s0[18]), .Q (new_AGEMA_signal_4826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2309 ( .C (clk), .D (plaintext_s1[18]), .Q (new_AGEMA_signal_4830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2313 ( .C (clk), .D (plaintext_s0[19]), .Q (new_AGEMA_signal_4834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2317 ( .C (clk), .D (plaintext_s1[19]), .Q (new_AGEMA_signal_4838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2321 ( .C (clk), .D (plaintext_s0[20]), .Q (new_AGEMA_signal_4842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2325 ( .C (clk), .D (plaintext_s1[20]), .Q (new_AGEMA_signal_4846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2329 ( .C (clk), .D (plaintext_s0[21]), .Q (new_AGEMA_signal_4850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2333 ( .C (clk), .D (plaintext_s1[21]), .Q (new_AGEMA_signal_4854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2337 ( .C (clk), .D (plaintext_s0[22]), .Q (new_AGEMA_signal_4858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2341 ( .C (clk), .D (plaintext_s1[22]), .Q (new_AGEMA_signal_4862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2345 ( .C (clk), .D (plaintext_s0[23]), .Q (new_AGEMA_signal_4866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2349 ( .C (clk), .D (plaintext_s1[23]), .Q (new_AGEMA_signal_4870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2353 ( .C (clk), .D (plaintext_s0[24]), .Q (new_AGEMA_signal_4874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2357 ( .C (clk), .D (plaintext_s1[24]), .Q (new_AGEMA_signal_4878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2361 ( .C (clk), .D (plaintext_s0[25]), .Q (new_AGEMA_signal_4882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2365 ( .C (clk), .D (plaintext_s1[25]), .Q (new_AGEMA_signal_4886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2369 ( .C (clk), .D (plaintext_s0[26]), .Q (new_AGEMA_signal_4890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2373 ( .C (clk), .D (plaintext_s1[26]), .Q (new_AGEMA_signal_4894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2377 ( .C (clk), .D (plaintext_s0[27]), .Q (new_AGEMA_signal_4898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2381 ( .C (clk), .D (plaintext_s1[27]), .Q (new_AGEMA_signal_4902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2385 ( .C (clk), .D (plaintext_s0[28]), .Q (new_AGEMA_signal_4906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2389 ( .C (clk), .D (plaintext_s1[28]), .Q (new_AGEMA_signal_4910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2393 ( .C (clk), .D (plaintext_s0[29]), .Q (new_AGEMA_signal_4914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2397 ( .C (clk), .D (plaintext_s1[29]), .Q (new_AGEMA_signal_4918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2401 ( .C (clk), .D (plaintext_s0[30]), .Q (new_AGEMA_signal_4922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2405 ( .C (clk), .D (plaintext_s1[30]), .Q (new_AGEMA_signal_4926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2409 ( .C (clk), .D (plaintext_s0[31]), .Q (new_AGEMA_signal_4930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2413 ( .C (clk), .D (plaintext_s1[31]), .Q (new_AGEMA_signal_4934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2417 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T6), .Q (new_AGEMA_signal_4938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2420 ( .C (clk), .D (new_AGEMA_signal_3082), .Q (new_AGEMA_signal_4941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2423 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T8), .Q (new_AGEMA_signal_4944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2426 ( .C (clk), .D (new_AGEMA_signal_3114), .Q (new_AGEMA_signal_4947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2429 ( .C (clk), .D (SubBytesInput[0]), .Q (new_AGEMA_signal_4950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2432 ( .C (clk), .D (new_AGEMA_signal_2723), .Q (new_AGEMA_signal_4953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2435 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T16), .Q (new_AGEMA_signal_4956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2438 ( .C (clk), .D (new_AGEMA_signal_3086), .Q (new_AGEMA_signal_4959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2441 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T9), .Q (new_AGEMA_signal_4962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2444 ( .C (clk), .D (new_AGEMA_signal_3083), .Q (new_AGEMA_signal_4965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2447 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T17), .Q (new_AGEMA_signal_4968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2450 ( .C (clk), .D (new_AGEMA_signal_3117), .Q (new_AGEMA_signal_4971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2453 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T15), .Q (new_AGEMA_signal_4974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2456 ( .C (clk), .D (new_AGEMA_signal_3085), .Q (new_AGEMA_signal_4977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2459 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T27), .Q (new_AGEMA_signal_4980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2462 ( .C (clk), .D (new_AGEMA_signal_3089), .Q (new_AGEMA_signal_4983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2465 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T10), .Q (new_AGEMA_signal_4986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2468 ( .C (clk), .D (new_AGEMA_signal_3115), .Q (new_AGEMA_signal_4989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2471 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T13), .Q (new_AGEMA_signal_4992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2474 ( .C (clk), .D (new_AGEMA_signal_3084), .Q (new_AGEMA_signal_4995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2477 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T23), .Q (new_AGEMA_signal_4998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2480 ( .C (clk), .D (new_AGEMA_signal_3119), .Q (new_AGEMA_signal_5001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2483 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T19), .Q (new_AGEMA_signal_5004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2486 ( .C (clk), .D (new_AGEMA_signal_3087), .Q (new_AGEMA_signal_5007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2489 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T3), .Q (new_AGEMA_signal_5010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2492 ( .C (clk), .D (new_AGEMA_signal_3044), .Q (new_AGEMA_signal_5013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2495 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T22), .Q (new_AGEMA_signal_5016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2498 ( .C (clk), .D (new_AGEMA_signal_3088), .Q (new_AGEMA_signal_5019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2501 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T20), .Q (new_AGEMA_signal_5022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2504 ( .C (clk), .D (new_AGEMA_signal_3118), .Q (new_AGEMA_signal_5025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2507 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T1), .Q (new_AGEMA_signal_5028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2510 ( .C (clk), .D (new_AGEMA_signal_3042), .Q (new_AGEMA_signal_5031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2513 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T4), .Q (new_AGEMA_signal_5034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2516 ( .C (clk), .D (new_AGEMA_signal_3045), .Q (new_AGEMA_signal_5037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2519 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_T2), .Q (new_AGEMA_signal_5040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2522 ( .C (clk), .D (new_AGEMA_signal_3043), .Q (new_AGEMA_signal_5043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2525 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T6), .Q (new_AGEMA_signal_5046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2528 ( .C (clk), .D (new_AGEMA_signal_3090), .Q (new_AGEMA_signal_5049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2531 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T8), .Q (new_AGEMA_signal_5052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2534 ( .C (clk), .D (new_AGEMA_signal_3127), .Q (new_AGEMA_signal_5055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2537 ( .C (clk), .D (SubBytesInput[8]), .Q (new_AGEMA_signal_5058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2540 ( .C (clk), .D (new_AGEMA_signal_2722), .Q (new_AGEMA_signal_5061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2543 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T16), .Q (new_AGEMA_signal_5064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2546 ( .C (clk), .D (new_AGEMA_signal_3094), .Q (new_AGEMA_signal_5067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2549 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T9), .Q (new_AGEMA_signal_5070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2552 ( .C (clk), .D (new_AGEMA_signal_3091), .Q (new_AGEMA_signal_5073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2555 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T17), .Q (new_AGEMA_signal_5076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2558 ( .C (clk), .D (new_AGEMA_signal_3130), .Q (new_AGEMA_signal_5079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2561 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T15), .Q (new_AGEMA_signal_5082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2564 ( .C (clk), .D (new_AGEMA_signal_3093), .Q (new_AGEMA_signal_5085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2567 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T27), .Q (new_AGEMA_signal_5088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2570 ( .C (clk), .D (new_AGEMA_signal_3097), .Q (new_AGEMA_signal_5091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2573 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T10), .Q (new_AGEMA_signal_5094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2576 ( .C (clk), .D (new_AGEMA_signal_3128), .Q (new_AGEMA_signal_5097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2579 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T13), .Q (new_AGEMA_signal_5100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2582 ( .C (clk), .D (new_AGEMA_signal_3092), .Q (new_AGEMA_signal_5103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2585 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T23), .Q (new_AGEMA_signal_5106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2588 ( .C (clk), .D (new_AGEMA_signal_3132), .Q (new_AGEMA_signal_5109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2591 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T19), .Q (new_AGEMA_signal_5112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2594 ( .C (clk), .D (new_AGEMA_signal_3095), .Q (new_AGEMA_signal_5115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2597 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T3), .Q (new_AGEMA_signal_5118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2600 ( .C (clk), .D (new_AGEMA_signal_3054), .Q (new_AGEMA_signal_5121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2603 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T22), .Q (new_AGEMA_signal_5124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2606 ( .C (clk), .D (new_AGEMA_signal_3096), .Q (new_AGEMA_signal_5127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2609 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T20), .Q (new_AGEMA_signal_5130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2612 ( .C (clk), .D (new_AGEMA_signal_3131), .Q (new_AGEMA_signal_5133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2615 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T1), .Q (new_AGEMA_signal_5136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2618 ( .C (clk), .D (new_AGEMA_signal_3052), .Q (new_AGEMA_signal_5139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2621 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T4), .Q (new_AGEMA_signal_5142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2624 ( .C (clk), .D (new_AGEMA_signal_3055), .Q (new_AGEMA_signal_5145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2627 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_T2), .Q (new_AGEMA_signal_5148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2630 ( .C (clk), .D (new_AGEMA_signal_3053), .Q (new_AGEMA_signal_5151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2633 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T6), .Q (new_AGEMA_signal_5154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2636 ( .C (clk), .D (new_AGEMA_signal_3098), .Q (new_AGEMA_signal_5157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2639 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T8), .Q (new_AGEMA_signal_5160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2642 ( .C (clk), .D (new_AGEMA_signal_3140), .Q (new_AGEMA_signal_5163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2645 ( .C (clk), .D (SubBytesInput[16]), .Q (new_AGEMA_signal_5166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2648 ( .C (clk), .D (new_AGEMA_signal_2738), .Q (new_AGEMA_signal_5169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2651 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T16), .Q (new_AGEMA_signal_5172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2654 ( .C (clk), .D (new_AGEMA_signal_3102), .Q (new_AGEMA_signal_5175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2657 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T9), .Q (new_AGEMA_signal_5178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2660 ( .C (clk), .D (new_AGEMA_signal_3099), .Q (new_AGEMA_signal_5181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2663 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T17), .Q (new_AGEMA_signal_5184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2666 ( .C (clk), .D (new_AGEMA_signal_3143), .Q (new_AGEMA_signal_5187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2669 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T15), .Q (new_AGEMA_signal_5190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2672 ( .C (clk), .D (new_AGEMA_signal_3101), .Q (new_AGEMA_signal_5193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2675 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T27), .Q (new_AGEMA_signal_5196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2678 ( .C (clk), .D (new_AGEMA_signal_3105), .Q (new_AGEMA_signal_5199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2681 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T10), .Q (new_AGEMA_signal_5202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2684 ( .C (clk), .D (new_AGEMA_signal_3141), .Q (new_AGEMA_signal_5205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2687 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T13), .Q (new_AGEMA_signal_5208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2690 ( .C (clk), .D (new_AGEMA_signal_3100), .Q (new_AGEMA_signal_5211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2693 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T23), .Q (new_AGEMA_signal_5214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2696 ( .C (clk), .D (new_AGEMA_signal_3145), .Q (new_AGEMA_signal_5217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2699 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T19), .Q (new_AGEMA_signal_5220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2702 ( .C (clk), .D (new_AGEMA_signal_3103), .Q (new_AGEMA_signal_5223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2705 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T3), .Q (new_AGEMA_signal_5226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2708 ( .C (clk), .D (new_AGEMA_signal_3064), .Q (new_AGEMA_signal_5229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2711 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T22), .Q (new_AGEMA_signal_5232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2714 ( .C (clk), .D (new_AGEMA_signal_3104), .Q (new_AGEMA_signal_5235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2717 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T20), .Q (new_AGEMA_signal_5238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2720 ( .C (clk), .D (new_AGEMA_signal_3144), .Q (new_AGEMA_signal_5241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2723 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T1), .Q (new_AGEMA_signal_5244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2726 ( .C (clk), .D (new_AGEMA_signal_3062), .Q (new_AGEMA_signal_5247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2729 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T4), .Q (new_AGEMA_signal_5250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2732 ( .C (clk), .D (new_AGEMA_signal_3065), .Q (new_AGEMA_signal_5253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2735 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_T2), .Q (new_AGEMA_signal_5256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2738 ( .C (clk), .D (new_AGEMA_signal_3063), .Q (new_AGEMA_signal_5259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2741 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T6), .Q (new_AGEMA_signal_5262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2744 ( .C (clk), .D (new_AGEMA_signal_3106), .Q (new_AGEMA_signal_5265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2747 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T8), .Q (new_AGEMA_signal_5268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2750 ( .C (clk), .D (new_AGEMA_signal_3153), .Q (new_AGEMA_signal_5271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2753 ( .C (clk), .D (SubBytesInput[24]), .Q (new_AGEMA_signal_5274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2756 ( .C (clk), .D (new_AGEMA_signal_2746), .Q (new_AGEMA_signal_5277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2759 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T16), .Q (new_AGEMA_signal_5280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2762 ( .C (clk), .D (new_AGEMA_signal_3110), .Q (new_AGEMA_signal_5283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2765 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T9), .Q (new_AGEMA_signal_5286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2768 ( .C (clk), .D (new_AGEMA_signal_3107), .Q (new_AGEMA_signal_5289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2771 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T17), .Q (new_AGEMA_signal_5292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2774 ( .C (clk), .D (new_AGEMA_signal_3156), .Q (new_AGEMA_signal_5295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2777 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T15), .Q (new_AGEMA_signal_5298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2780 ( .C (clk), .D (new_AGEMA_signal_3109), .Q (new_AGEMA_signal_5301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2783 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T27), .Q (new_AGEMA_signal_5304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2786 ( .C (clk), .D (new_AGEMA_signal_3113), .Q (new_AGEMA_signal_5307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2789 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T10), .Q (new_AGEMA_signal_5310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2792 ( .C (clk), .D (new_AGEMA_signal_3154), .Q (new_AGEMA_signal_5313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2795 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T13), .Q (new_AGEMA_signal_5316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2798 ( .C (clk), .D (new_AGEMA_signal_3108), .Q (new_AGEMA_signal_5319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2801 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T23), .Q (new_AGEMA_signal_5322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2804 ( .C (clk), .D (new_AGEMA_signal_3158), .Q (new_AGEMA_signal_5325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2807 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T19), .Q (new_AGEMA_signal_5328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2810 ( .C (clk), .D (new_AGEMA_signal_3111), .Q (new_AGEMA_signal_5331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2813 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T3), .Q (new_AGEMA_signal_5334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2816 ( .C (clk), .D (new_AGEMA_signal_3074), .Q (new_AGEMA_signal_5337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2819 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T22), .Q (new_AGEMA_signal_5340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2822 ( .C (clk), .D (new_AGEMA_signal_3112), .Q (new_AGEMA_signal_5343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2825 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T20), .Q (new_AGEMA_signal_5346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2828 ( .C (clk), .D (new_AGEMA_signal_3157), .Q (new_AGEMA_signal_5349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2831 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T1), .Q (new_AGEMA_signal_5352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2834 ( .C (clk), .D (new_AGEMA_signal_3072), .Q (new_AGEMA_signal_5355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2837 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T4), .Q (new_AGEMA_signal_5358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2840 ( .C (clk), .D (new_AGEMA_signal_3075), .Q (new_AGEMA_signal_5361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2843 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_T2), .Q (new_AGEMA_signal_5364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2846 ( .C (clk), .D (new_AGEMA_signal_3073), .Q (new_AGEMA_signal_5367) ) ;
    buf_clk new_AGEMA_reg_buffer_2849 ( .C (clk), .D (MuxMCOut_n5), .Q (new_AGEMA_signal_5370) ) ;
    buf_clk new_AGEMA_reg_buffer_2853 ( .C (clk), .D (LastRoundorDone), .Q (new_AGEMA_signal_5374) ) ;
    buf_clk new_AGEMA_reg_buffer_2857 ( .C (clk), .D (MuxMCOut_n4), .Q (new_AGEMA_signal_5378) ) ;
    buf_clk new_AGEMA_reg_buffer_2861 ( .C (clk), .D (AKSRnotDone), .Q (new_AGEMA_signal_5382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2865 ( .C (clk), .D (ShiftRowsOutput[0]), .Q (new_AGEMA_signal_5386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2869 ( .C (clk), .D (new_AGEMA_signal_2499), .Q (new_AGEMA_signal_5390) ) ;
    buf_clk new_AGEMA_reg_buffer_2873 ( .C (clk), .D (MuxRound_n13), .Q (new_AGEMA_signal_5394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2877 ( .C (clk), .D (ShiftRowsOutput[1]), .Q (new_AGEMA_signal_5398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2881 ( .C (clk), .D (new_AGEMA_signal_2502), .Q (new_AGEMA_signal_5402) ) ;
    buf_clk new_AGEMA_reg_buffer_2885 ( .C (clk), .D (MuxRound_n14), .Q (new_AGEMA_signal_5406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2889 ( .C (clk), .D (ShiftRowsOutput[2]), .Q (new_AGEMA_signal_5410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2893 ( .C (clk), .D (new_AGEMA_signal_2505), .Q (new_AGEMA_signal_5414) ) ;
    buf_clk new_AGEMA_reg_buffer_2897 ( .C (clk), .D (MuxRound_n15), .Q (new_AGEMA_signal_5418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2901 ( .C (clk), .D (ShiftRowsOutput[3]), .Q (new_AGEMA_signal_5422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2905 ( .C (clk), .D (new_AGEMA_signal_2508), .Q (new_AGEMA_signal_5426) ) ;
    buf_clk new_AGEMA_reg_buffer_2909 ( .C (clk), .D (MuxRound_n16), .Q (new_AGEMA_signal_5430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2913 ( .C (clk), .D (ShiftRowsOutput[4]), .Q (new_AGEMA_signal_5434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2917 ( .C (clk), .D (new_AGEMA_signal_2511), .Q (new_AGEMA_signal_5438) ) ;
    buf_clk new_AGEMA_reg_buffer_2921 ( .C (clk), .D (MuxRound_n17), .Q (new_AGEMA_signal_5442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2925 ( .C (clk), .D (ShiftRowsOutput[5]), .Q (new_AGEMA_signal_5446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2929 ( .C (clk), .D (new_AGEMA_signal_2514), .Q (new_AGEMA_signal_5450) ) ;
    buf_clk new_AGEMA_reg_buffer_2933 ( .C (clk), .D (MuxRound_n18), .Q (new_AGEMA_signal_5454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2937 ( .C (clk), .D (ShiftRowsOutput[6]), .Q (new_AGEMA_signal_5458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2941 ( .C (clk), .D (new_AGEMA_signal_2517), .Q (new_AGEMA_signal_5462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2945 ( .C (clk), .D (ShiftRowsOutput[7]), .Q (new_AGEMA_signal_5466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2949 ( .C (clk), .D (new_AGEMA_signal_2520), .Q (new_AGEMA_signal_5470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2953 ( .C (clk), .D (ShiftRowsOutput[8]), .Q (new_AGEMA_signal_5474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2957 ( .C (clk), .D (new_AGEMA_signal_2631), .Q (new_AGEMA_signal_5478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2961 ( .C (clk), .D (ShiftRowsOutput[9]), .Q (new_AGEMA_signal_5482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2965 ( .C (clk), .D (new_AGEMA_signal_2634), .Q (new_AGEMA_signal_5486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2969 ( .C (clk), .D (ShiftRowsOutput[10]), .Q (new_AGEMA_signal_5490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2973 ( .C (clk), .D (new_AGEMA_signal_2637), .Q (new_AGEMA_signal_5494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2977 ( .C (clk), .D (ShiftRowsOutput[11]), .Q (new_AGEMA_signal_5498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2981 ( .C (clk), .D (new_AGEMA_signal_2640), .Q (new_AGEMA_signal_5502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2985 ( .C (clk), .D (ShiftRowsOutput[12]), .Q (new_AGEMA_signal_5506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2989 ( .C (clk), .D (new_AGEMA_signal_2643), .Q (new_AGEMA_signal_5510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2993 ( .C (clk), .D (ShiftRowsOutput[13]), .Q (new_AGEMA_signal_5514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2997 ( .C (clk), .D (new_AGEMA_signal_2646), .Q (new_AGEMA_signal_5518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3001 ( .C (clk), .D (ShiftRowsOutput[14]), .Q (new_AGEMA_signal_5522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3005 ( .C (clk), .D (new_AGEMA_signal_2649), .Q (new_AGEMA_signal_5526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3009 ( .C (clk), .D (ShiftRowsOutput[15]), .Q (new_AGEMA_signal_5530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3013 ( .C (clk), .D (new_AGEMA_signal_2652), .Q (new_AGEMA_signal_5534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3017 ( .C (clk), .D (ShiftRowsOutput[16]), .Q (new_AGEMA_signal_5538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3021 ( .C (clk), .D (new_AGEMA_signal_2382), .Q (new_AGEMA_signal_5542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3025 ( .C (clk), .D (ShiftRowsOutput[17]), .Q (new_AGEMA_signal_5546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3029 ( .C (clk), .D (new_AGEMA_signal_2385), .Q (new_AGEMA_signal_5550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3033 ( .C (clk), .D (ShiftRowsOutput[18]), .Q (new_AGEMA_signal_5554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3037 ( .C (clk), .D (new_AGEMA_signal_2388), .Q (new_AGEMA_signal_5558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3041 ( .C (clk), .D (ShiftRowsOutput[19]), .Q (new_AGEMA_signal_5562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3045 ( .C (clk), .D (new_AGEMA_signal_2391), .Q (new_AGEMA_signal_5566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3049 ( .C (clk), .D (ShiftRowsOutput[20]), .Q (new_AGEMA_signal_5570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3053 ( .C (clk), .D (new_AGEMA_signal_2394), .Q (new_AGEMA_signal_5574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3057 ( .C (clk), .D (ShiftRowsOutput[21]), .Q (new_AGEMA_signal_5578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3061 ( .C (clk), .D (new_AGEMA_signal_2397), .Q (new_AGEMA_signal_5582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3065 ( .C (clk), .D (ShiftRowsOutput[22]), .Q (new_AGEMA_signal_5586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3069 ( .C (clk), .D (new_AGEMA_signal_2400), .Q (new_AGEMA_signal_5590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3073 ( .C (clk), .D (ShiftRowsOutput[23]), .Q (new_AGEMA_signal_5594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3077 ( .C (clk), .D (new_AGEMA_signal_2403), .Q (new_AGEMA_signal_5598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3081 ( .C (clk), .D (ShiftRowsOutput[24]), .Q (new_AGEMA_signal_5602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3085 ( .C (clk), .D (new_AGEMA_signal_2472), .Q (new_AGEMA_signal_5606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3089 ( .C (clk), .D (ShiftRowsOutput[25]), .Q (new_AGEMA_signal_5610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3093 ( .C (clk), .D (new_AGEMA_signal_2475), .Q (new_AGEMA_signal_5614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3097 ( .C (clk), .D (ShiftRowsOutput[26]), .Q (new_AGEMA_signal_5618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3101 ( .C (clk), .D (new_AGEMA_signal_2478), .Q (new_AGEMA_signal_5622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3105 ( .C (clk), .D (ShiftRowsOutput[27]), .Q (new_AGEMA_signal_5626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3109 ( .C (clk), .D (new_AGEMA_signal_2481), .Q (new_AGEMA_signal_5630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3113 ( .C (clk), .D (ShiftRowsOutput[28]), .Q (new_AGEMA_signal_5634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3117 ( .C (clk), .D (new_AGEMA_signal_2484), .Q (new_AGEMA_signal_5638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3121 ( .C (clk), .D (ShiftRowsOutput[29]), .Q (new_AGEMA_signal_5642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3125 ( .C (clk), .D (new_AGEMA_signal_2487), .Q (new_AGEMA_signal_5646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3129 ( .C (clk), .D (ShiftRowsOutput[30]), .Q (new_AGEMA_signal_5650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3133 ( .C (clk), .D (new_AGEMA_signal_2493), .Q (new_AGEMA_signal_5654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3137 ( .C (clk), .D (ShiftRowsOutput[31]), .Q (new_AGEMA_signal_5658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3141 ( .C (clk), .D (new_AGEMA_signal_2496), .Q (new_AGEMA_signal_5662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3145 ( .C (clk), .D (key_s0[0]), .Q (new_AGEMA_signal_5666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3149 ( .C (clk), .D (key_s1[0]), .Q (new_AGEMA_signal_5670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3153 ( .C (clk), .D (key_s0[1]), .Q (new_AGEMA_signal_5674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3157 ( .C (clk), .D (key_s1[1]), .Q (new_AGEMA_signal_5678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3161 ( .C (clk), .D (key_s0[2]), .Q (new_AGEMA_signal_5682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3165 ( .C (clk), .D (key_s1[2]), .Q (new_AGEMA_signal_5686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3169 ( .C (clk), .D (key_s0[3]), .Q (new_AGEMA_signal_5690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3173 ( .C (clk), .D (key_s1[3]), .Q (new_AGEMA_signal_5694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3177 ( .C (clk), .D (key_s0[4]), .Q (new_AGEMA_signal_5698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3181 ( .C (clk), .D (key_s1[4]), .Q (new_AGEMA_signal_5702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3185 ( .C (clk), .D (key_s0[5]), .Q (new_AGEMA_signal_5706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3189 ( .C (clk), .D (key_s1[5]), .Q (new_AGEMA_signal_5710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3193 ( .C (clk), .D (key_s0[6]), .Q (new_AGEMA_signal_5714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3197 ( .C (clk), .D (key_s1[6]), .Q (new_AGEMA_signal_5718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3201 ( .C (clk), .D (key_s0[7]), .Q (new_AGEMA_signal_5722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3205 ( .C (clk), .D (key_s1[7]), .Q (new_AGEMA_signal_5726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3209 ( .C (clk), .D (key_s0[8]), .Q (new_AGEMA_signal_5730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3213 ( .C (clk), .D (key_s1[8]), .Q (new_AGEMA_signal_5734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3217 ( .C (clk), .D (key_s0[9]), .Q (new_AGEMA_signal_5738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3221 ( .C (clk), .D (key_s1[9]), .Q (new_AGEMA_signal_5742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3225 ( .C (clk), .D (key_s0[10]), .Q (new_AGEMA_signal_5746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3229 ( .C (clk), .D (key_s1[10]), .Q (new_AGEMA_signal_5750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3233 ( .C (clk), .D (key_s0[11]), .Q (new_AGEMA_signal_5754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3237 ( .C (clk), .D (key_s1[11]), .Q (new_AGEMA_signal_5758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3241 ( .C (clk), .D (key_s0[12]), .Q (new_AGEMA_signal_5762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3245 ( .C (clk), .D (key_s1[12]), .Q (new_AGEMA_signal_5766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3249 ( .C (clk), .D (key_s0[13]), .Q (new_AGEMA_signal_5770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3253 ( .C (clk), .D (key_s1[13]), .Q (new_AGEMA_signal_5774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3257 ( .C (clk), .D (key_s0[14]), .Q (new_AGEMA_signal_5778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3261 ( .C (clk), .D (key_s1[14]), .Q (new_AGEMA_signal_5782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3265 ( .C (clk), .D (key_s0[15]), .Q (new_AGEMA_signal_5786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3269 ( .C (clk), .D (key_s1[15]), .Q (new_AGEMA_signal_5790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3273 ( .C (clk), .D (key_s0[16]), .Q (new_AGEMA_signal_5794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3277 ( .C (clk), .D (key_s1[16]), .Q (new_AGEMA_signal_5798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3281 ( .C (clk), .D (key_s0[17]), .Q (new_AGEMA_signal_5802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3285 ( .C (clk), .D (key_s1[17]), .Q (new_AGEMA_signal_5806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3289 ( .C (clk), .D (key_s0[18]), .Q (new_AGEMA_signal_5810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3293 ( .C (clk), .D (key_s1[18]), .Q (new_AGEMA_signal_5814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3297 ( .C (clk), .D (key_s0[19]), .Q (new_AGEMA_signal_5818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3301 ( .C (clk), .D (key_s1[19]), .Q (new_AGEMA_signal_5822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3305 ( .C (clk), .D (key_s0[20]), .Q (new_AGEMA_signal_5826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3309 ( .C (clk), .D (key_s1[20]), .Q (new_AGEMA_signal_5830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3313 ( .C (clk), .D (key_s0[21]), .Q (new_AGEMA_signal_5834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3317 ( .C (clk), .D (key_s1[21]), .Q (new_AGEMA_signal_5838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3321 ( .C (clk), .D (key_s0[22]), .Q (new_AGEMA_signal_5842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3325 ( .C (clk), .D (key_s1[22]), .Q (new_AGEMA_signal_5846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3329 ( .C (clk), .D (key_s0[23]), .Q (new_AGEMA_signal_5850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3333 ( .C (clk), .D (key_s1[23]), .Q (new_AGEMA_signal_5854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3337 ( .C (clk), .D (key_s0[24]), .Q (new_AGEMA_signal_5858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3341 ( .C (clk), .D (key_s1[24]), .Q (new_AGEMA_signal_5862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3345 ( .C (clk), .D (key_s0[25]), .Q (new_AGEMA_signal_5866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3349 ( .C (clk), .D (key_s1[25]), .Q (new_AGEMA_signal_5870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3353 ( .C (clk), .D (key_s0[26]), .Q (new_AGEMA_signal_5874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3357 ( .C (clk), .D (key_s1[26]), .Q (new_AGEMA_signal_5878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3361 ( .C (clk), .D (key_s0[27]), .Q (new_AGEMA_signal_5882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3365 ( .C (clk), .D (key_s1[27]), .Q (new_AGEMA_signal_5886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3369 ( .C (clk), .D (key_s0[28]), .Q (new_AGEMA_signal_5890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3373 ( .C (clk), .D (key_s1[28]), .Q (new_AGEMA_signal_5894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3377 ( .C (clk), .D (key_s0[29]), .Q (new_AGEMA_signal_5898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3381 ( .C (clk), .D (key_s1[29]), .Q (new_AGEMA_signal_5902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3385 ( .C (clk), .D (key_s0[30]), .Q (new_AGEMA_signal_5906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3389 ( .C (clk), .D (key_s1[30]), .Q (new_AGEMA_signal_5910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3393 ( .C (clk), .D (key_s0[31]), .Q (new_AGEMA_signal_5914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3397 ( .C (clk), .D (key_s1[31]), .Q (new_AGEMA_signal_5918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3401 ( .C (clk), .D (key_s0[32]), .Q (new_AGEMA_signal_5922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3405 ( .C (clk), .D (key_s1[32]), .Q (new_AGEMA_signal_5926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3409 ( .C (clk), .D (key_s0[33]), .Q (new_AGEMA_signal_5930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3413 ( .C (clk), .D (key_s1[33]), .Q (new_AGEMA_signal_5934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3417 ( .C (clk), .D (key_s0[34]), .Q (new_AGEMA_signal_5938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3421 ( .C (clk), .D (key_s1[34]), .Q (new_AGEMA_signal_5942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3425 ( .C (clk), .D (key_s0[35]), .Q (new_AGEMA_signal_5946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3429 ( .C (clk), .D (key_s1[35]), .Q (new_AGEMA_signal_5950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3433 ( .C (clk), .D (key_s0[36]), .Q (new_AGEMA_signal_5954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3437 ( .C (clk), .D (key_s1[36]), .Q (new_AGEMA_signal_5958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3441 ( .C (clk), .D (key_s0[37]), .Q (new_AGEMA_signal_5962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3445 ( .C (clk), .D (key_s1[37]), .Q (new_AGEMA_signal_5966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3449 ( .C (clk), .D (key_s0[38]), .Q (new_AGEMA_signal_5970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3453 ( .C (clk), .D (key_s1[38]), .Q (new_AGEMA_signal_5974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3457 ( .C (clk), .D (key_s0[39]), .Q (new_AGEMA_signal_5978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3461 ( .C (clk), .D (key_s1[39]), .Q (new_AGEMA_signal_5982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3465 ( .C (clk), .D (key_s0[40]), .Q (new_AGEMA_signal_5986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3469 ( .C (clk), .D (key_s1[40]), .Q (new_AGEMA_signal_5990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3473 ( .C (clk), .D (key_s0[41]), .Q (new_AGEMA_signal_5994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3477 ( .C (clk), .D (key_s1[41]), .Q (new_AGEMA_signal_5998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3481 ( .C (clk), .D (key_s0[42]), .Q (new_AGEMA_signal_6002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3485 ( .C (clk), .D (key_s1[42]), .Q (new_AGEMA_signal_6006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3489 ( .C (clk), .D (key_s0[43]), .Q (new_AGEMA_signal_6010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3493 ( .C (clk), .D (key_s1[43]), .Q (new_AGEMA_signal_6014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3497 ( .C (clk), .D (key_s0[44]), .Q (new_AGEMA_signal_6018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3501 ( .C (clk), .D (key_s1[44]), .Q (new_AGEMA_signal_6022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3505 ( .C (clk), .D (key_s0[45]), .Q (new_AGEMA_signal_6026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3509 ( .C (clk), .D (key_s1[45]), .Q (new_AGEMA_signal_6030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3513 ( .C (clk), .D (key_s0[46]), .Q (new_AGEMA_signal_6034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3517 ( .C (clk), .D (key_s1[46]), .Q (new_AGEMA_signal_6038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3521 ( .C (clk), .D (key_s0[47]), .Q (new_AGEMA_signal_6042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3525 ( .C (clk), .D (key_s1[47]), .Q (new_AGEMA_signal_6046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3529 ( .C (clk), .D (key_s0[48]), .Q (new_AGEMA_signal_6050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3533 ( .C (clk), .D (key_s1[48]), .Q (new_AGEMA_signal_6054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3537 ( .C (clk), .D (key_s0[49]), .Q (new_AGEMA_signal_6058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3541 ( .C (clk), .D (key_s1[49]), .Q (new_AGEMA_signal_6062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3545 ( .C (clk), .D (key_s0[50]), .Q (new_AGEMA_signal_6066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3549 ( .C (clk), .D (key_s1[50]), .Q (new_AGEMA_signal_6070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3553 ( .C (clk), .D (key_s0[51]), .Q (new_AGEMA_signal_6074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3557 ( .C (clk), .D (key_s1[51]), .Q (new_AGEMA_signal_6078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3561 ( .C (clk), .D (key_s0[52]), .Q (new_AGEMA_signal_6082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3565 ( .C (clk), .D (key_s1[52]), .Q (new_AGEMA_signal_6086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3569 ( .C (clk), .D (key_s0[53]), .Q (new_AGEMA_signal_6090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3573 ( .C (clk), .D (key_s1[53]), .Q (new_AGEMA_signal_6094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3577 ( .C (clk), .D (key_s0[54]), .Q (new_AGEMA_signal_6098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3581 ( .C (clk), .D (key_s1[54]), .Q (new_AGEMA_signal_6102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3585 ( .C (clk), .D (key_s0[55]), .Q (new_AGEMA_signal_6106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3589 ( .C (clk), .D (key_s1[55]), .Q (new_AGEMA_signal_6110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3593 ( .C (clk), .D (key_s0[56]), .Q (new_AGEMA_signal_6114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3597 ( .C (clk), .D (key_s1[56]), .Q (new_AGEMA_signal_6118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3601 ( .C (clk), .D (key_s0[57]), .Q (new_AGEMA_signal_6122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3605 ( .C (clk), .D (key_s1[57]), .Q (new_AGEMA_signal_6126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3609 ( .C (clk), .D (key_s0[58]), .Q (new_AGEMA_signal_6130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3613 ( .C (clk), .D (key_s1[58]), .Q (new_AGEMA_signal_6134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3617 ( .C (clk), .D (key_s0[59]), .Q (new_AGEMA_signal_6138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3621 ( .C (clk), .D (key_s1[59]), .Q (new_AGEMA_signal_6142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3625 ( .C (clk), .D (key_s0[60]), .Q (new_AGEMA_signal_6146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3629 ( .C (clk), .D (key_s1[60]), .Q (new_AGEMA_signal_6150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3633 ( .C (clk), .D (key_s0[61]), .Q (new_AGEMA_signal_6154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3637 ( .C (clk), .D (key_s1[61]), .Q (new_AGEMA_signal_6158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3641 ( .C (clk), .D (key_s0[62]), .Q (new_AGEMA_signal_6162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3645 ( .C (clk), .D (key_s1[62]), .Q (new_AGEMA_signal_6166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3649 ( .C (clk), .D (key_s0[63]), .Q (new_AGEMA_signal_6170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3653 ( .C (clk), .D (key_s1[63]), .Q (new_AGEMA_signal_6174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3657 ( .C (clk), .D (key_s0[64]), .Q (new_AGEMA_signal_6178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3661 ( .C (clk), .D (key_s1[64]), .Q (new_AGEMA_signal_6182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3665 ( .C (clk), .D (key_s0[65]), .Q (new_AGEMA_signal_6186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3669 ( .C (clk), .D (key_s1[65]), .Q (new_AGEMA_signal_6190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3673 ( .C (clk), .D (key_s0[66]), .Q (new_AGEMA_signal_6194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3677 ( .C (clk), .D (key_s1[66]), .Q (new_AGEMA_signal_6198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3681 ( .C (clk), .D (key_s0[67]), .Q (new_AGEMA_signal_6202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3685 ( .C (clk), .D (key_s1[67]), .Q (new_AGEMA_signal_6206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3689 ( .C (clk), .D (key_s0[68]), .Q (new_AGEMA_signal_6210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3693 ( .C (clk), .D (key_s1[68]), .Q (new_AGEMA_signal_6214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3697 ( .C (clk), .D (key_s0[69]), .Q (new_AGEMA_signal_6218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3701 ( .C (clk), .D (key_s1[69]), .Q (new_AGEMA_signal_6222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3705 ( .C (clk), .D (key_s0[70]), .Q (new_AGEMA_signal_6226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3709 ( .C (clk), .D (key_s1[70]), .Q (new_AGEMA_signal_6230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3713 ( .C (clk), .D (key_s0[71]), .Q (new_AGEMA_signal_6234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3717 ( .C (clk), .D (key_s1[71]), .Q (new_AGEMA_signal_6238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3721 ( .C (clk), .D (key_s0[72]), .Q (new_AGEMA_signal_6242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3725 ( .C (clk), .D (key_s1[72]), .Q (new_AGEMA_signal_6246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3729 ( .C (clk), .D (key_s0[73]), .Q (new_AGEMA_signal_6250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3733 ( .C (clk), .D (key_s1[73]), .Q (new_AGEMA_signal_6254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3737 ( .C (clk), .D (key_s0[74]), .Q (new_AGEMA_signal_6258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3741 ( .C (clk), .D (key_s1[74]), .Q (new_AGEMA_signal_6262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3745 ( .C (clk), .D (key_s0[75]), .Q (new_AGEMA_signal_6266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3749 ( .C (clk), .D (key_s1[75]), .Q (new_AGEMA_signal_6270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3753 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_6274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3757 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_6278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3761 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_6282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3765 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_6286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3769 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_6290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3773 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_6294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3777 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_6298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3781 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_6302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3785 ( .C (clk), .D (key_s0[80]), .Q (new_AGEMA_signal_6306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3789 ( .C (clk), .D (key_s1[80]), .Q (new_AGEMA_signal_6310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3793 ( .C (clk), .D (key_s0[81]), .Q (new_AGEMA_signal_6314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3797 ( .C (clk), .D (key_s1[81]), .Q (new_AGEMA_signal_6318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3801 ( .C (clk), .D (key_s0[82]), .Q (new_AGEMA_signal_6322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3805 ( .C (clk), .D (key_s1[82]), .Q (new_AGEMA_signal_6326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3809 ( .C (clk), .D (key_s0[83]), .Q (new_AGEMA_signal_6330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3813 ( .C (clk), .D (key_s1[83]), .Q (new_AGEMA_signal_6334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3817 ( .C (clk), .D (key_s0[84]), .Q (new_AGEMA_signal_6338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3821 ( .C (clk), .D (key_s1[84]), .Q (new_AGEMA_signal_6342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3825 ( .C (clk), .D (key_s0[85]), .Q (new_AGEMA_signal_6346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3829 ( .C (clk), .D (key_s1[85]), .Q (new_AGEMA_signal_6350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3833 ( .C (clk), .D (key_s0[86]), .Q (new_AGEMA_signal_6354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3837 ( .C (clk), .D (key_s1[86]), .Q (new_AGEMA_signal_6358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3841 ( .C (clk), .D (key_s0[87]), .Q (new_AGEMA_signal_6362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3845 ( .C (clk), .D (key_s1[87]), .Q (new_AGEMA_signal_6366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3849 ( .C (clk), .D (key_s0[88]), .Q (new_AGEMA_signal_6370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3853 ( .C (clk), .D (key_s1[88]), .Q (new_AGEMA_signal_6374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3857 ( .C (clk), .D (key_s0[89]), .Q (new_AGEMA_signal_6378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3861 ( .C (clk), .D (key_s1[89]), .Q (new_AGEMA_signal_6382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3865 ( .C (clk), .D (key_s0[90]), .Q (new_AGEMA_signal_6386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3869 ( .C (clk), .D (key_s1[90]), .Q (new_AGEMA_signal_6390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3873 ( .C (clk), .D (key_s0[91]), .Q (new_AGEMA_signal_6394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3877 ( .C (clk), .D (key_s1[91]), .Q (new_AGEMA_signal_6398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3881 ( .C (clk), .D (key_s0[92]), .Q (new_AGEMA_signal_6402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3885 ( .C (clk), .D (key_s1[92]), .Q (new_AGEMA_signal_6406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3889 ( .C (clk), .D (key_s0[93]), .Q (new_AGEMA_signal_6410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3893 ( .C (clk), .D (key_s1[93]), .Q (new_AGEMA_signal_6414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3897 ( .C (clk), .D (key_s0[94]), .Q (new_AGEMA_signal_6418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3901 ( .C (clk), .D (key_s1[94]), .Q (new_AGEMA_signal_6422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3905 ( .C (clk), .D (key_s0[95]), .Q (new_AGEMA_signal_6426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3909 ( .C (clk), .D (key_s1[95]), .Q (new_AGEMA_signal_6430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3913 ( .C (clk), .D (key_s0[96]), .Q (new_AGEMA_signal_6434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3917 ( .C (clk), .D (key_s1[96]), .Q (new_AGEMA_signal_6438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3921 ( .C (clk), .D (key_s0[97]), .Q (new_AGEMA_signal_6442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3925 ( .C (clk), .D (key_s1[97]), .Q (new_AGEMA_signal_6446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3929 ( .C (clk), .D (key_s0[98]), .Q (new_AGEMA_signal_6450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3933 ( .C (clk), .D (key_s1[98]), .Q (new_AGEMA_signal_6454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3937 ( .C (clk), .D (key_s0[99]), .Q (new_AGEMA_signal_6458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3941 ( .C (clk), .D (key_s1[99]), .Q (new_AGEMA_signal_6462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3945 ( .C (clk), .D (key_s0[100]), .Q (new_AGEMA_signal_6466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3949 ( .C (clk), .D (key_s1[100]), .Q (new_AGEMA_signal_6470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3953 ( .C (clk), .D (key_s0[101]), .Q (new_AGEMA_signal_6474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3957 ( .C (clk), .D (key_s1[101]), .Q (new_AGEMA_signal_6478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3961 ( .C (clk), .D (key_s0[102]), .Q (new_AGEMA_signal_6482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3965 ( .C (clk), .D (key_s1[102]), .Q (new_AGEMA_signal_6486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3969 ( .C (clk), .D (key_s0[103]), .Q (new_AGEMA_signal_6490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3973 ( .C (clk), .D (key_s1[103]), .Q (new_AGEMA_signal_6494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3977 ( .C (clk), .D (key_s0[104]), .Q (new_AGEMA_signal_6498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3981 ( .C (clk), .D (key_s1[104]), .Q (new_AGEMA_signal_6502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3985 ( .C (clk), .D (key_s0[105]), .Q (new_AGEMA_signal_6506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3989 ( .C (clk), .D (key_s1[105]), .Q (new_AGEMA_signal_6510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3993 ( .C (clk), .D (key_s0[106]), .Q (new_AGEMA_signal_6514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3997 ( .C (clk), .D (key_s1[106]), .Q (new_AGEMA_signal_6518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4001 ( .C (clk), .D (key_s0[107]), .Q (new_AGEMA_signal_6522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4005 ( .C (clk), .D (key_s1[107]), .Q (new_AGEMA_signal_6526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4009 ( .C (clk), .D (key_s0[108]), .Q (new_AGEMA_signal_6530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4013 ( .C (clk), .D (key_s1[108]), .Q (new_AGEMA_signal_6534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4017 ( .C (clk), .D (key_s0[109]), .Q (new_AGEMA_signal_6538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4021 ( .C (clk), .D (key_s1[109]), .Q (new_AGEMA_signal_6542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4025 ( .C (clk), .D (key_s0[110]), .Q (new_AGEMA_signal_6546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4029 ( .C (clk), .D (key_s1[110]), .Q (new_AGEMA_signal_6550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4033 ( .C (clk), .D (key_s0[111]), .Q (new_AGEMA_signal_6554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4037 ( .C (clk), .D (key_s1[111]), .Q (new_AGEMA_signal_6558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4041 ( .C (clk), .D (key_s0[112]), .Q (new_AGEMA_signal_6562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4045 ( .C (clk), .D (key_s1[112]), .Q (new_AGEMA_signal_6566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4049 ( .C (clk), .D (key_s0[113]), .Q (new_AGEMA_signal_6570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4053 ( .C (clk), .D (key_s1[113]), .Q (new_AGEMA_signal_6574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4057 ( .C (clk), .D (key_s0[114]), .Q (new_AGEMA_signal_6578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4061 ( .C (clk), .D (key_s1[114]), .Q (new_AGEMA_signal_6582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4065 ( .C (clk), .D (key_s0[115]), .Q (new_AGEMA_signal_6586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4069 ( .C (clk), .D (key_s1[115]), .Q (new_AGEMA_signal_6590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4073 ( .C (clk), .D (key_s0[116]), .Q (new_AGEMA_signal_6594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4077 ( .C (clk), .D (key_s1[116]), .Q (new_AGEMA_signal_6598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4081 ( .C (clk), .D (key_s0[117]), .Q (new_AGEMA_signal_6602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4085 ( .C (clk), .D (key_s1[117]), .Q (new_AGEMA_signal_6606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4089 ( .C (clk), .D (key_s0[118]), .Q (new_AGEMA_signal_6610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4093 ( .C (clk), .D (key_s1[118]), .Q (new_AGEMA_signal_6614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4097 ( .C (clk), .D (key_s0[119]), .Q (new_AGEMA_signal_6618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4101 ( .C (clk), .D (key_s1[119]), .Q (new_AGEMA_signal_6622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4105 ( .C (clk), .D (key_s0[120]), .Q (new_AGEMA_signal_6626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4109 ( .C (clk), .D (key_s1[120]), .Q (new_AGEMA_signal_6630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4113 ( .C (clk), .D (key_s0[121]), .Q (new_AGEMA_signal_6634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4117 ( .C (clk), .D (key_s1[121]), .Q (new_AGEMA_signal_6638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4121 ( .C (clk), .D (key_s0[122]), .Q (new_AGEMA_signal_6642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4125 ( .C (clk), .D (key_s1[122]), .Q (new_AGEMA_signal_6646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4129 ( .C (clk), .D (key_s0[123]), .Q (new_AGEMA_signal_6650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4133 ( .C (clk), .D (key_s1[123]), .Q (new_AGEMA_signal_6654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4137 ( .C (clk), .D (key_s0[124]), .Q (new_AGEMA_signal_6658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4141 ( .C (clk), .D (key_s1[124]), .Q (new_AGEMA_signal_6662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4145 ( .C (clk), .D (key_s0[125]), .Q (new_AGEMA_signal_6666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4149 ( .C (clk), .D (key_s1[125]), .Q (new_AGEMA_signal_6670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4153 ( .C (clk), .D (key_s0[126]), .Q (new_AGEMA_signal_6674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4157 ( .C (clk), .D (key_s1[126]), .Q (new_AGEMA_signal_6678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4161 ( .C (clk), .D (key_s0[127]), .Q (new_AGEMA_signal_6682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4165 ( .C (clk), .D (key_s1[127]), .Q (new_AGEMA_signal_6686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4169 ( .C (clk), .D (KSSubBytesInput[9]), .Q (new_AGEMA_signal_6690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4173 ( .C (clk), .D (new_AGEMA_signal_2720), .Q (new_AGEMA_signal_6694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4177 ( .C (clk), .D (KSSubBytesInput[8]), .Q (new_AGEMA_signal_6698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4181 ( .C (clk), .D (new_AGEMA_signal_2687), .Q (new_AGEMA_signal_6702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4185 ( .C (clk), .D (KSSubBytesInput[23]), .Q (new_AGEMA_signal_6706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4189 ( .C (clk), .D (new_AGEMA_signal_2654), .Q (new_AGEMA_signal_6710) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4193 ( .C (clk), .D (KSSubBytesInput[22]), .Q (new_AGEMA_signal_6714) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4197 ( .C (clk), .D (new_AGEMA_signal_2621), .Q (new_AGEMA_signal_6718) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4201 ( .C (clk), .D (KSSubBytesInput[21]), .Q (new_AGEMA_signal_6722) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4205 ( .C (clk), .D (new_AGEMA_signal_2588), .Q (new_AGEMA_signal_6726) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4209 ( .C (clk), .D (KSSubBytesInput[20]), .Q (new_AGEMA_signal_6730) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4213 ( .C (clk), .D (new_AGEMA_signal_2555), .Q (new_AGEMA_signal_6734) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4217 ( .C (clk), .D (RoundKey[41]), .Q (new_AGEMA_signal_6738) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4221 ( .C (clk), .D (new_AGEMA_signal_2528), .Q (new_AGEMA_signal_6742) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4225 ( .C (clk), .D (RoundKey[73]), .Q (new_AGEMA_signal_6746) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4229 ( .C (clk), .D (new_AGEMA_signal_2633), .Q (new_AGEMA_signal_6750) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4233 ( .C (clk), .D (RoundKey[40]), .Q (new_AGEMA_signal_6754) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4237 ( .C (clk), .D (new_AGEMA_signal_2525), .Q (new_AGEMA_signal_6758) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4241 ( .C (clk), .D (RoundKey[72]), .Q (new_AGEMA_signal_6762) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4245 ( .C (clk), .D (new_AGEMA_signal_2630), .Q (new_AGEMA_signal_6766) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4249 ( .C (clk), .D (KSSubBytesInput[19]), .Q (new_AGEMA_signal_6770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4253 ( .C (clk), .D (new_AGEMA_signal_2522), .Q (new_AGEMA_signal_6774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4257 ( .C (clk), .D (RoundKey[39]), .Q (new_AGEMA_signal_6778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4261 ( .C (clk), .D (new_AGEMA_signal_2519), .Q (new_AGEMA_signal_6782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4265 ( .C (clk), .D (RoundKey[71]), .Q (new_AGEMA_signal_6786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4269 ( .C (clk), .D (new_AGEMA_signal_2627), .Q (new_AGEMA_signal_6790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4273 ( .C (clk), .D (RoundKey[38]), .Q (new_AGEMA_signal_6794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4277 ( .C (clk), .D (new_AGEMA_signal_2516), .Q (new_AGEMA_signal_6798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4281 ( .C (clk), .D (RoundKey[70]), .Q (new_AGEMA_signal_6802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4285 ( .C (clk), .D (new_AGEMA_signal_2624), .Q (new_AGEMA_signal_6806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4289 ( .C (clk), .D (RoundKey[37]), .Q (new_AGEMA_signal_6810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4293 ( .C (clk), .D (new_AGEMA_signal_2513), .Q (new_AGEMA_signal_6814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4297 ( .C (clk), .D (RoundKey[69]), .Q (new_AGEMA_signal_6818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4301 ( .C (clk), .D (new_AGEMA_signal_2618), .Q (new_AGEMA_signal_6822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4305 ( .C (clk), .D (RoundKey[36]), .Q (new_AGEMA_signal_6826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4309 ( .C (clk), .D (new_AGEMA_signal_2510), .Q (new_AGEMA_signal_6830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4313 ( .C (clk), .D (RoundKey[68]), .Q (new_AGEMA_signal_6834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4317 ( .C (clk), .D (new_AGEMA_signal_2615), .Q (new_AGEMA_signal_6838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4321 ( .C (clk), .D (RoundKey[35]), .Q (new_AGEMA_signal_6842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4325 ( .C (clk), .D (new_AGEMA_signal_2507), .Q (new_AGEMA_signal_6846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4329 ( .C (clk), .D (RoundKey[67]), .Q (new_AGEMA_signal_6850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4333 ( .C (clk), .D (new_AGEMA_signal_2612), .Q (new_AGEMA_signal_6854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4337 ( .C (clk), .D (RoundKey[99]), .Q (new_AGEMA_signal_6858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4341 ( .C (clk), .D (new_AGEMA_signal_2717), .Q (new_AGEMA_signal_6862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4345 ( .C (clk), .D (KSSubBytesInput[31]), .Q (new_AGEMA_signal_6866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4349 ( .C (clk), .D (new_AGEMA_signal_2495), .Q (new_AGEMA_signal_6870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4353 ( .C (clk), .D (RoundKey[63]), .Q (new_AGEMA_signal_6874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4357 ( .C (clk), .D (new_AGEMA_signal_2600), .Q (new_AGEMA_signal_6878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4361 ( .C (clk), .D (RoundKey[95]), .Q (new_AGEMA_signal_6882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4365 ( .C (clk), .D (new_AGEMA_signal_2705), .Q (new_AGEMA_signal_6886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4369 ( .C (clk), .D (KSSubBytesInput[30]), .Q (new_AGEMA_signal_6890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4373 ( .C (clk), .D (new_AGEMA_signal_2492), .Q (new_AGEMA_signal_6894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4377 ( .C (clk), .D (RoundKey[62]), .Q (new_AGEMA_signal_6898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4381 ( .C (clk), .D (new_AGEMA_signal_2597), .Q (new_AGEMA_signal_6902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4385 ( .C (clk), .D (RoundKey[94]), .Q (new_AGEMA_signal_6906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4389 ( .C (clk), .D (new_AGEMA_signal_2702), .Q (new_AGEMA_signal_6910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4393 ( .C (clk), .D (KSSubBytesInput[18]), .Q (new_AGEMA_signal_6914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4397 ( .C (clk), .D (new_AGEMA_signal_2489), .Q (new_AGEMA_signal_6918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4401 ( .C (clk), .D (RoundKey[34]), .Q (new_AGEMA_signal_6922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4405 ( .C (clk), .D (new_AGEMA_signal_2504), .Q (new_AGEMA_signal_6926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4409 ( .C (clk), .D (RoundKey[66]), .Q (new_AGEMA_signal_6930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4413 ( .C (clk), .D (new_AGEMA_signal_2609), .Q (new_AGEMA_signal_6934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4417 ( .C (clk), .D (RoundKey[98]), .Q (new_AGEMA_signal_6938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4421 ( .C (clk), .D (new_AGEMA_signal_2714), .Q (new_AGEMA_signal_6942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4425 ( .C (clk), .D (KSSubBytesInput[29]), .Q (new_AGEMA_signal_6946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4429 ( .C (clk), .D (new_AGEMA_signal_2486), .Q (new_AGEMA_signal_6950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4433 ( .C (clk), .D (RoundKey[61]), .Q (new_AGEMA_signal_6954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4437 ( .C (clk), .D (new_AGEMA_signal_2594), .Q (new_AGEMA_signal_6958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4441 ( .C (clk), .D (RoundKey[93]), .Q (new_AGEMA_signal_6962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4445 ( .C (clk), .D (new_AGEMA_signal_2699), .Q (new_AGEMA_signal_6966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4449 ( .C (clk), .D (KSSubBytesInput[28]), .Q (new_AGEMA_signal_6970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4453 ( .C (clk), .D (new_AGEMA_signal_2483), .Q (new_AGEMA_signal_6974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4457 ( .C (clk), .D (RoundKey[60]), .Q (new_AGEMA_signal_6978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4461 ( .C (clk), .D (new_AGEMA_signal_2591), .Q (new_AGEMA_signal_6982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4465 ( .C (clk), .D (RoundKey[92]), .Q (new_AGEMA_signal_6986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4469 ( .C (clk), .D (new_AGEMA_signal_2696), .Q (new_AGEMA_signal_6990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4473 ( .C (clk), .D (KSSubBytesInput[27]), .Q (new_AGEMA_signal_6994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4477 ( .C (clk), .D (new_AGEMA_signal_2480), .Q (new_AGEMA_signal_6998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4481 ( .C (clk), .D (RoundKey[59]), .Q (new_AGEMA_signal_7002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4485 ( .C (clk), .D (new_AGEMA_signal_2585), .Q (new_AGEMA_signal_7006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4489 ( .C (clk), .D (RoundKey[91]), .Q (new_AGEMA_signal_7010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4493 ( .C (clk), .D (new_AGEMA_signal_2693), .Q (new_AGEMA_signal_7014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4497 ( .C (clk), .D (KSSubBytesInput[26]), .Q (new_AGEMA_signal_7018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4501 ( .C (clk), .D (new_AGEMA_signal_2477), .Q (new_AGEMA_signal_7022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4505 ( .C (clk), .D (RoundKey[58]), .Q (new_AGEMA_signal_7026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4509 ( .C (clk), .D (new_AGEMA_signal_2582), .Q (new_AGEMA_signal_7030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4513 ( .C (clk), .D (RoundKey[90]), .Q (new_AGEMA_signal_7034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4517 ( .C (clk), .D (new_AGEMA_signal_2690), .Q (new_AGEMA_signal_7038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4521 ( .C (clk), .D (KSSubBytesInput[25]), .Q (new_AGEMA_signal_7042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4525 ( .C (clk), .D (new_AGEMA_signal_2474), .Q (new_AGEMA_signal_7046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4529 ( .C (clk), .D (RoundKey[57]), .Q (new_AGEMA_signal_7050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4533 ( .C (clk), .D (new_AGEMA_signal_2579), .Q (new_AGEMA_signal_7054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4537 ( .C (clk), .D (RoundKey[89]), .Q (new_AGEMA_signal_7058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4541 ( .C (clk), .D (new_AGEMA_signal_2684), .Q (new_AGEMA_signal_7062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4545 ( .C (clk), .D (KSSubBytesInput[24]), .Q (new_AGEMA_signal_7066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4549 ( .C (clk), .D (new_AGEMA_signal_2471), .Q (new_AGEMA_signal_7070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4553 ( .C (clk), .D (RoundKey[56]), .Q (new_AGEMA_signal_7074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4557 ( .C (clk), .D (new_AGEMA_signal_2576), .Q (new_AGEMA_signal_7078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4561 ( .C (clk), .D (RoundKey[88]), .Q (new_AGEMA_signal_7082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4565 ( .C (clk), .D (new_AGEMA_signal_2681), .Q (new_AGEMA_signal_7086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4569 ( .C (clk), .D (KSSubBytesInput[7]), .Q (new_AGEMA_signal_7090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4573 ( .C (clk), .D (new_AGEMA_signal_2468), .Q (new_AGEMA_signal_7094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4577 ( .C (clk), .D (RoundKey[55]), .Q (new_AGEMA_signal_7098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4581 ( .C (clk), .D (new_AGEMA_signal_2573), .Q (new_AGEMA_signal_7102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4585 ( .C (clk), .D (RoundKey[87]), .Q (new_AGEMA_signal_7106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4589 ( .C (clk), .D (new_AGEMA_signal_2678), .Q (new_AGEMA_signal_7110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4593 ( .C (clk), .D (KSSubBytesInput[6]), .Q (new_AGEMA_signal_7114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4597 ( .C (clk), .D (new_AGEMA_signal_2465), .Q (new_AGEMA_signal_7118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4601 ( .C (clk), .D (RoundKey[54]), .Q (new_AGEMA_signal_7122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4605 ( .C (clk), .D (new_AGEMA_signal_2570), .Q (new_AGEMA_signal_7126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4609 ( .C (clk), .D (RoundKey[86]), .Q (new_AGEMA_signal_7130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4613 ( .C (clk), .D (new_AGEMA_signal_2675), .Q (new_AGEMA_signal_7134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4617 ( .C (clk), .D (KSSubBytesInput[5]), .Q (new_AGEMA_signal_7138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4621 ( .C (clk), .D (new_AGEMA_signal_2462), .Q (new_AGEMA_signal_7142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4625 ( .C (clk), .D (RoundKey[53]), .Q (new_AGEMA_signal_7146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4629 ( .C (clk), .D (new_AGEMA_signal_2567), .Q (new_AGEMA_signal_7150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4633 ( .C (clk), .D (RoundKey[85]), .Q (new_AGEMA_signal_7154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4637 ( .C (clk), .D (new_AGEMA_signal_2672), .Q (new_AGEMA_signal_7158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4641 ( .C (clk), .D (KSSubBytesInput[4]), .Q (new_AGEMA_signal_7162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4645 ( .C (clk), .D (new_AGEMA_signal_2459), .Q (new_AGEMA_signal_7166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4649 ( .C (clk), .D (RoundKey[52]), .Q (new_AGEMA_signal_7170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4653 ( .C (clk), .D (new_AGEMA_signal_2564), .Q (new_AGEMA_signal_7174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4657 ( .C (clk), .D (RoundKey[84]), .Q (new_AGEMA_signal_7178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4661 ( .C (clk), .D (new_AGEMA_signal_2669), .Q (new_AGEMA_signal_7182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4665 ( .C (clk), .D (KSSubBytesInput[17]), .Q (new_AGEMA_signal_7186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4669 ( .C (clk), .D (new_AGEMA_signal_2456), .Q (new_AGEMA_signal_7190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4673 ( .C (clk), .D (RoundKey[33]), .Q (new_AGEMA_signal_7194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4677 ( .C (clk), .D (new_AGEMA_signal_2501), .Q (new_AGEMA_signal_7198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4681 ( .C (clk), .D (RoundKey[65]), .Q (new_AGEMA_signal_7202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4685 ( .C (clk), .D (new_AGEMA_signal_2606), .Q (new_AGEMA_signal_7206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4689 ( .C (clk), .D (RoundKey[97]), .Q (new_AGEMA_signal_7210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4693 ( .C (clk), .D (new_AGEMA_signal_2711), .Q (new_AGEMA_signal_7214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4697 ( .C (clk), .D (KSSubBytesInput[3]), .Q (new_AGEMA_signal_7218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4701 ( .C (clk), .D (new_AGEMA_signal_2453), .Q (new_AGEMA_signal_7222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4705 ( .C (clk), .D (RoundKey[51]), .Q (new_AGEMA_signal_7226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4709 ( .C (clk), .D (new_AGEMA_signal_2561), .Q (new_AGEMA_signal_7230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4713 ( .C (clk), .D (RoundKey[83]), .Q (new_AGEMA_signal_7234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4717 ( .C (clk), .D (new_AGEMA_signal_2666), .Q (new_AGEMA_signal_7238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4721 ( .C (clk), .D (KSSubBytesInput[2]), .Q (new_AGEMA_signal_7242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4725 ( .C (clk), .D (new_AGEMA_signal_2450), .Q (new_AGEMA_signal_7246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4729 ( .C (clk), .D (RoundKey[50]), .Q (new_AGEMA_signal_7250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4733 ( .C (clk), .D (new_AGEMA_signal_2558), .Q (new_AGEMA_signal_7254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4737 ( .C (clk), .D (RoundKey[82]), .Q (new_AGEMA_signal_7258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4741 ( .C (clk), .D (new_AGEMA_signal_2663), .Q (new_AGEMA_signal_7262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4745 ( .C (clk), .D (KSSubBytesInput[1]), .Q (new_AGEMA_signal_7266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4749 ( .C (clk), .D (new_AGEMA_signal_2447), .Q (new_AGEMA_signal_7270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4753 ( .C (clk), .D (RoundKey[49]), .Q (new_AGEMA_signal_7274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4757 ( .C (clk), .D (new_AGEMA_signal_2552), .Q (new_AGEMA_signal_7278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4761 ( .C (clk), .D (RoundKey[81]), .Q (new_AGEMA_signal_7282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4765 ( .C (clk), .D (new_AGEMA_signal_2660), .Q (new_AGEMA_signal_7286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4769 ( .C (clk), .D (KSSubBytesInput[0]), .Q (new_AGEMA_signal_7290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4773 ( .C (clk), .D (new_AGEMA_signal_2444), .Q (new_AGEMA_signal_7294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4777 ( .C (clk), .D (RoundKey[48]), .Q (new_AGEMA_signal_7298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4781 ( .C (clk), .D (new_AGEMA_signal_2549), .Q (new_AGEMA_signal_7302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4785 ( .C (clk), .D (RoundKey[80]), .Q (new_AGEMA_signal_7306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4789 ( .C (clk), .D (new_AGEMA_signal_2657), .Q (new_AGEMA_signal_7310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4793 ( .C (clk), .D (KSSubBytesInput[15]), .Q (new_AGEMA_signal_7314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4797 ( .C (clk), .D (new_AGEMA_signal_2441), .Q (new_AGEMA_signal_7318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4801 ( .C (clk), .D (RoundKey[47]), .Q (new_AGEMA_signal_7322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4805 ( .C (clk), .D (new_AGEMA_signal_2546), .Q (new_AGEMA_signal_7326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4809 ( .C (clk), .D (RoundKey[79]), .Q (new_AGEMA_signal_7330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4813 ( .C (clk), .D (new_AGEMA_signal_2651), .Q (new_AGEMA_signal_7334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4817 ( .C (clk), .D (KSSubBytesInput[14]), .Q (new_AGEMA_signal_7338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4821 ( .C (clk), .D (new_AGEMA_signal_2438), .Q (new_AGEMA_signal_7342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4825 ( .C (clk), .D (RoundKey[46]), .Q (new_AGEMA_signal_7346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4829 ( .C (clk), .D (new_AGEMA_signal_2543), .Q (new_AGEMA_signal_7350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4833 ( .C (clk), .D (RoundKey[78]), .Q (new_AGEMA_signal_7354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4837 ( .C (clk), .D (new_AGEMA_signal_2648), .Q (new_AGEMA_signal_7358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4841 ( .C (clk), .D (KSSubBytesInput[13]), .Q (new_AGEMA_signal_7362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4845 ( .C (clk), .D (new_AGEMA_signal_2435), .Q (new_AGEMA_signal_7366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4849 ( .C (clk), .D (RoundKey[45]), .Q (new_AGEMA_signal_7370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4853 ( .C (clk), .D (new_AGEMA_signal_2540), .Q (new_AGEMA_signal_7374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4857 ( .C (clk), .D (RoundKey[77]), .Q (new_AGEMA_signal_7378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4861 ( .C (clk), .D (new_AGEMA_signal_2645), .Q (new_AGEMA_signal_7382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4865 ( .C (clk), .D (KSSubBytesInput[12]), .Q (new_AGEMA_signal_7386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4869 ( .C (clk), .D (new_AGEMA_signal_2432), .Q (new_AGEMA_signal_7390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4873 ( .C (clk), .D (RoundKey[44]), .Q (new_AGEMA_signal_7394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4877 ( .C (clk), .D (new_AGEMA_signal_2537), .Q (new_AGEMA_signal_7398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4881 ( .C (clk), .D (RoundKey[76]), .Q (new_AGEMA_signal_7402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4885 ( .C (clk), .D (new_AGEMA_signal_2642), .Q (new_AGEMA_signal_7406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4889 ( .C (clk), .D (RoundKey[127]), .Q (new_AGEMA_signal_7410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4893 ( .C (clk), .D (new_AGEMA_signal_2429), .Q (new_AGEMA_signal_7414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4897 ( .C (clk), .D (RoundKey[126]), .Q (new_AGEMA_signal_7418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4901 ( .C (clk), .D (new_AGEMA_signal_2426), .Q (new_AGEMA_signal_7422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4905 ( .C (clk), .D (RoundKey[125]), .Q (new_AGEMA_signal_7426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4909 ( .C (clk), .D (new_AGEMA_signal_2423), .Q (new_AGEMA_signal_7430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4913 ( .C (clk), .D (RoundKey[124]), .Q (new_AGEMA_signal_7434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4917 ( .C (clk), .D (new_AGEMA_signal_2420), .Q (new_AGEMA_signal_7438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4921 ( .C (clk), .D (RoundKey[123]), .Q (new_AGEMA_signal_7442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4925 ( .C (clk), .D (new_AGEMA_signal_2417), .Q (new_AGEMA_signal_7446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4929 ( .C (clk), .D (RoundKey[122]), .Q (new_AGEMA_signal_7450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4933 ( .C (clk), .D (new_AGEMA_signal_2414), .Q (new_AGEMA_signal_7454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4937 ( .C (clk), .D (RoundKey[121]), .Q (new_AGEMA_signal_7458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4941 ( .C (clk), .D (new_AGEMA_signal_2411), .Q (new_AGEMA_signal_7462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4945 ( .C (clk), .D (RoundKey[120]), .Q (new_AGEMA_signal_7466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4949 ( .C (clk), .D (new_AGEMA_signal_2408), .Q (new_AGEMA_signal_7470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4953 ( .C (clk), .D (KSSubBytesInput[11]), .Q (new_AGEMA_signal_7474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4957 ( .C (clk), .D (new_AGEMA_signal_2405), .Q (new_AGEMA_signal_7478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4961 ( .C (clk), .D (RoundKey[43]), .Q (new_AGEMA_signal_7482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4965 ( .C (clk), .D (new_AGEMA_signal_2534), .Q (new_AGEMA_signal_7486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4969 ( .C (clk), .D (RoundKey[75]), .Q (new_AGEMA_signal_7490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4973 ( .C (clk), .D (new_AGEMA_signal_2639), .Q (new_AGEMA_signal_7494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4977 ( .C (clk), .D (RoundKey[119]), .Q (new_AGEMA_signal_7498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4981 ( .C (clk), .D (new_AGEMA_signal_2402), .Q (new_AGEMA_signal_7502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4985 ( .C (clk), .D (RoundKey[118]), .Q (new_AGEMA_signal_7506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4989 ( .C (clk), .D (new_AGEMA_signal_2399), .Q (new_AGEMA_signal_7510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4993 ( .C (clk), .D (RoundKey[117]), .Q (new_AGEMA_signal_7514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4997 ( .C (clk), .D (new_AGEMA_signal_2396), .Q (new_AGEMA_signal_7518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5001 ( .C (clk), .D (RoundKey[116]), .Q (new_AGEMA_signal_7522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5005 ( .C (clk), .D (new_AGEMA_signal_2393), .Q (new_AGEMA_signal_7526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5009 ( .C (clk), .D (RoundKey[115]), .Q (new_AGEMA_signal_7530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5013 ( .C (clk), .D (new_AGEMA_signal_2390), .Q (new_AGEMA_signal_7534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5017 ( .C (clk), .D (RoundKey[114]), .Q (new_AGEMA_signal_7538) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5021 ( .C (clk), .D (new_AGEMA_signal_2387), .Q (new_AGEMA_signal_7542) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5025 ( .C (clk), .D (RoundKey[113]), .Q (new_AGEMA_signal_7546) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5029 ( .C (clk), .D (new_AGEMA_signal_2384), .Q (new_AGEMA_signal_7550) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5033 ( .C (clk), .D (RoundKey[112]), .Q (new_AGEMA_signal_7554) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5037 ( .C (clk), .D (new_AGEMA_signal_2381), .Q (new_AGEMA_signal_7558) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5041 ( .C (clk), .D (RoundKey[111]), .Q (new_AGEMA_signal_7562) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5045 ( .C (clk), .D (new_AGEMA_signal_2378), .Q (new_AGEMA_signal_7566) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5049 ( .C (clk), .D (RoundKey[110]), .Q (new_AGEMA_signal_7570) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5053 ( .C (clk), .D (new_AGEMA_signal_2375), .Q (new_AGEMA_signal_7574) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5057 ( .C (clk), .D (KSSubBytesInput[10]), .Q (new_AGEMA_signal_7578) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5061 ( .C (clk), .D (new_AGEMA_signal_2372), .Q (new_AGEMA_signal_7582) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5065 ( .C (clk), .D (RoundKey[42]), .Q (new_AGEMA_signal_7586) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5069 ( .C (clk), .D (new_AGEMA_signal_2531), .Q (new_AGEMA_signal_7590) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5073 ( .C (clk), .D (RoundKey[74]), .Q (new_AGEMA_signal_7594) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5077 ( .C (clk), .D (new_AGEMA_signal_2636), .Q (new_AGEMA_signal_7598) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5081 ( .C (clk), .D (RoundKey[109]), .Q (new_AGEMA_signal_7602) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5085 ( .C (clk), .D (new_AGEMA_signal_2369), .Q (new_AGEMA_signal_7606) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5089 ( .C (clk), .D (RoundKey[108]), .Q (new_AGEMA_signal_7610) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5093 ( .C (clk), .D (new_AGEMA_signal_2366), .Q (new_AGEMA_signal_7614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5097 ( .C (clk), .D (RoundKey[107]), .Q (new_AGEMA_signal_7618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5101 ( .C (clk), .D (new_AGEMA_signal_2363), .Q (new_AGEMA_signal_7622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5105 ( .C (clk), .D (RoundKey[106]), .Q (new_AGEMA_signal_7626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5109 ( .C (clk), .D (new_AGEMA_signal_2360), .Q (new_AGEMA_signal_7630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5113 ( .C (clk), .D (RoundKey[105]), .Q (new_AGEMA_signal_7634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5117 ( .C (clk), .D (new_AGEMA_signal_2357), .Q (new_AGEMA_signal_7638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5121 ( .C (clk), .D (RoundKey[104]), .Q (new_AGEMA_signal_7642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5125 ( .C (clk), .D (new_AGEMA_signal_2354), .Q (new_AGEMA_signal_7646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5129 ( .C (clk), .D (RoundKey[103]), .Q (new_AGEMA_signal_7650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5133 ( .C (clk), .D (new_AGEMA_signal_2351), .Q (new_AGEMA_signal_7654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5137 ( .C (clk), .D (RoundKey[102]), .Q (new_AGEMA_signal_7658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5141 ( .C (clk), .D (new_AGEMA_signal_2348), .Q (new_AGEMA_signal_7662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5145 ( .C (clk), .D (RoundKey[101]), .Q (new_AGEMA_signal_7666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5149 ( .C (clk), .D (new_AGEMA_signal_2345), .Q (new_AGEMA_signal_7670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5153 ( .C (clk), .D (RoundKey[100]), .Q (new_AGEMA_signal_7674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5157 ( .C (clk), .D (new_AGEMA_signal_2342), .Q (new_AGEMA_signal_7678) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5161 ( .C (clk), .D (KSSubBytesInput[16]), .Q (new_AGEMA_signal_7682) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5165 ( .C (clk), .D (new_AGEMA_signal_2339), .Q (new_AGEMA_signal_7686) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5169 ( .C (clk), .D (RoundKey[32]), .Q (new_AGEMA_signal_7690) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5173 ( .C (clk), .D (new_AGEMA_signal_2498), .Q (new_AGEMA_signal_7694) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5177 ( .C (clk), .D (RoundKey[64]), .Q (new_AGEMA_signal_7698) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5181 ( .C (clk), .D (new_AGEMA_signal_2603), .Q (new_AGEMA_signal_7702) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5185 ( .C (clk), .D (RoundKey[96]), .Q (new_AGEMA_signal_7706) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5189 ( .C (clk), .D (new_AGEMA_signal_2708), .Q (new_AGEMA_signal_7710) ) ;
    buf_clk new_AGEMA_reg_buffer_5193 ( .C (clk), .D (Rcon[7]), .Q (new_AGEMA_signal_7714) ) ;
    buf_clk new_AGEMA_reg_buffer_5197 ( .C (clk), .D (Rcon[6]), .Q (new_AGEMA_signal_7718) ) ;
    buf_clk new_AGEMA_reg_buffer_5201 ( .C (clk), .D (Rcon[5]), .Q (new_AGEMA_signal_7722) ) ;
    buf_clk new_AGEMA_reg_buffer_5205 ( .C (clk), .D (Rcon[4]), .Q (new_AGEMA_signal_7726) ) ;
    buf_clk new_AGEMA_reg_buffer_5209 ( .C (clk), .D (Rcon[3]), .Q (new_AGEMA_signal_7730) ) ;
    buf_clk new_AGEMA_reg_buffer_5213 ( .C (clk), .D (Rcon[2]), .Q (new_AGEMA_signal_7734) ) ;
    buf_clk new_AGEMA_reg_buffer_5217 ( .C (clk), .D (Rcon[1]), .Q (new_AGEMA_signal_7738) ) ;
    buf_clk new_AGEMA_reg_buffer_5221 ( .C (clk), .D (Rcon[0]), .Q (new_AGEMA_signal_7742) ) ;
    buf_clk new_AGEMA_reg_buffer_5225 ( .C (clk), .D (MuxKeyExpansion_n15), .Q (new_AGEMA_signal_7746) ) ;
    buf_clk new_AGEMA_reg_buffer_5229 ( .C (clk), .D (MuxKeyExpansion_n16), .Q (new_AGEMA_signal_7750) ) ;
    buf_clk new_AGEMA_reg_buffer_5233 ( .C (clk), .D (MuxKeyExpansion_n17), .Q (new_AGEMA_signal_7754) ) ;
    buf_clk new_AGEMA_reg_buffer_5237 ( .C (clk), .D (MuxKeyExpansion_n18), .Q (new_AGEMA_signal_7758) ) ;
    buf_clk new_AGEMA_reg_buffer_5241 ( .C (clk), .D (MuxKeyExpansion_n19), .Q (new_AGEMA_signal_7762) ) ;
    buf_clk new_AGEMA_reg_buffer_5245 ( .C (clk), .D (MuxKeyExpansion_n20), .Q (new_AGEMA_signal_7766) ) ;
    buf_clk new_AGEMA_reg_buffer_5249 ( .C (clk), .D (MuxKeyExpansion_n14), .Q (new_AGEMA_signal_7770) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5253 ( .C (clk), .D (RoundReg_Inst_ff_SDE_32_next_state), .Q (new_AGEMA_signal_7774) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5257 ( .C (clk), .D (new_AGEMA_signal_2851), .Q (new_AGEMA_signal_7778) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5261 ( .C (clk), .D (RoundReg_Inst_ff_SDE_33_next_state), .Q (new_AGEMA_signal_7782) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5265 ( .C (clk), .D (new_AGEMA_signal_2853), .Q (new_AGEMA_signal_7786) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5269 ( .C (clk), .D (RoundReg_Inst_ff_SDE_34_next_state), .Q (new_AGEMA_signal_7790) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5273 ( .C (clk), .D (new_AGEMA_signal_2855), .Q (new_AGEMA_signal_7794) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5277 ( .C (clk), .D (RoundReg_Inst_ff_SDE_35_next_state), .Q (new_AGEMA_signal_7798) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5281 ( .C (clk), .D (new_AGEMA_signal_2857), .Q (new_AGEMA_signal_7802) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5285 ( .C (clk), .D (RoundReg_Inst_ff_SDE_36_next_state), .Q (new_AGEMA_signal_7806) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5289 ( .C (clk), .D (new_AGEMA_signal_2859), .Q (new_AGEMA_signal_7810) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5293 ( .C (clk), .D (RoundReg_Inst_ff_SDE_37_next_state), .Q (new_AGEMA_signal_7814) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5297 ( .C (clk), .D (new_AGEMA_signal_2861), .Q (new_AGEMA_signal_7818) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5301 ( .C (clk), .D (RoundReg_Inst_ff_SDE_38_next_state), .Q (new_AGEMA_signal_7822) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5305 ( .C (clk), .D (new_AGEMA_signal_2863), .Q (new_AGEMA_signal_7826) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5309 ( .C (clk), .D (RoundReg_Inst_ff_SDE_39_next_state), .Q (new_AGEMA_signal_7830) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5313 ( .C (clk), .D (new_AGEMA_signal_2865), .Q (new_AGEMA_signal_7834) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5317 ( .C (clk), .D (RoundReg_Inst_ff_SDE_40_next_state), .Q (new_AGEMA_signal_7838) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5321 ( .C (clk), .D (new_AGEMA_signal_2867), .Q (new_AGEMA_signal_7842) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5325 ( .C (clk), .D (RoundReg_Inst_ff_SDE_41_next_state), .Q (new_AGEMA_signal_7846) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5329 ( .C (clk), .D (new_AGEMA_signal_2869), .Q (new_AGEMA_signal_7850) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5333 ( .C (clk), .D (RoundReg_Inst_ff_SDE_42_next_state), .Q (new_AGEMA_signal_7854) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5337 ( .C (clk), .D (new_AGEMA_signal_2871), .Q (new_AGEMA_signal_7858) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5341 ( .C (clk), .D (RoundReg_Inst_ff_SDE_43_next_state), .Q (new_AGEMA_signal_7862) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5345 ( .C (clk), .D (new_AGEMA_signal_2873), .Q (new_AGEMA_signal_7866) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5349 ( .C (clk), .D (RoundReg_Inst_ff_SDE_44_next_state), .Q (new_AGEMA_signal_7870) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5353 ( .C (clk), .D (new_AGEMA_signal_2875), .Q (new_AGEMA_signal_7874) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5357 ( .C (clk), .D (RoundReg_Inst_ff_SDE_45_next_state), .Q (new_AGEMA_signal_7878) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5361 ( .C (clk), .D (new_AGEMA_signal_2877), .Q (new_AGEMA_signal_7882) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5365 ( .C (clk), .D (RoundReg_Inst_ff_SDE_46_next_state), .Q (new_AGEMA_signal_7886) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5369 ( .C (clk), .D (new_AGEMA_signal_2879), .Q (new_AGEMA_signal_7890) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5373 ( .C (clk), .D (RoundReg_Inst_ff_SDE_47_next_state), .Q (new_AGEMA_signal_7894) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5377 ( .C (clk), .D (new_AGEMA_signal_2881), .Q (new_AGEMA_signal_7898) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5381 ( .C (clk), .D (RoundReg_Inst_ff_SDE_48_next_state), .Q (new_AGEMA_signal_7902) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5385 ( .C (clk), .D (new_AGEMA_signal_2883), .Q (new_AGEMA_signal_7906) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5389 ( .C (clk), .D (RoundReg_Inst_ff_SDE_49_next_state), .Q (new_AGEMA_signal_7910) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5393 ( .C (clk), .D (new_AGEMA_signal_2885), .Q (new_AGEMA_signal_7914) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5397 ( .C (clk), .D (RoundReg_Inst_ff_SDE_50_next_state), .Q (new_AGEMA_signal_7918) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5401 ( .C (clk), .D (new_AGEMA_signal_2887), .Q (new_AGEMA_signal_7922) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5405 ( .C (clk), .D (RoundReg_Inst_ff_SDE_51_next_state), .Q (new_AGEMA_signal_7926) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5409 ( .C (clk), .D (new_AGEMA_signal_2889), .Q (new_AGEMA_signal_7930) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5413 ( .C (clk), .D (RoundReg_Inst_ff_SDE_52_next_state), .Q (new_AGEMA_signal_7934) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5417 ( .C (clk), .D (new_AGEMA_signal_2891), .Q (new_AGEMA_signal_7938) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5421 ( .C (clk), .D (RoundReg_Inst_ff_SDE_53_next_state), .Q (new_AGEMA_signal_7942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5425 ( .C (clk), .D (new_AGEMA_signal_2893), .Q (new_AGEMA_signal_7946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5429 ( .C (clk), .D (RoundReg_Inst_ff_SDE_54_next_state), .Q (new_AGEMA_signal_7950) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5433 ( .C (clk), .D (new_AGEMA_signal_2895), .Q (new_AGEMA_signal_7954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5437 ( .C (clk), .D (RoundReg_Inst_ff_SDE_55_next_state), .Q (new_AGEMA_signal_7958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5441 ( .C (clk), .D (new_AGEMA_signal_2897), .Q (new_AGEMA_signal_7962) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5445 ( .C (clk), .D (RoundReg_Inst_ff_SDE_56_next_state), .Q (new_AGEMA_signal_7966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5449 ( .C (clk), .D (new_AGEMA_signal_2899), .Q (new_AGEMA_signal_7970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5453 ( .C (clk), .D (RoundReg_Inst_ff_SDE_57_next_state), .Q (new_AGEMA_signal_7974) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5457 ( .C (clk), .D (new_AGEMA_signal_2901), .Q (new_AGEMA_signal_7978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5461 ( .C (clk), .D (RoundReg_Inst_ff_SDE_58_next_state), .Q (new_AGEMA_signal_7982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5465 ( .C (clk), .D (new_AGEMA_signal_2903), .Q (new_AGEMA_signal_7986) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5469 ( .C (clk), .D (RoundReg_Inst_ff_SDE_59_next_state), .Q (new_AGEMA_signal_7990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5473 ( .C (clk), .D (new_AGEMA_signal_2905), .Q (new_AGEMA_signal_7994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5477 ( .C (clk), .D (RoundReg_Inst_ff_SDE_60_next_state), .Q (new_AGEMA_signal_7998) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5481 ( .C (clk), .D (new_AGEMA_signal_2907), .Q (new_AGEMA_signal_8002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5485 ( .C (clk), .D (RoundReg_Inst_ff_SDE_61_next_state), .Q (new_AGEMA_signal_8006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5489 ( .C (clk), .D (new_AGEMA_signal_2909), .Q (new_AGEMA_signal_8010) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5493 ( .C (clk), .D (RoundReg_Inst_ff_SDE_62_next_state), .Q (new_AGEMA_signal_8014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5497 ( .C (clk), .D (new_AGEMA_signal_2911), .Q (new_AGEMA_signal_8018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5501 ( .C (clk), .D (RoundReg_Inst_ff_SDE_63_next_state), .Q (new_AGEMA_signal_8022) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5505 ( .C (clk), .D (new_AGEMA_signal_2913), .Q (new_AGEMA_signal_8026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5509 ( .C (clk), .D (RoundReg_Inst_ff_SDE_64_next_state), .Q (new_AGEMA_signal_8030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5513 ( .C (clk), .D (new_AGEMA_signal_2915), .Q (new_AGEMA_signal_8034) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5517 ( .C (clk), .D (RoundReg_Inst_ff_SDE_65_next_state), .Q (new_AGEMA_signal_8038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5521 ( .C (clk), .D (new_AGEMA_signal_2917), .Q (new_AGEMA_signal_8042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5525 ( .C (clk), .D (RoundReg_Inst_ff_SDE_66_next_state), .Q (new_AGEMA_signal_8046) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5529 ( .C (clk), .D (new_AGEMA_signal_2919), .Q (new_AGEMA_signal_8050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5533 ( .C (clk), .D (RoundReg_Inst_ff_SDE_67_next_state), .Q (new_AGEMA_signal_8054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5537 ( .C (clk), .D (new_AGEMA_signal_2921), .Q (new_AGEMA_signal_8058) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5541 ( .C (clk), .D (RoundReg_Inst_ff_SDE_68_next_state), .Q (new_AGEMA_signal_8062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5545 ( .C (clk), .D (new_AGEMA_signal_2923), .Q (new_AGEMA_signal_8066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5549 ( .C (clk), .D (RoundReg_Inst_ff_SDE_69_next_state), .Q (new_AGEMA_signal_8070) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5553 ( .C (clk), .D (new_AGEMA_signal_2925), .Q (new_AGEMA_signal_8074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5557 ( .C (clk), .D (RoundReg_Inst_ff_SDE_70_next_state), .Q (new_AGEMA_signal_8078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5561 ( .C (clk), .D (new_AGEMA_signal_2927), .Q (new_AGEMA_signal_8082) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5565 ( .C (clk), .D (RoundReg_Inst_ff_SDE_71_next_state), .Q (new_AGEMA_signal_8086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5569 ( .C (clk), .D (new_AGEMA_signal_2929), .Q (new_AGEMA_signal_8090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5573 ( .C (clk), .D (RoundReg_Inst_ff_SDE_72_next_state), .Q (new_AGEMA_signal_8094) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5577 ( .C (clk), .D (new_AGEMA_signal_2931), .Q (new_AGEMA_signal_8098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5581 ( .C (clk), .D (RoundReg_Inst_ff_SDE_73_next_state), .Q (new_AGEMA_signal_8102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5585 ( .C (clk), .D (new_AGEMA_signal_2933), .Q (new_AGEMA_signal_8106) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5589 ( .C (clk), .D (RoundReg_Inst_ff_SDE_74_next_state), .Q (new_AGEMA_signal_8110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5593 ( .C (clk), .D (new_AGEMA_signal_2935), .Q (new_AGEMA_signal_8114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5597 ( .C (clk), .D (RoundReg_Inst_ff_SDE_75_next_state), .Q (new_AGEMA_signal_8118) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5601 ( .C (clk), .D (new_AGEMA_signal_2937), .Q (new_AGEMA_signal_8122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5605 ( .C (clk), .D (RoundReg_Inst_ff_SDE_76_next_state), .Q (new_AGEMA_signal_8126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5609 ( .C (clk), .D (new_AGEMA_signal_2939), .Q (new_AGEMA_signal_8130) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5613 ( .C (clk), .D (RoundReg_Inst_ff_SDE_77_next_state), .Q (new_AGEMA_signal_8134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5617 ( .C (clk), .D (new_AGEMA_signal_2941), .Q (new_AGEMA_signal_8138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5621 ( .C (clk), .D (RoundReg_Inst_ff_SDE_78_next_state), .Q (new_AGEMA_signal_8142) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5625 ( .C (clk), .D (new_AGEMA_signal_2943), .Q (new_AGEMA_signal_8146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5629 ( .C (clk), .D (RoundReg_Inst_ff_SDE_79_next_state), .Q (new_AGEMA_signal_8150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5633 ( .C (clk), .D (new_AGEMA_signal_2945), .Q (new_AGEMA_signal_8154) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5637 ( .C (clk), .D (RoundReg_Inst_ff_SDE_80_next_state), .Q (new_AGEMA_signal_8158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5641 ( .C (clk), .D (new_AGEMA_signal_2947), .Q (new_AGEMA_signal_8162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5645 ( .C (clk), .D (RoundReg_Inst_ff_SDE_81_next_state), .Q (new_AGEMA_signal_8166) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5649 ( .C (clk), .D (new_AGEMA_signal_2949), .Q (new_AGEMA_signal_8170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5653 ( .C (clk), .D (RoundReg_Inst_ff_SDE_82_next_state), .Q (new_AGEMA_signal_8174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5657 ( .C (clk), .D (new_AGEMA_signal_2951), .Q (new_AGEMA_signal_8178) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5661 ( .C (clk), .D (RoundReg_Inst_ff_SDE_83_next_state), .Q (new_AGEMA_signal_8182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5665 ( .C (clk), .D (new_AGEMA_signal_2953), .Q (new_AGEMA_signal_8186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5669 ( .C (clk), .D (RoundReg_Inst_ff_SDE_84_next_state), .Q (new_AGEMA_signal_8190) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5673 ( .C (clk), .D (new_AGEMA_signal_2955), .Q (new_AGEMA_signal_8194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5677 ( .C (clk), .D (RoundReg_Inst_ff_SDE_85_next_state), .Q (new_AGEMA_signal_8198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5681 ( .C (clk), .D (new_AGEMA_signal_2957), .Q (new_AGEMA_signal_8202) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5685 ( .C (clk), .D (RoundReg_Inst_ff_SDE_86_next_state), .Q (new_AGEMA_signal_8206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5689 ( .C (clk), .D (new_AGEMA_signal_2959), .Q (new_AGEMA_signal_8210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5693 ( .C (clk), .D (RoundReg_Inst_ff_SDE_87_next_state), .Q (new_AGEMA_signal_8214) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5697 ( .C (clk), .D (new_AGEMA_signal_2961), .Q (new_AGEMA_signal_8218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5701 ( .C (clk), .D (RoundReg_Inst_ff_SDE_88_next_state), .Q (new_AGEMA_signal_8222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5705 ( .C (clk), .D (new_AGEMA_signal_2963), .Q (new_AGEMA_signal_8226) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5709 ( .C (clk), .D (RoundReg_Inst_ff_SDE_89_next_state), .Q (new_AGEMA_signal_8230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5713 ( .C (clk), .D (new_AGEMA_signal_2965), .Q (new_AGEMA_signal_8234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5717 ( .C (clk), .D (RoundReg_Inst_ff_SDE_90_next_state), .Q (new_AGEMA_signal_8238) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5721 ( .C (clk), .D (new_AGEMA_signal_2967), .Q (new_AGEMA_signal_8242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5725 ( .C (clk), .D (RoundReg_Inst_ff_SDE_91_next_state), .Q (new_AGEMA_signal_8246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5729 ( .C (clk), .D (new_AGEMA_signal_2969), .Q (new_AGEMA_signal_8250) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5733 ( .C (clk), .D (RoundReg_Inst_ff_SDE_92_next_state), .Q (new_AGEMA_signal_8254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5737 ( .C (clk), .D (new_AGEMA_signal_2971), .Q (new_AGEMA_signal_8258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5741 ( .C (clk), .D (RoundReg_Inst_ff_SDE_93_next_state), .Q (new_AGEMA_signal_8262) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5745 ( .C (clk), .D (new_AGEMA_signal_2973), .Q (new_AGEMA_signal_8266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5749 ( .C (clk), .D (RoundReg_Inst_ff_SDE_94_next_state), .Q (new_AGEMA_signal_8270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5753 ( .C (clk), .D (new_AGEMA_signal_2975), .Q (new_AGEMA_signal_8274) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5757 ( .C (clk), .D (RoundReg_Inst_ff_SDE_95_next_state), .Q (new_AGEMA_signal_8278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5761 ( .C (clk), .D (new_AGEMA_signal_2977), .Q (new_AGEMA_signal_8282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5765 ( .C (clk), .D (RoundReg_Inst_ff_SDE_96_next_state), .Q (new_AGEMA_signal_8286) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5769 ( .C (clk), .D (new_AGEMA_signal_2979), .Q (new_AGEMA_signal_8290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5773 ( .C (clk), .D (RoundReg_Inst_ff_SDE_97_next_state), .Q (new_AGEMA_signal_8294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5777 ( .C (clk), .D (new_AGEMA_signal_2981), .Q (new_AGEMA_signal_8298) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5781 ( .C (clk), .D (RoundReg_Inst_ff_SDE_98_next_state), .Q (new_AGEMA_signal_8302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5785 ( .C (clk), .D (new_AGEMA_signal_2983), .Q (new_AGEMA_signal_8306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5789 ( .C (clk), .D (RoundReg_Inst_ff_SDE_99_next_state), .Q (new_AGEMA_signal_8310) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5793 ( .C (clk), .D (new_AGEMA_signal_2985), .Q (new_AGEMA_signal_8314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5797 ( .C (clk), .D (RoundReg_Inst_ff_SDE_100_next_state), .Q (new_AGEMA_signal_8318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5801 ( .C (clk), .D (new_AGEMA_signal_2987), .Q (new_AGEMA_signal_8322) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5805 ( .C (clk), .D (RoundReg_Inst_ff_SDE_101_next_state), .Q (new_AGEMA_signal_8326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5809 ( .C (clk), .D (new_AGEMA_signal_2989), .Q (new_AGEMA_signal_8330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5813 ( .C (clk), .D (RoundReg_Inst_ff_SDE_102_next_state), .Q (new_AGEMA_signal_8334) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5817 ( .C (clk), .D (new_AGEMA_signal_2991), .Q (new_AGEMA_signal_8338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5821 ( .C (clk), .D (RoundReg_Inst_ff_SDE_103_next_state), .Q (new_AGEMA_signal_8342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5825 ( .C (clk), .D (new_AGEMA_signal_2993), .Q (new_AGEMA_signal_8346) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5829 ( .C (clk), .D (RoundReg_Inst_ff_SDE_104_next_state), .Q (new_AGEMA_signal_8350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5833 ( .C (clk), .D (new_AGEMA_signal_2995), .Q (new_AGEMA_signal_8354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5837 ( .C (clk), .D (RoundReg_Inst_ff_SDE_105_next_state), .Q (new_AGEMA_signal_8358) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5841 ( .C (clk), .D (new_AGEMA_signal_2997), .Q (new_AGEMA_signal_8362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5845 ( .C (clk), .D (RoundReg_Inst_ff_SDE_106_next_state), .Q (new_AGEMA_signal_8366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5849 ( .C (clk), .D (new_AGEMA_signal_2999), .Q (new_AGEMA_signal_8370) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5853 ( .C (clk), .D (RoundReg_Inst_ff_SDE_107_next_state), .Q (new_AGEMA_signal_8374) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5857 ( .C (clk), .D (new_AGEMA_signal_3001), .Q (new_AGEMA_signal_8378) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5861 ( .C (clk), .D (RoundReg_Inst_ff_SDE_108_next_state), .Q (new_AGEMA_signal_8382) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5865 ( .C (clk), .D (new_AGEMA_signal_3003), .Q (new_AGEMA_signal_8386) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5869 ( .C (clk), .D (RoundReg_Inst_ff_SDE_109_next_state), .Q (new_AGEMA_signal_8390) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5873 ( .C (clk), .D (new_AGEMA_signal_3005), .Q (new_AGEMA_signal_8394) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5877 ( .C (clk), .D (RoundReg_Inst_ff_SDE_110_next_state), .Q (new_AGEMA_signal_8398) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5881 ( .C (clk), .D (new_AGEMA_signal_3007), .Q (new_AGEMA_signal_8402) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5885 ( .C (clk), .D (RoundReg_Inst_ff_SDE_111_next_state), .Q (new_AGEMA_signal_8406) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5889 ( .C (clk), .D (new_AGEMA_signal_3009), .Q (new_AGEMA_signal_8410) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5893 ( .C (clk), .D (RoundReg_Inst_ff_SDE_112_next_state), .Q (new_AGEMA_signal_8414) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5897 ( .C (clk), .D (new_AGEMA_signal_3011), .Q (new_AGEMA_signal_8418) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5901 ( .C (clk), .D (RoundReg_Inst_ff_SDE_113_next_state), .Q (new_AGEMA_signal_8422) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5905 ( .C (clk), .D (new_AGEMA_signal_3013), .Q (new_AGEMA_signal_8426) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5909 ( .C (clk), .D (RoundReg_Inst_ff_SDE_114_next_state), .Q (new_AGEMA_signal_8430) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5913 ( .C (clk), .D (new_AGEMA_signal_3015), .Q (new_AGEMA_signal_8434) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5917 ( .C (clk), .D (RoundReg_Inst_ff_SDE_115_next_state), .Q (new_AGEMA_signal_8438) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5921 ( .C (clk), .D (new_AGEMA_signal_3017), .Q (new_AGEMA_signal_8442) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5925 ( .C (clk), .D (RoundReg_Inst_ff_SDE_116_next_state), .Q (new_AGEMA_signal_8446) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5929 ( .C (clk), .D (new_AGEMA_signal_3019), .Q (new_AGEMA_signal_8450) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5933 ( .C (clk), .D (RoundReg_Inst_ff_SDE_117_next_state), .Q (new_AGEMA_signal_8454) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5937 ( .C (clk), .D (new_AGEMA_signal_3021), .Q (new_AGEMA_signal_8458) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5941 ( .C (clk), .D (RoundReg_Inst_ff_SDE_118_next_state), .Q (new_AGEMA_signal_8462) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5945 ( .C (clk), .D (new_AGEMA_signal_3023), .Q (new_AGEMA_signal_8466) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5949 ( .C (clk), .D (RoundReg_Inst_ff_SDE_119_next_state), .Q (new_AGEMA_signal_8470) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5953 ( .C (clk), .D (new_AGEMA_signal_3025), .Q (new_AGEMA_signal_8474) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5957 ( .C (clk), .D (RoundReg_Inst_ff_SDE_120_next_state), .Q (new_AGEMA_signal_8478) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5961 ( .C (clk), .D (new_AGEMA_signal_3027), .Q (new_AGEMA_signal_8482) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5965 ( .C (clk), .D (RoundReg_Inst_ff_SDE_121_next_state), .Q (new_AGEMA_signal_8486) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5969 ( .C (clk), .D (new_AGEMA_signal_3029), .Q (new_AGEMA_signal_8490) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5973 ( .C (clk), .D (RoundReg_Inst_ff_SDE_122_next_state), .Q (new_AGEMA_signal_8494) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5977 ( .C (clk), .D (new_AGEMA_signal_3031), .Q (new_AGEMA_signal_8498) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5981 ( .C (clk), .D (RoundReg_Inst_ff_SDE_123_next_state), .Q (new_AGEMA_signal_8502) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5985 ( .C (clk), .D (new_AGEMA_signal_3033), .Q (new_AGEMA_signal_8506) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5989 ( .C (clk), .D (RoundReg_Inst_ff_SDE_124_next_state), .Q (new_AGEMA_signal_8510) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5993 ( .C (clk), .D (new_AGEMA_signal_3035), .Q (new_AGEMA_signal_8514) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5997 ( .C (clk), .D (RoundReg_Inst_ff_SDE_125_next_state), .Q (new_AGEMA_signal_8518) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6001 ( .C (clk), .D (new_AGEMA_signal_3037), .Q (new_AGEMA_signal_8522) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6005 ( .C (clk), .D (RoundReg_Inst_ff_SDE_126_next_state), .Q (new_AGEMA_signal_8526) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6009 ( .C (clk), .D (new_AGEMA_signal_3039), .Q (new_AGEMA_signal_8530) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6013 ( .C (clk), .D (RoundReg_Inst_ff_SDE_127_next_state), .Q (new_AGEMA_signal_8534) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6017 ( .C (clk), .D (new_AGEMA_signal_3041), .Q (new_AGEMA_signal_8538) ) ;
    buf_clk new_AGEMA_reg_buffer_6021 ( .C (clk), .D (RoundCounterIns_n45), .Q (new_AGEMA_signal_8542) ) ;
    buf_clk new_AGEMA_reg_buffer_6025 ( .C (clk), .D (RoundCounterIns_n44), .Q (new_AGEMA_signal_8546) ) ;
    buf_clk new_AGEMA_reg_buffer_6029 ( .C (clk), .D (RoundCounterIns_n1), .Q (new_AGEMA_signal_8550) ) ;
    buf_clk new_AGEMA_reg_buffer_6033 ( .C (clk), .D (RoundCounterIns_n42), .Q (new_AGEMA_signal_8554) ) ;
    buf_clk new_AGEMA_reg_buffer_6037 ( .C (clk), .D (InRoundCounterIns_n41), .Q (new_AGEMA_signal_8558) ) ;
    buf_clk new_AGEMA_reg_buffer_6041 ( .C (clk), .D (InRoundCounterIns_n40), .Q (new_AGEMA_signal_8562) ) ;
    buf_clk new_AGEMA_reg_buffer_6045 ( .C (clk), .D (InRoundCounterIns_n39), .Q (new_AGEMA_signal_8566) ) ;

    /* cells in depth 2 */
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_4615, new_AGEMA_signal_4614}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3255, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_4617, new_AGEMA_signal_4616}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3256, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_3223, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_3238, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[75], Fresh[74]}), .c ({new_AGEMA_signal_3257, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_4619, new_AGEMA_signal_4618}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3258, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_3224, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_3225, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[77], Fresh[76]}), .c ({new_AGEMA_signal_3241, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_4621, new_AGEMA_signal_4620}), .b ({new_AGEMA_signal_3239, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_3278, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_4623, new_AGEMA_signal_4622}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3260, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_4625, new_AGEMA_signal_4624}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3261, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_3227, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_3242, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_3262, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4626}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3263, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_3228, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_3229, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[83], Fresh[82]}), .c ({new_AGEMA_signal_3245, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_4629, new_AGEMA_signal_4628}), .b ({new_AGEMA_signal_3243, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_3283, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_4631, new_AGEMA_signal_4630}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3265, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_4633, new_AGEMA_signal_4632}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3266, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_3231, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_3246, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[87], Fresh[86]}), .c ({new_AGEMA_signal_3267, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_4635, new_AGEMA_signal_4634}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3268, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_3232, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_3233, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[89], Fresh[88]}), .c ({new_AGEMA_signal_3249, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_4637, new_AGEMA_signal_4636}), .b ({new_AGEMA_signal_3247, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_3288, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_4639, new_AGEMA_signal_4638}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3270, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_4641, new_AGEMA_signal_4640}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3271, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_3235, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_3250, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[93], Fresh[92]}), .c ({new_AGEMA_signal_3272, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_4643, new_AGEMA_signal_4642}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3273, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_3236, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_3237, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[95], Fresh[94]}), .c ({new_AGEMA_signal_3253, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_4645, new_AGEMA_signal_4644}), .b ({new_AGEMA_signal_3251, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_3293, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2093 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M21), .Q (new_AGEMA_signal_4614) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2094 ( .C (clk), .D (new_AGEMA_signal_3224), .Q (new_AGEMA_signal_4615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2095 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M23), .Q (new_AGEMA_signal_4616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2096 ( .C (clk), .D (new_AGEMA_signal_3238), .Q (new_AGEMA_signal_4617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2097 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M27), .Q (new_AGEMA_signal_4618) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2098 ( .C (clk), .D (new_AGEMA_signal_3240), .Q (new_AGEMA_signal_4619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2099 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M24), .Q (new_AGEMA_signal_4620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2100 ( .C (clk), .D (new_AGEMA_signal_3254), .Q (new_AGEMA_signal_4621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2101 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M21), .Q (new_AGEMA_signal_4622) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2102 ( .C (clk), .D (new_AGEMA_signal_3228), .Q (new_AGEMA_signal_4623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2103 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M23), .Q (new_AGEMA_signal_4624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2104 ( .C (clk), .D (new_AGEMA_signal_3242), .Q (new_AGEMA_signal_4625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2105 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M27), .Q (new_AGEMA_signal_4626) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2106 ( .C (clk), .D (new_AGEMA_signal_3244), .Q (new_AGEMA_signal_4627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2107 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M24), .Q (new_AGEMA_signal_4628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2108 ( .C (clk), .D (new_AGEMA_signal_3259), .Q (new_AGEMA_signal_4629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2109 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M21), .Q (new_AGEMA_signal_4630) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2110 ( .C (clk), .D (new_AGEMA_signal_3232), .Q (new_AGEMA_signal_4631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2111 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M23), .Q (new_AGEMA_signal_4632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2112 ( .C (clk), .D (new_AGEMA_signal_3246), .Q (new_AGEMA_signal_4633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2113 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M27), .Q (new_AGEMA_signal_4634) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2114 ( .C (clk), .D (new_AGEMA_signal_3248), .Q (new_AGEMA_signal_4635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2115 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M24), .Q (new_AGEMA_signal_4636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2116 ( .C (clk), .D (new_AGEMA_signal_3264), .Q (new_AGEMA_signal_4637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2117 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M21), .Q (new_AGEMA_signal_4638) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2118 ( .C (clk), .D (new_AGEMA_signal_3236), .Q (new_AGEMA_signal_4639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2119 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M23), .Q (new_AGEMA_signal_4640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2120 ( .C (clk), .D (new_AGEMA_signal_3250), .Q (new_AGEMA_signal_4641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2121 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M27), .Q (new_AGEMA_signal_4642) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2122 ( .C (clk), .D (new_AGEMA_signal_3252), .Q (new_AGEMA_signal_4643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2123 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M24), .Q (new_AGEMA_signal_4644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2124 ( .C (clk), .D (new_AGEMA_signal_3269), .Q (new_AGEMA_signal_4645) ) ;
    buf_clk new_AGEMA_reg_buffer_2158 ( .C (clk), .D (new_AGEMA_signal_4678), .Q (new_AGEMA_signal_4679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2162 ( .C (clk), .D (new_AGEMA_signal_4682), .Q (new_AGEMA_signal_4683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2166 ( .C (clk), .D (new_AGEMA_signal_4686), .Q (new_AGEMA_signal_4687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2170 ( .C (clk), .D (new_AGEMA_signal_4690), .Q (new_AGEMA_signal_4691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2174 ( .C (clk), .D (new_AGEMA_signal_4694), .Q (new_AGEMA_signal_4695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2178 ( .C (clk), .D (new_AGEMA_signal_4698), .Q (new_AGEMA_signal_4699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2182 ( .C (clk), .D (new_AGEMA_signal_4702), .Q (new_AGEMA_signal_4703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2186 ( .C (clk), .D (new_AGEMA_signal_4706), .Q (new_AGEMA_signal_4707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2190 ( .C (clk), .D (new_AGEMA_signal_4710), .Q (new_AGEMA_signal_4711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2194 ( .C (clk), .D (new_AGEMA_signal_4714), .Q (new_AGEMA_signal_4715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2198 ( .C (clk), .D (new_AGEMA_signal_4718), .Q (new_AGEMA_signal_4719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2202 ( .C (clk), .D (new_AGEMA_signal_4722), .Q (new_AGEMA_signal_4723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2206 ( .C (clk), .D (new_AGEMA_signal_4726), .Q (new_AGEMA_signal_4727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2210 ( .C (clk), .D (new_AGEMA_signal_4730), .Q (new_AGEMA_signal_4731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2214 ( .C (clk), .D (new_AGEMA_signal_4734), .Q (new_AGEMA_signal_4735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2218 ( .C (clk), .D (new_AGEMA_signal_4738), .Q (new_AGEMA_signal_4739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2222 ( .C (clk), .D (new_AGEMA_signal_4742), .Q (new_AGEMA_signal_4743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2226 ( .C (clk), .D (new_AGEMA_signal_4746), .Q (new_AGEMA_signal_4747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2230 ( .C (clk), .D (new_AGEMA_signal_4750), .Q (new_AGEMA_signal_4751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2234 ( .C (clk), .D (new_AGEMA_signal_4754), .Q (new_AGEMA_signal_4755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2238 ( .C (clk), .D (new_AGEMA_signal_4758), .Q (new_AGEMA_signal_4759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2242 ( .C (clk), .D (new_AGEMA_signal_4762), .Q (new_AGEMA_signal_4763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2246 ( .C (clk), .D (new_AGEMA_signal_4766), .Q (new_AGEMA_signal_4767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2250 ( .C (clk), .D (new_AGEMA_signal_4770), .Q (new_AGEMA_signal_4771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2254 ( .C (clk), .D (new_AGEMA_signal_4774), .Q (new_AGEMA_signal_4775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2258 ( .C (clk), .D (new_AGEMA_signal_4778), .Q (new_AGEMA_signal_4779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2262 ( .C (clk), .D (new_AGEMA_signal_4782), .Q (new_AGEMA_signal_4783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2266 ( .C (clk), .D (new_AGEMA_signal_4786), .Q (new_AGEMA_signal_4787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2270 ( .C (clk), .D (new_AGEMA_signal_4790), .Q (new_AGEMA_signal_4791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2274 ( .C (clk), .D (new_AGEMA_signal_4794), .Q (new_AGEMA_signal_4795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2278 ( .C (clk), .D (new_AGEMA_signal_4798), .Q (new_AGEMA_signal_4799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2282 ( .C (clk), .D (new_AGEMA_signal_4802), .Q (new_AGEMA_signal_4803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2286 ( .C (clk), .D (new_AGEMA_signal_4806), .Q (new_AGEMA_signal_4807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2290 ( .C (clk), .D (new_AGEMA_signal_4810), .Q (new_AGEMA_signal_4811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2294 ( .C (clk), .D (new_AGEMA_signal_4814), .Q (new_AGEMA_signal_4815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2298 ( .C (clk), .D (new_AGEMA_signal_4818), .Q (new_AGEMA_signal_4819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2302 ( .C (clk), .D (new_AGEMA_signal_4822), .Q (new_AGEMA_signal_4823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2306 ( .C (clk), .D (new_AGEMA_signal_4826), .Q (new_AGEMA_signal_4827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2310 ( .C (clk), .D (new_AGEMA_signal_4830), .Q (new_AGEMA_signal_4831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2314 ( .C (clk), .D (new_AGEMA_signal_4834), .Q (new_AGEMA_signal_4835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2318 ( .C (clk), .D (new_AGEMA_signal_4838), .Q (new_AGEMA_signal_4839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2322 ( .C (clk), .D (new_AGEMA_signal_4842), .Q (new_AGEMA_signal_4843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2326 ( .C (clk), .D (new_AGEMA_signal_4846), .Q (new_AGEMA_signal_4847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2330 ( .C (clk), .D (new_AGEMA_signal_4850), .Q (new_AGEMA_signal_4851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2334 ( .C (clk), .D (new_AGEMA_signal_4854), .Q (new_AGEMA_signal_4855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2338 ( .C (clk), .D (new_AGEMA_signal_4858), .Q (new_AGEMA_signal_4859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2342 ( .C (clk), .D (new_AGEMA_signal_4862), .Q (new_AGEMA_signal_4863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2346 ( .C (clk), .D (new_AGEMA_signal_4866), .Q (new_AGEMA_signal_4867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2350 ( .C (clk), .D (new_AGEMA_signal_4870), .Q (new_AGEMA_signal_4871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2354 ( .C (clk), .D (new_AGEMA_signal_4874), .Q (new_AGEMA_signal_4875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2358 ( .C (clk), .D (new_AGEMA_signal_4878), .Q (new_AGEMA_signal_4879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2362 ( .C (clk), .D (new_AGEMA_signal_4882), .Q (new_AGEMA_signal_4883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2366 ( .C (clk), .D (new_AGEMA_signal_4886), .Q (new_AGEMA_signal_4887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2370 ( .C (clk), .D (new_AGEMA_signal_4890), .Q (new_AGEMA_signal_4891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2374 ( .C (clk), .D (new_AGEMA_signal_4894), .Q (new_AGEMA_signal_4895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2378 ( .C (clk), .D (new_AGEMA_signal_4898), .Q (new_AGEMA_signal_4899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2382 ( .C (clk), .D (new_AGEMA_signal_4902), .Q (new_AGEMA_signal_4903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2386 ( .C (clk), .D (new_AGEMA_signal_4906), .Q (new_AGEMA_signal_4907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2390 ( .C (clk), .D (new_AGEMA_signal_4910), .Q (new_AGEMA_signal_4911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2394 ( .C (clk), .D (new_AGEMA_signal_4914), .Q (new_AGEMA_signal_4915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2398 ( .C (clk), .D (new_AGEMA_signal_4918), .Q (new_AGEMA_signal_4919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2402 ( .C (clk), .D (new_AGEMA_signal_4922), .Q (new_AGEMA_signal_4923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2406 ( .C (clk), .D (new_AGEMA_signal_4926), .Q (new_AGEMA_signal_4927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2410 ( .C (clk), .D (new_AGEMA_signal_4930), .Q (new_AGEMA_signal_4931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2414 ( .C (clk), .D (new_AGEMA_signal_4934), .Q (new_AGEMA_signal_4935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2418 ( .C (clk), .D (new_AGEMA_signal_4938), .Q (new_AGEMA_signal_4939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2421 ( .C (clk), .D (new_AGEMA_signal_4941), .Q (new_AGEMA_signal_4942) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2424 ( .C (clk), .D (new_AGEMA_signal_4944), .Q (new_AGEMA_signal_4945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2427 ( .C (clk), .D (new_AGEMA_signal_4947), .Q (new_AGEMA_signal_4948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2430 ( .C (clk), .D (new_AGEMA_signal_4950), .Q (new_AGEMA_signal_4951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2433 ( .C (clk), .D (new_AGEMA_signal_4953), .Q (new_AGEMA_signal_4954) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2436 ( .C (clk), .D (new_AGEMA_signal_4956), .Q (new_AGEMA_signal_4957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2439 ( .C (clk), .D (new_AGEMA_signal_4959), .Q (new_AGEMA_signal_4960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2442 ( .C (clk), .D (new_AGEMA_signal_4962), .Q (new_AGEMA_signal_4963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2445 ( .C (clk), .D (new_AGEMA_signal_4965), .Q (new_AGEMA_signal_4966) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2448 ( .C (clk), .D (new_AGEMA_signal_4968), .Q (new_AGEMA_signal_4969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2451 ( .C (clk), .D (new_AGEMA_signal_4971), .Q (new_AGEMA_signal_4972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2454 ( .C (clk), .D (new_AGEMA_signal_4974), .Q (new_AGEMA_signal_4975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2457 ( .C (clk), .D (new_AGEMA_signal_4977), .Q (new_AGEMA_signal_4978) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2460 ( .C (clk), .D (new_AGEMA_signal_4980), .Q (new_AGEMA_signal_4981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2463 ( .C (clk), .D (new_AGEMA_signal_4983), .Q (new_AGEMA_signal_4984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2466 ( .C (clk), .D (new_AGEMA_signal_4986), .Q (new_AGEMA_signal_4987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2469 ( .C (clk), .D (new_AGEMA_signal_4989), .Q (new_AGEMA_signal_4990) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2472 ( .C (clk), .D (new_AGEMA_signal_4992), .Q (new_AGEMA_signal_4993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2475 ( .C (clk), .D (new_AGEMA_signal_4995), .Q (new_AGEMA_signal_4996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2478 ( .C (clk), .D (new_AGEMA_signal_4998), .Q (new_AGEMA_signal_4999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2481 ( .C (clk), .D (new_AGEMA_signal_5001), .Q (new_AGEMA_signal_5002) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2484 ( .C (clk), .D (new_AGEMA_signal_5004), .Q (new_AGEMA_signal_5005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2487 ( .C (clk), .D (new_AGEMA_signal_5007), .Q (new_AGEMA_signal_5008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2490 ( .C (clk), .D (new_AGEMA_signal_5010), .Q (new_AGEMA_signal_5011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2493 ( .C (clk), .D (new_AGEMA_signal_5013), .Q (new_AGEMA_signal_5014) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2496 ( .C (clk), .D (new_AGEMA_signal_5016), .Q (new_AGEMA_signal_5017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2499 ( .C (clk), .D (new_AGEMA_signal_5019), .Q (new_AGEMA_signal_5020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2502 ( .C (clk), .D (new_AGEMA_signal_5022), .Q (new_AGEMA_signal_5023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2505 ( .C (clk), .D (new_AGEMA_signal_5025), .Q (new_AGEMA_signal_5026) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2508 ( .C (clk), .D (new_AGEMA_signal_5028), .Q (new_AGEMA_signal_5029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2511 ( .C (clk), .D (new_AGEMA_signal_5031), .Q (new_AGEMA_signal_5032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2514 ( .C (clk), .D (new_AGEMA_signal_5034), .Q (new_AGEMA_signal_5035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2517 ( .C (clk), .D (new_AGEMA_signal_5037), .Q (new_AGEMA_signal_5038) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2520 ( .C (clk), .D (new_AGEMA_signal_5040), .Q (new_AGEMA_signal_5041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2523 ( .C (clk), .D (new_AGEMA_signal_5043), .Q (new_AGEMA_signal_5044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2526 ( .C (clk), .D (new_AGEMA_signal_5046), .Q (new_AGEMA_signal_5047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2529 ( .C (clk), .D (new_AGEMA_signal_5049), .Q (new_AGEMA_signal_5050) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2532 ( .C (clk), .D (new_AGEMA_signal_5052), .Q (new_AGEMA_signal_5053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2535 ( .C (clk), .D (new_AGEMA_signal_5055), .Q (new_AGEMA_signal_5056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2538 ( .C (clk), .D (new_AGEMA_signal_5058), .Q (new_AGEMA_signal_5059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2541 ( .C (clk), .D (new_AGEMA_signal_5061), .Q (new_AGEMA_signal_5062) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2544 ( .C (clk), .D (new_AGEMA_signal_5064), .Q (new_AGEMA_signal_5065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2547 ( .C (clk), .D (new_AGEMA_signal_5067), .Q (new_AGEMA_signal_5068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2550 ( .C (clk), .D (new_AGEMA_signal_5070), .Q (new_AGEMA_signal_5071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2553 ( .C (clk), .D (new_AGEMA_signal_5073), .Q (new_AGEMA_signal_5074) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2556 ( .C (clk), .D (new_AGEMA_signal_5076), .Q (new_AGEMA_signal_5077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2559 ( .C (clk), .D (new_AGEMA_signal_5079), .Q (new_AGEMA_signal_5080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2562 ( .C (clk), .D (new_AGEMA_signal_5082), .Q (new_AGEMA_signal_5083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2565 ( .C (clk), .D (new_AGEMA_signal_5085), .Q (new_AGEMA_signal_5086) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2568 ( .C (clk), .D (new_AGEMA_signal_5088), .Q (new_AGEMA_signal_5089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2571 ( .C (clk), .D (new_AGEMA_signal_5091), .Q (new_AGEMA_signal_5092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2574 ( .C (clk), .D (new_AGEMA_signal_5094), .Q (new_AGEMA_signal_5095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2577 ( .C (clk), .D (new_AGEMA_signal_5097), .Q (new_AGEMA_signal_5098) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2580 ( .C (clk), .D (new_AGEMA_signal_5100), .Q (new_AGEMA_signal_5101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2583 ( .C (clk), .D (new_AGEMA_signal_5103), .Q (new_AGEMA_signal_5104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2586 ( .C (clk), .D (new_AGEMA_signal_5106), .Q (new_AGEMA_signal_5107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2589 ( .C (clk), .D (new_AGEMA_signal_5109), .Q (new_AGEMA_signal_5110) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2592 ( .C (clk), .D (new_AGEMA_signal_5112), .Q (new_AGEMA_signal_5113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2595 ( .C (clk), .D (new_AGEMA_signal_5115), .Q (new_AGEMA_signal_5116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2598 ( .C (clk), .D (new_AGEMA_signal_5118), .Q (new_AGEMA_signal_5119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2601 ( .C (clk), .D (new_AGEMA_signal_5121), .Q (new_AGEMA_signal_5122) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2604 ( .C (clk), .D (new_AGEMA_signal_5124), .Q (new_AGEMA_signal_5125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2607 ( .C (clk), .D (new_AGEMA_signal_5127), .Q (new_AGEMA_signal_5128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2610 ( .C (clk), .D (new_AGEMA_signal_5130), .Q (new_AGEMA_signal_5131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2613 ( .C (clk), .D (new_AGEMA_signal_5133), .Q (new_AGEMA_signal_5134) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2616 ( .C (clk), .D (new_AGEMA_signal_5136), .Q (new_AGEMA_signal_5137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2619 ( .C (clk), .D (new_AGEMA_signal_5139), .Q (new_AGEMA_signal_5140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2622 ( .C (clk), .D (new_AGEMA_signal_5142), .Q (new_AGEMA_signal_5143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2625 ( .C (clk), .D (new_AGEMA_signal_5145), .Q (new_AGEMA_signal_5146) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2628 ( .C (clk), .D (new_AGEMA_signal_5148), .Q (new_AGEMA_signal_5149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2631 ( .C (clk), .D (new_AGEMA_signal_5151), .Q (new_AGEMA_signal_5152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2634 ( .C (clk), .D (new_AGEMA_signal_5154), .Q (new_AGEMA_signal_5155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2637 ( .C (clk), .D (new_AGEMA_signal_5157), .Q (new_AGEMA_signal_5158) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2640 ( .C (clk), .D (new_AGEMA_signal_5160), .Q (new_AGEMA_signal_5161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2643 ( .C (clk), .D (new_AGEMA_signal_5163), .Q (new_AGEMA_signal_5164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2646 ( .C (clk), .D (new_AGEMA_signal_5166), .Q (new_AGEMA_signal_5167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2649 ( .C (clk), .D (new_AGEMA_signal_5169), .Q (new_AGEMA_signal_5170) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2652 ( .C (clk), .D (new_AGEMA_signal_5172), .Q (new_AGEMA_signal_5173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2655 ( .C (clk), .D (new_AGEMA_signal_5175), .Q (new_AGEMA_signal_5176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2658 ( .C (clk), .D (new_AGEMA_signal_5178), .Q (new_AGEMA_signal_5179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2661 ( .C (clk), .D (new_AGEMA_signal_5181), .Q (new_AGEMA_signal_5182) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2664 ( .C (clk), .D (new_AGEMA_signal_5184), .Q (new_AGEMA_signal_5185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2667 ( .C (clk), .D (new_AGEMA_signal_5187), .Q (new_AGEMA_signal_5188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2670 ( .C (clk), .D (new_AGEMA_signal_5190), .Q (new_AGEMA_signal_5191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2673 ( .C (clk), .D (new_AGEMA_signal_5193), .Q (new_AGEMA_signal_5194) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2676 ( .C (clk), .D (new_AGEMA_signal_5196), .Q (new_AGEMA_signal_5197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2679 ( .C (clk), .D (new_AGEMA_signal_5199), .Q (new_AGEMA_signal_5200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2682 ( .C (clk), .D (new_AGEMA_signal_5202), .Q (new_AGEMA_signal_5203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2685 ( .C (clk), .D (new_AGEMA_signal_5205), .Q (new_AGEMA_signal_5206) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2688 ( .C (clk), .D (new_AGEMA_signal_5208), .Q (new_AGEMA_signal_5209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2691 ( .C (clk), .D (new_AGEMA_signal_5211), .Q (new_AGEMA_signal_5212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2694 ( .C (clk), .D (new_AGEMA_signal_5214), .Q (new_AGEMA_signal_5215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2697 ( .C (clk), .D (new_AGEMA_signal_5217), .Q (new_AGEMA_signal_5218) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2700 ( .C (clk), .D (new_AGEMA_signal_5220), .Q (new_AGEMA_signal_5221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2703 ( .C (clk), .D (new_AGEMA_signal_5223), .Q (new_AGEMA_signal_5224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2706 ( .C (clk), .D (new_AGEMA_signal_5226), .Q (new_AGEMA_signal_5227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2709 ( .C (clk), .D (new_AGEMA_signal_5229), .Q (new_AGEMA_signal_5230) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2712 ( .C (clk), .D (new_AGEMA_signal_5232), .Q (new_AGEMA_signal_5233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2715 ( .C (clk), .D (new_AGEMA_signal_5235), .Q (new_AGEMA_signal_5236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2718 ( .C (clk), .D (new_AGEMA_signal_5238), .Q (new_AGEMA_signal_5239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2721 ( .C (clk), .D (new_AGEMA_signal_5241), .Q (new_AGEMA_signal_5242) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2724 ( .C (clk), .D (new_AGEMA_signal_5244), .Q (new_AGEMA_signal_5245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2727 ( .C (clk), .D (new_AGEMA_signal_5247), .Q (new_AGEMA_signal_5248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2730 ( .C (clk), .D (new_AGEMA_signal_5250), .Q (new_AGEMA_signal_5251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2733 ( .C (clk), .D (new_AGEMA_signal_5253), .Q (new_AGEMA_signal_5254) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2736 ( .C (clk), .D (new_AGEMA_signal_5256), .Q (new_AGEMA_signal_5257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2739 ( .C (clk), .D (new_AGEMA_signal_5259), .Q (new_AGEMA_signal_5260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2742 ( .C (clk), .D (new_AGEMA_signal_5262), .Q (new_AGEMA_signal_5263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2745 ( .C (clk), .D (new_AGEMA_signal_5265), .Q (new_AGEMA_signal_5266) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2748 ( .C (clk), .D (new_AGEMA_signal_5268), .Q (new_AGEMA_signal_5269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2751 ( .C (clk), .D (new_AGEMA_signal_5271), .Q (new_AGEMA_signal_5272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2754 ( .C (clk), .D (new_AGEMA_signal_5274), .Q (new_AGEMA_signal_5275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2757 ( .C (clk), .D (new_AGEMA_signal_5277), .Q (new_AGEMA_signal_5278) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2760 ( .C (clk), .D (new_AGEMA_signal_5280), .Q (new_AGEMA_signal_5281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2763 ( .C (clk), .D (new_AGEMA_signal_5283), .Q (new_AGEMA_signal_5284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2766 ( .C (clk), .D (new_AGEMA_signal_5286), .Q (new_AGEMA_signal_5287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2769 ( .C (clk), .D (new_AGEMA_signal_5289), .Q (new_AGEMA_signal_5290) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2772 ( .C (clk), .D (new_AGEMA_signal_5292), .Q (new_AGEMA_signal_5293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2775 ( .C (clk), .D (new_AGEMA_signal_5295), .Q (new_AGEMA_signal_5296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2778 ( .C (clk), .D (new_AGEMA_signal_5298), .Q (new_AGEMA_signal_5299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2781 ( .C (clk), .D (new_AGEMA_signal_5301), .Q (new_AGEMA_signal_5302) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2784 ( .C (clk), .D (new_AGEMA_signal_5304), .Q (new_AGEMA_signal_5305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2787 ( .C (clk), .D (new_AGEMA_signal_5307), .Q (new_AGEMA_signal_5308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2790 ( .C (clk), .D (new_AGEMA_signal_5310), .Q (new_AGEMA_signal_5311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2793 ( .C (clk), .D (new_AGEMA_signal_5313), .Q (new_AGEMA_signal_5314) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2796 ( .C (clk), .D (new_AGEMA_signal_5316), .Q (new_AGEMA_signal_5317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2799 ( .C (clk), .D (new_AGEMA_signal_5319), .Q (new_AGEMA_signal_5320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2802 ( .C (clk), .D (new_AGEMA_signal_5322), .Q (new_AGEMA_signal_5323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2805 ( .C (clk), .D (new_AGEMA_signal_5325), .Q (new_AGEMA_signal_5326) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2808 ( .C (clk), .D (new_AGEMA_signal_5328), .Q (new_AGEMA_signal_5329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2811 ( .C (clk), .D (new_AGEMA_signal_5331), .Q (new_AGEMA_signal_5332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2814 ( .C (clk), .D (new_AGEMA_signal_5334), .Q (new_AGEMA_signal_5335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2817 ( .C (clk), .D (new_AGEMA_signal_5337), .Q (new_AGEMA_signal_5338) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2820 ( .C (clk), .D (new_AGEMA_signal_5340), .Q (new_AGEMA_signal_5341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2823 ( .C (clk), .D (new_AGEMA_signal_5343), .Q (new_AGEMA_signal_5344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2826 ( .C (clk), .D (new_AGEMA_signal_5346), .Q (new_AGEMA_signal_5347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2829 ( .C (clk), .D (new_AGEMA_signal_5349), .Q (new_AGEMA_signal_5350) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2832 ( .C (clk), .D (new_AGEMA_signal_5352), .Q (new_AGEMA_signal_5353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2835 ( .C (clk), .D (new_AGEMA_signal_5355), .Q (new_AGEMA_signal_5356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2838 ( .C (clk), .D (new_AGEMA_signal_5358), .Q (new_AGEMA_signal_5359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2841 ( .C (clk), .D (new_AGEMA_signal_5361), .Q (new_AGEMA_signal_5362) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2844 ( .C (clk), .D (new_AGEMA_signal_5364), .Q (new_AGEMA_signal_5365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2847 ( .C (clk), .D (new_AGEMA_signal_5367), .Q (new_AGEMA_signal_5368) ) ;
    buf_clk new_AGEMA_reg_buffer_2850 ( .C (clk), .D (new_AGEMA_signal_5370), .Q (new_AGEMA_signal_5371) ) ;
    buf_clk new_AGEMA_reg_buffer_2854 ( .C (clk), .D (new_AGEMA_signal_5374), .Q (new_AGEMA_signal_5375) ) ;
    buf_clk new_AGEMA_reg_buffer_2858 ( .C (clk), .D (new_AGEMA_signal_5378), .Q (new_AGEMA_signal_5379) ) ;
    buf_clk new_AGEMA_reg_buffer_2862 ( .C (clk), .D (new_AGEMA_signal_5382), .Q (new_AGEMA_signal_5383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2866 ( .C (clk), .D (new_AGEMA_signal_5386), .Q (new_AGEMA_signal_5387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2870 ( .C (clk), .D (new_AGEMA_signal_5390), .Q (new_AGEMA_signal_5391) ) ;
    buf_clk new_AGEMA_reg_buffer_2874 ( .C (clk), .D (new_AGEMA_signal_5394), .Q (new_AGEMA_signal_5395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2878 ( .C (clk), .D (new_AGEMA_signal_5398), .Q (new_AGEMA_signal_5399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2882 ( .C (clk), .D (new_AGEMA_signal_5402), .Q (new_AGEMA_signal_5403) ) ;
    buf_clk new_AGEMA_reg_buffer_2886 ( .C (clk), .D (new_AGEMA_signal_5406), .Q (new_AGEMA_signal_5407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2890 ( .C (clk), .D (new_AGEMA_signal_5410), .Q (new_AGEMA_signal_5411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2894 ( .C (clk), .D (new_AGEMA_signal_5414), .Q (new_AGEMA_signal_5415) ) ;
    buf_clk new_AGEMA_reg_buffer_2898 ( .C (clk), .D (new_AGEMA_signal_5418), .Q (new_AGEMA_signal_5419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2902 ( .C (clk), .D (new_AGEMA_signal_5422), .Q (new_AGEMA_signal_5423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2906 ( .C (clk), .D (new_AGEMA_signal_5426), .Q (new_AGEMA_signal_5427) ) ;
    buf_clk new_AGEMA_reg_buffer_2910 ( .C (clk), .D (new_AGEMA_signal_5430), .Q (new_AGEMA_signal_5431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2914 ( .C (clk), .D (new_AGEMA_signal_5434), .Q (new_AGEMA_signal_5435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2918 ( .C (clk), .D (new_AGEMA_signal_5438), .Q (new_AGEMA_signal_5439) ) ;
    buf_clk new_AGEMA_reg_buffer_2922 ( .C (clk), .D (new_AGEMA_signal_5442), .Q (new_AGEMA_signal_5443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2926 ( .C (clk), .D (new_AGEMA_signal_5446), .Q (new_AGEMA_signal_5447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2930 ( .C (clk), .D (new_AGEMA_signal_5450), .Q (new_AGEMA_signal_5451) ) ;
    buf_clk new_AGEMA_reg_buffer_2934 ( .C (clk), .D (new_AGEMA_signal_5454), .Q (new_AGEMA_signal_5455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2938 ( .C (clk), .D (new_AGEMA_signal_5458), .Q (new_AGEMA_signal_5459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2942 ( .C (clk), .D (new_AGEMA_signal_5462), .Q (new_AGEMA_signal_5463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2946 ( .C (clk), .D (new_AGEMA_signal_5466), .Q (new_AGEMA_signal_5467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2950 ( .C (clk), .D (new_AGEMA_signal_5470), .Q (new_AGEMA_signal_5471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2954 ( .C (clk), .D (new_AGEMA_signal_5474), .Q (new_AGEMA_signal_5475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2958 ( .C (clk), .D (new_AGEMA_signal_5478), .Q (new_AGEMA_signal_5479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2962 ( .C (clk), .D (new_AGEMA_signal_5482), .Q (new_AGEMA_signal_5483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2966 ( .C (clk), .D (new_AGEMA_signal_5486), .Q (new_AGEMA_signal_5487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2970 ( .C (clk), .D (new_AGEMA_signal_5490), .Q (new_AGEMA_signal_5491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2974 ( .C (clk), .D (new_AGEMA_signal_5494), .Q (new_AGEMA_signal_5495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2978 ( .C (clk), .D (new_AGEMA_signal_5498), .Q (new_AGEMA_signal_5499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2982 ( .C (clk), .D (new_AGEMA_signal_5502), .Q (new_AGEMA_signal_5503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2986 ( .C (clk), .D (new_AGEMA_signal_5506), .Q (new_AGEMA_signal_5507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2990 ( .C (clk), .D (new_AGEMA_signal_5510), .Q (new_AGEMA_signal_5511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2994 ( .C (clk), .D (new_AGEMA_signal_5514), .Q (new_AGEMA_signal_5515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2998 ( .C (clk), .D (new_AGEMA_signal_5518), .Q (new_AGEMA_signal_5519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3002 ( .C (clk), .D (new_AGEMA_signal_5522), .Q (new_AGEMA_signal_5523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3006 ( .C (clk), .D (new_AGEMA_signal_5526), .Q (new_AGEMA_signal_5527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3010 ( .C (clk), .D (new_AGEMA_signal_5530), .Q (new_AGEMA_signal_5531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3014 ( .C (clk), .D (new_AGEMA_signal_5534), .Q (new_AGEMA_signal_5535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3018 ( .C (clk), .D (new_AGEMA_signal_5538), .Q (new_AGEMA_signal_5539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3022 ( .C (clk), .D (new_AGEMA_signal_5542), .Q (new_AGEMA_signal_5543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3026 ( .C (clk), .D (new_AGEMA_signal_5546), .Q (new_AGEMA_signal_5547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3030 ( .C (clk), .D (new_AGEMA_signal_5550), .Q (new_AGEMA_signal_5551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3034 ( .C (clk), .D (new_AGEMA_signal_5554), .Q (new_AGEMA_signal_5555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3038 ( .C (clk), .D (new_AGEMA_signal_5558), .Q (new_AGEMA_signal_5559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3042 ( .C (clk), .D (new_AGEMA_signal_5562), .Q (new_AGEMA_signal_5563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3046 ( .C (clk), .D (new_AGEMA_signal_5566), .Q (new_AGEMA_signal_5567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3050 ( .C (clk), .D (new_AGEMA_signal_5570), .Q (new_AGEMA_signal_5571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3054 ( .C (clk), .D (new_AGEMA_signal_5574), .Q (new_AGEMA_signal_5575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3058 ( .C (clk), .D (new_AGEMA_signal_5578), .Q (new_AGEMA_signal_5579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3062 ( .C (clk), .D (new_AGEMA_signal_5582), .Q (new_AGEMA_signal_5583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3066 ( .C (clk), .D (new_AGEMA_signal_5586), .Q (new_AGEMA_signal_5587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3070 ( .C (clk), .D (new_AGEMA_signal_5590), .Q (new_AGEMA_signal_5591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3074 ( .C (clk), .D (new_AGEMA_signal_5594), .Q (new_AGEMA_signal_5595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3078 ( .C (clk), .D (new_AGEMA_signal_5598), .Q (new_AGEMA_signal_5599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3082 ( .C (clk), .D (new_AGEMA_signal_5602), .Q (new_AGEMA_signal_5603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3086 ( .C (clk), .D (new_AGEMA_signal_5606), .Q (new_AGEMA_signal_5607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3090 ( .C (clk), .D (new_AGEMA_signal_5610), .Q (new_AGEMA_signal_5611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3094 ( .C (clk), .D (new_AGEMA_signal_5614), .Q (new_AGEMA_signal_5615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3098 ( .C (clk), .D (new_AGEMA_signal_5618), .Q (new_AGEMA_signal_5619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3102 ( .C (clk), .D (new_AGEMA_signal_5622), .Q (new_AGEMA_signal_5623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3106 ( .C (clk), .D (new_AGEMA_signal_5626), .Q (new_AGEMA_signal_5627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3110 ( .C (clk), .D (new_AGEMA_signal_5630), .Q (new_AGEMA_signal_5631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3114 ( .C (clk), .D (new_AGEMA_signal_5634), .Q (new_AGEMA_signal_5635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3118 ( .C (clk), .D (new_AGEMA_signal_5638), .Q (new_AGEMA_signal_5639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3122 ( .C (clk), .D (new_AGEMA_signal_5642), .Q (new_AGEMA_signal_5643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3126 ( .C (clk), .D (new_AGEMA_signal_5646), .Q (new_AGEMA_signal_5647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3130 ( .C (clk), .D (new_AGEMA_signal_5650), .Q (new_AGEMA_signal_5651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3134 ( .C (clk), .D (new_AGEMA_signal_5654), .Q (new_AGEMA_signal_5655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3138 ( .C (clk), .D (new_AGEMA_signal_5658), .Q (new_AGEMA_signal_5659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3142 ( .C (clk), .D (new_AGEMA_signal_5662), .Q (new_AGEMA_signal_5663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3146 ( .C (clk), .D (new_AGEMA_signal_5666), .Q (new_AGEMA_signal_5667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3150 ( .C (clk), .D (new_AGEMA_signal_5670), .Q (new_AGEMA_signal_5671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3154 ( .C (clk), .D (new_AGEMA_signal_5674), .Q (new_AGEMA_signal_5675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3158 ( .C (clk), .D (new_AGEMA_signal_5678), .Q (new_AGEMA_signal_5679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3162 ( .C (clk), .D (new_AGEMA_signal_5682), .Q (new_AGEMA_signal_5683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3166 ( .C (clk), .D (new_AGEMA_signal_5686), .Q (new_AGEMA_signal_5687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3170 ( .C (clk), .D (new_AGEMA_signal_5690), .Q (new_AGEMA_signal_5691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3174 ( .C (clk), .D (new_AGEMA_signal_5694), .Q (new_AGEMA_signal_5695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3178 ( .C (clk), .D (new_AGEMA_signal_5698), .Q (new_AGEMA_signal_5699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3182 ( .C (clk), .D (new_AGEMA_signal_5702), .Q (new_AGEMA_signal_5703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3186 ( .C (clk), .D (new_AGEMA_signal_5706), .Q (new_AGEMA_signal_5707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3190 ( .C (clk), .D (new_AGEMA_signal_5710), .Q (new_AGEMA_signal_5711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3194 ( .C (clk), .D (new_AGEMA_signal_5714), .Q (new_AGEMA_signal_5715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3198 ( .C (clk), .D (new_AGEMA_signal_5718), .Q (new_AGEMA_signal_5719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3202 ( .C (clk), .D (new_AGEMA_signal_5722), .Q (new_AGEMA_signal_5723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3206 ( .C (clk), .D (new_AGEMA_signal_5726), .Q (new_AGEMA_signal_5727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3210 ( .C (clk), .D (new_AGEMA_signal_5730), .Q (new_AGEMA_signal_5731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3214 ( .C (clk), .D (new_AGEMA_signal_5734), .Q (new_AGEMA_signal_5735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3218 ( .C (clk), .D (new_AGEMA_signal_5738), .Q (new_AGEMA_signal_5739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3222 ( .C (clk), .D (new_AGEMA_signal_5742), .Q (new_AGEMA_signal_5743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3226 ( .C (clk), .D (new_AGEMA_signal_5746), .Q (new_AGEMA_signal_5747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3230 ( .C (clk), .D (new_AGEMA_signal_5750), .Q (new_AGEMA_signal_5751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3234 ( .C (clk), .D (new_AGEMA_signal_5754), .Q (new_AGEMA_signal_5755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3238 ( .C (clk), .D (new_AGEMA_signal_5758), .Q (new_AGEMA_signal_5759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3242 ( .C (clk), .D (new_AGEMA_signal_5762), .Q (new_AGEMA_signal_5763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3246 ( .C (clk), .D (new_AGEMA_signal_5766), .Q (new_AGEMA_signal_5767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3250 ( .C (clk), .D (new_AGEMA_signal_5770), .Q (new_AGEMA_signal_5771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3254 ( .C (clk), .D (new_AGEMA_signal_5774), .Q (new_AGEMA_signal_5775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3258 ( .C (clk), .D (new_AGEMA_signal_5778), .Q (new_AGEMA_signal_5779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3262 ( .C (clk), .D (new_AGEMA_signal_5782), .Q (new_AGEMA_signal_5783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3266 ( .C (clk), .D (new_AGEMA_signal_5786), .Q (new_AGEMA_signal_5787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3270 ( .C (clk), .D (new_AGEMA_signal_5790), .Q (new_AGEMA_signal_5791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3274 ( .C (clk), .D (new_AGEMA_signal_5794), .Q (new_AGEMA_signal_5795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3278 ( .C (clk), .D (new_AGEMA_signal_5798), .Q (new_AGEMA_signal_5799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3282 ( .C (clk), .D (new_AGEMA_signal_5802), .Q (new_AGEMA_signal_5803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3286 ( .C (clk), .D (new_AGEMA_signal_5806), .Q (new_AGEMA_signal_5807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3290 ( .C (clk), .D (new_AGEMA_signal_5810), .Q (new_AGEMA_signal_5811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3294 ( .C (clk), .D (new_AGEMA_signal_5814), .Q (new_AGEMA_signal_5815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3298 ( .C (clk), .D (new_AGEMA_signal_5818), .Q (new_AGEMA_signal_5819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3302 ( .C (clk), .D (new_AGEMA_signal_5822), .Q (new_AGEMA_signal_5823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3306 ( .C (clk), .D (new_AGEMA_signal_5826), .Q (new_AGEMA_signal_5827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3310 ( .C (clk), .D (new_AGEMA_signal_5830), .Q (new_AGEMA_signal_5831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3314 ( .C (clk), .D (new_AGEMA_signal_5834), .Q (new_AGEMA_signal_5835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3318 ( .C (clk), .D (new_AGEMA_signal_5838), .Q (new_AGEMA_signal_5839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3322 ( .C (clk), .D (new_AGEMA_signal_5842), .Q (new_AGEMA_signal_5843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3326 ( .C (clk), .D (new_AGEMA_signal_5846), .Q (new_AGEMA_signal_5847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3330 ( .C (clk), .D (new_AGEMA_signal_5850), .Q (new_AGEMA_signal_5851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3334 ( .C (clk), .D (new_AGEMA_signal_5854), .Q (new_AGEMA_signal_5855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3338 ( .C (clk), .D (new_AGEMA_signal_5858), .Q (new_AGEMA_signal_5859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3342 ( .C (clk), .D (new_AGEMA_signal_5862), .Q (new_AGEMA_signal_5863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3346 ( .C (clk), .D (new_AGEMA_signal_5866), .Q (new_AGEMA_signal_5867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3350 ( .C (clk), .D (new_AGEMA_signal_5870), .Q (new_AGEMA_signal_5871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3354 ( .C (clk), .D (new_AGEMA_signal_5874), .Q (new_AGEMA_signal_5875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3358 ( .C (clk), .D (new_AGEMA_signal_5878), .Q (new_AGEMA_signal_5879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3362 ( .C (clk), .D (new_AGEMA_signal_5882), .Q (new_AGEMA_signal_5883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3366 ( .C (clk), .D (new_AGEMA_signal_5886), .Q (new_AGEMA_signal_5887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3370 ( .C (clk), .D (new_AGEMA_signal_5890), .Q (new_AGEMA_signal_5891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3374 ( .C (clk), .D (new_AGEMA_signal_5894), .Q (new_AGEMA_signal_5895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3378 ( .C (clk), .D (new_AGEMA_signal_5898), .Q (new_AGEMA_signal_5899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3382 ( .C (clk), .D (new_AGEMA_signal_5902), .Q (new_AGEMA_signal_5903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3386 ( .C (clk), .D (new_AGEMA_signal_5906), .Q (new_AGEMA_signal_5907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3390 ( .C (clk), .D (new_AGEMA_signal_5910), .Q (new_AGEMA_signal_5911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3394 ( .C (clk), .D (new_AGEMA_signal_5914), .Q (new_AGEMA_signal_5915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3398 ( .C (clk), .D (new_AGEMA_signal_5918), .Q (new_AGEMA_signal_5919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3402 ( .C (clk), .D (new_AGEMA_signal_5922), .Q (new_AGEMA_signal_5923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3406 ( .C (clk), .D (new_AGEMA_signal_5926), .Q (new_AGEMA_signal_5927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3410 ( .C (clk), .D (new_AGEMA_signal_5930), .Q (new_AGEMA_signal_5931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3414 ( .C (clk), .D (new_AGEMA_signal_5934), .Q (new_AGEMA_signal_5935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3418 ( .C (clk), .D (new_AGEMA_signal_5938), .Q (new_AGEMA_signal_5939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3422 ( .C (clk), .D (new_AGEMA_signal_5942), .Q (new_AGEMA_signal_5943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3426 ( .C (clk), .D (new_AGEMA_signal_5946), .Q (new_AGEMA_signal_5947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3430 ( .C (clk), .D (new_AGEMA_signal_5950), .Q (new_AGEMA_signal_5951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3434 ( .C (clk), .D (new_AGEMA_signal_5954), .Q (new_AGEMA_signal_5955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3438 ( .C (clk), .D (new_AGEMA_signal_5958), .Q (new_AGEMA_signal_5959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3442 ( .C (clk), .D (new_AGEMA_signal_5962), .Q (new_AGEMA_signal_5963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3446 ( .C (clk), .D (new_AGEMA_signal_5966), .Q (new_AGEMA_signal_5967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3450 ( .C (clk), .D (new_AGEMA_signal_5970), .Q (new_AGEMA_signal_5971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3454 ( .C (clk), .D (new_AGEMA_signal_5974), .Q (new_AGEMA_signal_5975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3458 ( .C (clk), .D (new_AGEMA_signal_5978), .Q (new_AGEMA_signal_5979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3462 ( .C (clk), .D (new_AGEMA_signal_5982), .Q (new_AGEMA_signal_5983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3466 ( .C (clk), .D (new_AGEMA_signal_5986), .Q (new_AGEMA_signal_5987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3470 ( .C (clk), .D (new_AGEMA_signal_5990), .Q (new_AGEMA_signal_5991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3474 ( .C (clk), .D (new_AGEMA_signal_5994), .Q (new_AGEMA_signal_5995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3478 ( .C (clk), .D (new_AGEMA_signal_5998), .Q (new_AGEMA_signal_5999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3482 ( .C (clk), .D (new_AGEMA_signal_6002), .Q (new_AGEMA_signal_6003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3486 ( .C (clk), .D (new_AGEMA_signal_6006), .Q (new_AGEMA_signal_6007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3490 ( .C (clk), .D (new_AGEMA_signal_6010), .Q (new_AGEMA_signal_6011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3494 ( .C (clk), .D (new_AGEMA_signal_6014), .Q (new_AGEMA_signal_6015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3498 ( .C (clk), .D (new_AGEMA_signal_6018), .Q (new_AGEMA_signal_6019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3502 ( .C (clk), .D (new_AGEMA_signal_6022), .Q (new_AGEMA_signal_6023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3506 ( .C (clk), .D (new_AGEMA_signal_6026), .Q (new_AGEMA_signal_6027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3510 ( .C (clk), .D (new_AGEMA_signal_6030), .Q (new_AGEMA_signal_6031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3514 ( .C (clk), .D (new_AGEMA_signal_6034), .Q (new_AGEMA_signal_6035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3518 ( .C (clk), .D (new_AGEMA_signal_6038), .Q (new_AGEMA_signal_6039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3522 ( .C (clk), .D (new_AGEMA_signal_6042), .Q (new_AGEMA_signal_6043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3526 ( .C (clk), .D (new_AGEMA_signal_6046), .Q (new_AGEMA_signal_6047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3530 ( .C (clk), .D (new_AGEMA_signal_6050), .Q (new_AGEMA_signal_6051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3534 ( .C (clk), .D (new_AGEMA_signal_6054), .Q (new_AGEMA_signal_6055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3538 ( .C (clk), .D (new_AGEMA_signal_6058), .Q (new_AGEMA_signal_6059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3542 ( .C (clk), .D (new_AGEMA_signal_6062), .Q (new_AGEMA_signal_6063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3546 ( .C (clk), .D (new_AGEMA_signal_6066), .Q (new_AGEMA_signal_6067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3550 ( .C (clk), .D (new_AGEMA_signal_6070), .Q (new_AGEMA_signal_6071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3554 ( .C (clk), .D (new_AGEMA_signal_6074), .Q (new_AGEMA_signal_6075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3558 ( .C (clk), .D (new_AGEMA_signal_6078), .Q (new_AGEMA_signal_6079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3562 ( .C (clk), .D (new_AGEMA_signal_6082), .Q (new_AGEMA_signal_6083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3566 ( .C (clk), .D (new_AGEMA_signal_6086), .Q (new_AGEMA_signal_6087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3570 ( .C (clk), .D (new_AGEMA_signal_6090), .Q (new_AGEMA_signal_6091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3574 ( .C (clk), .D (new_AGEMA_signal_6094), .Q (new_AGEMA_signal_6095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3578 ( .C (clk), .D (new_AGEMA_signal_6098), .Q (new_AGEMA_signal_6099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3582 ( .C (clk), .D (new_AGEMA_signal_6102), .Q (new_AGEMA_signal_6103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3586 ( .C (clk), .D (new_AGEMA_signal_6106), .Q (new_AGEMA_signal_6107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3590 ( .C (clk), .D (new_AGEMA_signal_6110), .Q (new_AGEMA_signal_6111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3594 ( .C (clk), .D (new_AGEMA_signal_6114), .Q (new_AGEMA_signal_6115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3598 ( .C (clk), .D (new_AGEMA_signal_6118), .Q (new_AGEMA_signal_6119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3602 ( .C (clk), .D (new_AGEMA_signal_6122), .Q (new_AGEMA_signal_6123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3606 ( .C (clk), .D (new_AGEMA_signal_6126), .Q (new_AGEMA_signal_6127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3610 ( .C (clk), .D (new_AGEMA_signal_6130), .Q (new_AGEMA_signal_6131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3614 ( .C (clk), .D (new_AGEMA_signal_6134), .Q (new_AGEMA_signal_6135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3618 ( .C (clk), .D (new_AGEMA_signal_6138), .Q (new_AGEMA_signal_6139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3622 ( .C (clk), .D (new_AGEMA_signal_6142), .Q (new_AGEMA_signal_6143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3626 ( .C (clk), .D (new_AGEMA_signal_6146), .Q (new_AGEMA_signal_6147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3630 ( .C (clk), .D (new_AGEMA_signal_6150), .Q (new_AGEMA_signal_6151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3634 ( .C (clk), .D (new_AGEMA_signal_6154), .Q (new_AGEMA_signal_6155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3638 ( .C (clk), .D (new_AGEMA_signal_6158), .Q (new_AGEMA_signal_6159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3642 ( .C (clk), .D (new_AGEMA_signal_6162), .Q (new_AGEMA_signal_6163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3646 ( .C (clk), .D (new_AGEMA_signal_6166), .Q (new_AGEMA_signal_6167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3650 ( .C (clk), .D (new_AGEMA_signal_6170), .Q (new_AGEMA_signal_6171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3654 ( .C (clk), .D (new_AGEMA_signal_6174), .Q (new_AGEMA_signal_6175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3658 ( .C (clk), .D (new_AGEMA_signal_6178), .Q (new_AGEMA_signal_6179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3662 ( .C (clk), .D (new_AGEMA_signal_6182), .Q (new_AGEMA_signal_6183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3666 ( .C (clk), .D (new_AGEMA_signal_6186), .Q (new_AGEMA_signal_6187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3670 ( .C (clk), .D (new_AGEMA_signal_6190), .Q (new_AGEMA_signal_6191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3674 ( .C (clk), .D (new_AGEMA_signal_6194), .Q (new_AGEMA_signal_6195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3678 ( .C (clk), .D (new_AGEMA_signal_6198), .Q (new_AGEMA_signal_6199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3682 ( .C (clk), .D (new_AGEMA_signal_6202), .Q (new_AGEMA_signal_6203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3686 ( .C (clk), .D (new_AGEMA_signal_6206), .Q (new_AGEMA_signal_6207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3690 ( .C (clk), .D (new_AGEMA_signal_6210), .Q (new_AGEMA_signal_6211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3694 ( .C (clk), .D (new_AGEMA_signal_6214), .Q (new_AGEMA_signal_6215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3698 ( .C (clk), .D (new_AGEMA_signal_6218), .Q (new_AGEMA_signal_6219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3702 ( .C (clk), .D (new_AGEMA_signal_6222), .Q (new_AGEMA_signal_6223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3706 ( .C (clk), .D (new_AGEMA_signal_6226), .Q (new_AGEMA_signal_6227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3710 ( .C (clk), .D (new_AGEMA_signal_6230), .Q (new_AGEMA_signal_6231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3714 ( .C (clk), .D (new_AGEMA_signal_6234), .Q (new_AGEMA_signal_6235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3718 ( .C (clk), .D (new_AGEMA_signal_6238), .Q (new_AGEMA_signal_6239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3722 ( .C (clk), .D (new_AGEMA_signal_6242), .Q (new_AGEMA_signal_6243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3726 ( .C (clk), .D (new_AGEMA_signal_6246), .Q (new_AGEMA_signal_6247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3730 ( .C (clk), .D (new_AGEMA_signal_6250), .Q (new_AGEMA_signal_6251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3734 ( .C (clk), .D (new_AGEMA_signal_6254), .Q (new_AGEMA_signal_6255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3738 ( .C (clk), .D (new_AGEMA_signal_6258), .Q (new_AGEMA_signal_6259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3742 ( .C (clk), .D (new_AGEMA_signal_6262), .Q (new_AGEMA_signal_6263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3746 ( .C (clk), .D (new_AGEMA_signal_6266), .Q (new_AGEMA_signal_6267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3750 ( .C (clk), .D (new_AGEMA_signal_6270), .Q (new_AGEMA_signal_6271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3754 ( .C (clk), .D (new_AGEMA_signal_6274), .Q (new_AGEMA_signal_6275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3758 ( .C (clk), .D (new_AGEMA_signal_6278), .Q (new_AGEMA_signal_6279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3762 ( .C (clk), .D (new_AGEMA_signal_6282), .Q (new_AGEMA_signal_6283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3766 ( .C (clk), .D (new_AGEMA_signal_6286), .Q (new_AGEMA_signal_6287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3770 ( .C (clk), .D (new_AGEMA_signal_6290), .Q (new_AGEMA_signal_6291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3774 ( .C (clk), .D (new_AGEMA_signal_6294), .Q (new_AGEMA_signal_6295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3778 ( .C (clk), .D (new_AGEMA_signal_6298), .Q (new_AGEMA_signal_6299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3782 ( .C (clk), .D (new_AGEMA_signal_6302), .Q (new_AGEMA_signal_6303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3786 ( .C (clk), .D (new_AGEMA_signal_6306), .Q (new_AGEMA_signal_6307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3790 ( .C (clk), .D (new_AGEMA_signal_6310), .Q (new_AGEMA_signal_6311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3794 ( .C (clk), .D (new_AGEMA_signal_6314), .Q (new_AGEMA_signal_6315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3798 ( .C (clk), .D (new_AGEMA_signal_6318), .Q (new_AGEMA_signal_6319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3802 ( .C (clk), .D (new_AGEMA_signal_6322), .Q (new_AGEMA_signal_6323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3806 ( .C (clk), .D (new_AGEMA_signal_6326), .Q (new_AGEMA_signal_6327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3810 ( .C (clk), .D (new_AGEMA_signal_6330), .Q (new_AGEMA_signal_6331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3814 ( .C (clk), .D (new_AGEMA_signal_6334), .Q (new_AGEMA_signal_6335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3818 ( .C (clk), .D (new_AGEMA_signal_6338), .Q (new_AGEMA_signal_6339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3822 ( .C (clk), .D (new_AGEMA_signal_6342), .Q (new_AGEMA_signal_6343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3826 ( .C (clk), .D (new_AGEMA_signal_6346), .Q (new_AGEMA_signal_6347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3830 ( .C (clk), .D (new_AGEMA_signal_6350), .Q (new_AGEMA_signal_6351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3834 ( .C (clk), .D (new_AGEMA_signal_6354), .Q (new_AGEMA_signal_6355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3838 ( .C (clk), .D (new_AGEMA_signal_6358), .Q (new_AGEMA_signal_6359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3842 ( .C (clk), .D (new_AGEMA_signal_6362), .Q (new_AGEMA_signal_6363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3846 ( .C (clk), .D (new_AGEMA_signal_6366), .Q (new_AGEMA_signal_6367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3850 ( .C (clk), .D (new_AGEMA_signal_6370), .Q (new_AGEMA_signal_6371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3854 ( .C (clk), .D (new_AGEMA_signal_6374), .Q (new_AGEMA_signal_6375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3858 ( .C (clk), .D (new_AGEMA_signal_6378), .Q (new_AGEMA_signal_6379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3862 ( .C (clk), .D (new_AGEMA_signal_6382), .Q (new_AGEMA_signal_6383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3866 ( .C (clk), .D (new_AGEMA_signal_6386), .Q (new_AGEMA_signal_6387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3870 ( .C (clk), .D (new_AGEMA_signal_6390), .Q (new_AGEMA_signal_6391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3874 ( .C (clk), .D (new_AGEMA_signal_6394), .Q (new_AGEMA_signal_6395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3878 ( .C (clk), .D (new_AGEMA_signal_6398), .Q (new_AGEMA_signal_6399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3882 ( .C (clk), .D (new_AGEMA_signal_6402), .Q (new_AGEMA_signal_6403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3886 ( .C (clk), .D (new_AGEMA_signal_6406), .Q (new_AGEMA_signal_6407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3890 ( .C (clk), .D (new_AGEMA_signal_6410), .Q (new_AGEMA_signal_6411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3894 ( .C (clk), .D (new_AGEMA_signal_6414), .Q (new_AGEMA_signal_6415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3898 ( .C (clk), .D (new_AGEMA_signal_6418), .Q (new_AGEMA_signal_6419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3902 ( .C (clk), .D (new_AGEMA_signal_6422), .Q (new_AGEMA_signal_6423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3906 ( .C (clk), .D (new_AGEMA_signal_6426), .Q (new_AGEMA_signal_6427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3910 ( .C (clk), .D (new_AGEMA_signal_6430), .Q (new_AGEMA_signal_6431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3914 ( .C (clk), .D (new_AGEMA_signal_6434), .Q (new_AGEMA_signal_6435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3918 ( .C (clk), .D (new_AGEMA_signal_6438), .Q (new_AGEMA_signal_6439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3922 ( .C (clk), .D (new_AGEMA_signal_6442), .Q (new_AGEMA_signal_6443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3926 ( .C (clk), .D (new_AGEMA_signal_6446), .Q (new_AGEMA_signal_6447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3930 ( .C (clk), .D (new_AGEMA_signal_6450), .Q (new_AGEMA_signal_6451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3934 ( .C (clk), .D (new_AGEMA_signal_6454), .Q (new_AGEMA_signal_6455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3938 ( .C (clk), .D (new_AGEMA_signal_6458), .Q (new_AGEMA_signal_6459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3942 ( .C (clk), .D (new_AGEMA_signal_6462), .Q (new_AGEMA_signal_6463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3946 ( .C (clk), .D (new_AGEMA_signal_6466), .Q (new_AGEMA_signal_6467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3950 ( .C (clk), .D (new_AGEMA_signal_6470), .Q (new_AGEMA_signal_6471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3954 ( .C (clk), .D (new_AGEMA_signal_6474), .Q (new_AGEMA_signal_6475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3958 ( .C (clk), .D (new_AGEMA_signal_6478), .Q (new_AGEMA_signal_6479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3962 ( .C (clk), .D (new_AGEMA_signal_6482), .Q (new_AGEMA_signal_6483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3966 ( .C (clk), .D (new_AGEMA_signal_6486), .Q (new_AGEMA_signal_6487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3970 ( .C (clk), .D (new_AGEMA_signal_6490), .Q (new_AGEMA_signal_6491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3974 ( .C (clk), .D (new_AGEMA_signal_6494), .Q (new_AGEMA_signal_6495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3978 ( .C (clk), .D (new_AGEMA_signal_6498), .Q (new_AGEMA_signal_6499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3982 ( .C (clk), .D (new_AGEMA_signal_6502), .Q (new_AGEMA_signal_6503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3986 ( .C (clk), .D (new_AGEMA_signal_6506), .Q (new_AGEMA_signal_6507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3990 ( .C (clk), .D (new_AGEMA_signal_6510), .Q (new_AGEMA_signal_6511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3994 ( .C (clk), .D (new_AGEMA_signal_6514), .Q (new_AGEMA_signal_6515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3998 ( .C (clk), .D (new_AGEMA_signal_6518), .Q (new_AGEMA_signal_6519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4002 ( .C (clk), .D (new_AGEMA_signal_6522), .Q (new_AGEMA_signal_6523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4006 ( .C (clk), .D (new_AGEMA_signal_6526), .Q (new_AGEMA_signal_6527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4010 ( .C (clk), .D (new_AGEMA_signal_6530), .Q (new_AGEMA_signal_6531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4014 ( .C (clk), .D (new_AGEMA_signal_6534), .Q (new_AGEMA_signal_6535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4018 ( .C (clk), .D (new_AGEMA_signal_6538), .Q (new_AGEMA_signal_6539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4022 ( .C (clk), .D (new_AGEMA_signal_6542), .Q (new_AGEMA_signal_6543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4026 ( .C (clk), .D (new_AGEMA_signal_6546), .Q (new_AGEMA_signal_6547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4030 ( .C (clk), .D (new_AGEMA_signal_6550), .Q (new_AGEMA_signal_6551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4034 ( .C (clk), .D (new_AGEMA_signal_6554), .Q (new_AGEMA_signal_6555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4038 ( .C (clk), .D (new_AGEMA_signal_6558), .Q (new_AGEMA_signal_6559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4042 ( .C (clk), .D (new_AGEMA_signal_6562), .Q (new_AGEMA_signal_6563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4046 ( .C (clk), .D (new_AGEMA_signal_6566), .Q (new_AGEMA_signal_6567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4050 ( .C (clk), .D (new_AGEMA_signal_6570), .Q (new_AGEMA_signal_6571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4054 ( .C (clk), .D (new_AGEMA_signal_6574), .Q (new_AGEMA_signal_6575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4058 ( .C (clk), .D (new_AGEMA_signal_6578), .Q (new_AGEMA_signal_6579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4062 ( .C (clk), .D (new_AGEMA_signal_6582), .Q (new_AGEMA_signal_6583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4066 ( .C (clk), .D (new_AGEMA_signal_6586), .Q (new_AGEMA_signal_6587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4070 ( .C (clk), .D (new_AGEMA_signal_6590), .Q (new_AGEMA_signal_6591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4074 ( .C (clk), .D (new_AGEMA_signal_6594), .Q (new_AGEMA_signal_6595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4078 ( .C (clk), .D (new_AGEMA_signal_6598), .Q (new_AGEMA_signal_6599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4082 ( .C (clk), .D (new_AGEMA_signal_6602), .Q (new_AGEMA_signal_6603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4086 ( .C (clk), .D (new_AGEMA_signal_6606), .Q (new_AGEMA_signal_6607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4090 ( .C (clk), .D (new_AGEMA_signal_6610), .Q (new_AGEMA_signal_6611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4094 ( .C (clk), .D (new_AGEMA_signal_6614), .Q (new_AGEMA_signal_6615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4098 ( .C (clk), .D (new_AGEMA_signal_6618), .Q (new_AGEMA_signal_6619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4102 ( .C (clk), .D (new_AGEMA_signal_6622), .Q (new_AGEMA_signal_6623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4106 ( .C (clk), .D (new_AGEMA_signal_6626), .Q (new_AGEMA_signal_6627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4110 ( .C (clk), .D (new_AGEMA_signal_6630), .Q (new_AGEMA_signal_6631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4114 ( .C (clk), .D (new_AGEMA_signal_6634), .Q (new_AGEMA_signal_6635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4118 ( .C (clk), .D (new_AGEMA_signal_6638), .Q (new_AGEMA_signal_6639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4122 ( .C (clk), .D (new_AGEMA_signal_6642), .Q (new_AGEMA_signal_6643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4126 ( .C (clk), .D (new_AGEMA_signal_6646), .Q (new_AGEMA_signal_6647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4130 ( .C (clk), .D (new_AGEMA_signal_6650), .Q (new_AGEMA_signal_6651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4134 ( .C (clk), .D (new_AGEMA_signal_6654), .Q (new_AGEMA_signal_6655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4138 ( .C (clk), .D (new_AGEMA_signal_6658), .Q (new_AGEMA_signal_6659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4142 ( .C (clk), .D (new_AGEMA_signal_6662), .Q (new_AGEMA_signal_6663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4146 ( .C (clk), .D (new_AGEMA_signal_6666), .Q (new_AGEMA_signal_6667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4150 ( .C (clk), .D (new_AGEMA_signal_6670), .Q (new_AGEMA_signal_6671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4154 ( .C (clk), .D (new_AGEMA_signal_6674), .Q (new_AGEMA_signal_6675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4158 ( .C (clk), .D (new_AGEMA_signal_6678), .Q (new_AGEMA_signal_6679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4162 ( .C (clk), .D (new_AGEMA_signal_6682), .Q (new_AGEMA_signal_6683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4166 ( .C (clk), .D (new_AGEMA_signal_6686), .Q (new_AGEMA_signal_6687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4170 ( .C (clk), .D (new_AGEMA_signal_6690), .Q (new_AGEMA_signal_6691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4174 ( .C (clk), .D (new_AGEMA_signal_6694), .Q (new_AGEMA_signal_6695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4178 ( .C (clk), .D (new_AGEMA_signal_6698), .Q (new_AGEMA_signal_6699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4182 ( .C (clk), .D (new_AGEMA_signal_6702), .Q (new_AGEMA_signal_6703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4186 ( .C (clk), .D (new_AGEMA_signal_6706), .Q (new_AGEMA_signal_6707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4190 ( .C (clk), .D (new_AGEMA_signal_6710), .Q (new_AGEMA_signal_6711) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4194 ( .C (clk), .D (new_AGEMA_signal_6714), .Q (new_AGEMA_signal_6715) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4198 ( .C (clk), .D (new_AGEMA_signal_6718), .Q (new_AGEMA_signal_6719) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4202 ( .C (clk), .D (new_AGEMA_signal_6722), .Q (new_AGEMA_signal_6723) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4206 ( .C (clk), .D (new_AGEMA_signal_6726), .Q (new_AGEMA_signal_6727) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4210 ( .C (clk), .D (new_AGEMA_signal_6730), .Q (new_AGEMA_signal_6731) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4214 ( .C (clk), .D (new_AGEMA_signal_6734), .Q (new_AGEMA_signal_6735) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4218 ( .C (clk), .D (new_AGEMA_signal_6738), .Q (new_AGEMA_signal_6739) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4222 ( .C (clk), .D (new_AGEMA_signal_6742), .Q (new_AGEMA_signal_6743) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4226 ( .C (clk), .D (new_AGEMA_signal_6746), .Q (new_AGEMA_signal_6747) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4230 ( .C (clk), .D (new_AGEMA_signal_6750), .Q (new_AGEMA_signal_6751) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4234 ( .C (clk), .D (new_AGEMA_signal_6754), .Q (new_AGEMA_signal_6755) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4238 ( .C (clk), .D (new_AGEMA_signal_6758), .Q (new_AGEMA_signal_6759) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4242 ( .C (clk), .D (new_AGEMA_signal_6762), .Q (new_AGEMA_signal_6763) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4246 ( .C (clk), .D (new_AGEMA_signal_6766), .Q (new_AGEMA_signal_6767) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4250 ( .C (clk), .D (new_AGEMA_signal_6770), .Q (new_AGEMA_signal_6771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4254 ( .C (clk), .D (new_AGEMA_signal_6774), .Q (new_AGEMA_signal_6775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4258 ( .C (clk), .D (new_AGEMA_signal_6778), .Q (new_AGEMA_signal_6779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4262 ( .C (clk), .D (new_AGEMA_signal_6782), .Q (new_AGEMA_signal_6783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4266 ( .C (clk), .D (new_AGEMA_signal_6786), .Q (new_AGEMA_signal_6787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4270 ( .C (clk), .D (new_AGEMA_signal_6790), .Q (new_AGEMA_signal_6791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4274 ( .C (clk), .D (new_AGEMA_signal_6794), .Q (new_AGEMA_signal_6795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4278 ( .C (clk), .D (new_AGEMA_signal_6798), .Q (new_AGEMA_signal_6799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4282 ( .C (clk), .D (new_AGEMA_signal_6802), .Q (new_AGEMA_signal_6803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4286 ( .C (clk), .D (new_AGEMA_signal_6806), .Q (new_AGEMA_signal_6807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4290 ( .C (clk), .D (new_AGEMA_signal_6810), .Q (new_AGEMA_signal_6811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4294 ( .C (clk), .D (new_AGEMA_signal_6814), .Q (new_AGEMA_signal_6815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4298 ( .C (clk), .D (new_AGEMA_signal_6818), .Q (new_AGEMA_signal_6819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4302 ( .C (clk), .D (new_AGEMA_signal_6822), .Q (new_AGEMA_signal_6823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4306 ( .C (clk), .D (new_AGEMA_signal_6826), .Q (new_AGEMA_signal_6827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4310 ( .C (clk), .D (new_AGEMA_signal_6830), .Q (new_AGEMA_signal_6831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4314 ( .C (clk), .D (new_AGEMA_signal_6834), .Q (new_AGEMA_signal_6835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4318 ( .C (clk), .D (new_AGEMA_signal_6838), .Q (new_AGEMA_signal_6839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4322 ( .C (clk), .D (new_AGEMA_signal_6842), .Q (new_AGEMA_signal_6843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4326 ( .C (clk), .D (new_AGEMA_signal_6846), .Q (new_AGEMA_signal_6847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4330 ( .C (clk), .D (new_AGEMA_signal_6850), .Q (new_AGEMA_signal_6851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4334 ( .C (clk), .D (new_AGEMA_signal_6854), .Q (new_AGEMA_signal_6855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4338 ( .C (clk), .D (new_AGEMA_signal_6858), .Q (new_AGEMA_signal_6859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4342 ( .C (clk), .D (new_AGEMA_signal_6862), .Q (new_AGEMA_signal_6863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4346 ( .C (clk), .D (new_AGEMA_signal_6866), .Q (new_AGEMA_signal_6867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4350 ( .C (clk), .D (new_AGEMA_signal_6870), .Q (new_AGEMA_signal_6871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4354 ( .C (clk), .D (new_AGEMA_signal_6874), .Q (new_AGEMA_signal_6875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4358 ( .C (clk), .D (new_AGEMA_signal_6878), .Q (new_AGEMA_signal_6879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4362 ( .C (clk), .D (new_AGEMA_signal_6882), .Q (new_AGEMA_signal_6883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4366 ( .C (clk), .D (new_AGEMA_signal_6886), .Q (new_AGEMA_signal_6887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4370 ( .C (clk), .D (new_AGEMA_signal_6890), .Q (new_AGEMA_signal_6891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4374 ( .C (clk), .D (new_AGEMA_signal_6894), .Q (new_AGEMA_signal_6895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4378 ( .C (clk), .D (new_AGEMA_signal_6898), .Q (new_AGEMA_signal_6899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4382 ( .C (clk), .D (new_AGEMA_signal_6902), .Q (new_AGEMA_signal_6903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4386 ( .C (clk), .D (new_AGEMA_signal_6906), .Q (new_AGEMA_signal_6907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4390 ( .C (clk), .D (new_AGEMA_signal_6910), .Q (new_AGEMA_signal_6911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4394 ( .C (clk), .D (new_AGEMA_signal_6914), .Q (new_AGEMA_signal_6915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4398 ( .C (clk), .D (new_AGEMA_signal_6918), .Q (new_AGEMA_signal_6919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4402 ( .C (clk), .D (new_AGEMA_signal_6922), .Q (new_AGEMA_signal_6923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4406 ( .C (clk), .D (new_AGEMA_signal_6926), .Q (new_AGEMA_signal_6927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4410 ( .C (clk), .D (new_AGEMA_signal_6930), .Q (new_AGEMA_signal_6931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4414 ( .C (clk), .D (new_AGEMA_signal_6934), .Q (new_AGEMA_signal_6935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4418 ( .C (clk), .D (new_AGEMA_signal_6938), .Q (new_AGEMA_signal_6939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4422 ( .C (clk), .D (new_AGEMA_signal_6942), .Q (new_AGEMA_signal_6943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4426 ( .C (clk), .D (new_AGEMA_signal_6946), .Q (new_AGEMA_signal_6947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4430 ( .C (clk), .D (new_AGEMA_signal_6950), .Q (new_AGEMA_signal_6951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4434 ( .C (clk), .D (new_AGEMA_signal_6954), .Q (new_AGEMA_signal_6955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4438 ( .C (clk), .D (new_AGEMA_signal_6958), .Q (new_AGEMA_signal_6959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4442 ( .C (clk), .D (new_AGEMA_signal_6962), .Q (new_AGEMA_signal_6963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4446 ( .C (clk), .D (new_AGEMA_signal_6966), .Q (new_AGEMA_signal_6967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4450 ( .C (clk), .D (new_AGEMA_signal_6970), .Q (new_AGEMA_signal_6971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4454 ( .C (clk), .D (new_AGEMA_signal_6974), .Q (new_AGEMA_signal_6975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4458 ( .C (clk), .D (new_AGEMA_signal_6978), .Q (new_AGEMA_signal_6979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4462 ( .C (clk), .D (new_AGEMA_signal_6982), .Q (new_AGEMA_signal_6983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4466 ( .C (clk), .D (new_AGEMA_signal_6986), .Q (new_AGEMA_signal_6987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4470 ( .C (clk), .D (new_AGEMA_signal_6990), .Q (new_AGEMA_signal_6991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4474 ( .C (clk), .D (new_AGEMA_signal_6994), .Q (new_AGEMA_signal_6995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4478 ( .C (clk), .D (new_AGEMA_signal_6998), .Q (new_AGEMA_signal_6999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4482 ( .C (clk), .D (new_AGEMA_signal_7002), .Q (new_AGEMA_signal_7003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4486 ( .C (clk), .D (new_AGEMA_signal_7006), .Q (new_AGEMA_signal_7007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4490 ( .C (clk), .D (new_AGEMA_signal_7010), .Q (new_AGEMA_signal_7011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4494 ( .C (clk), .D (new_AGEMA_signal_7014), .Q (new_AGEMA_signal_7015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4498 ( .C (clk), .D (new_AGEMA_signal_7018), .Q (new_AGEMA_signal_7019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4502 ( .C (clk), .D (new_AGEMA_signal_7022), .Q (new_AGEMA_signal_7023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4506 ( .C (clk), .D (new_AGEMA_signal_7026), .Q (new_AGEMA_signal_7027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4510 ( .C (clk), .D (new_AGEMA_signal_7030), .Q (new_AGEMA_signal_7031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4514 ( .C (clk), .D (new_AGEMA_signal_7034), .Q (new_AGEMA_signal_7035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4518 ( .C (clk), .D (new_AGEMA_signal_7038), .Q (new_AGEMA_signal_7039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4522 ( .C (clk), .D (new_AGEMA_signal_7042), .Q (new_AGEMA_signal_7043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4526 ( .C (clk), .D (new_AGEMA_signal_7046), .Q (new_AGEMA_signal_7047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4530 ( .C (clk), .D (new_AGEMA_signal_7050), .Q (new_AGEMA_signal_7051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4534 ( .C (clk), .D (new_AGEMA_signal_7054), .Q (new_AGEMA_signal_7055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4538 ( .C (clk), .D (new_AGEMA_signal_7058), .Q (new_AGEMA_signal_7059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4542 ( .C (clk), .D (new_AGEMA_signal_7062), .Q (new_AGEMA_signal_7063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4546 ( .C (clk), .D (new_AGEMA_signal_7066), .Q (new_AGEMA_signal_7067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4550 ( .C (clk), .D (new_AGEMA_signal_7070), .Q (new_AGEMA_signal_7071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4554 ( .C (clk), .D (new_AGEMA_signal_7074), .Q (new_AGEMA_signal_7075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4558 ( .C (clk), .D (new_AGEMA_signal_7078), .Q (new_AGEMA_signal_7079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4562 ( .C (clk), .D (new_AGEMA_signal_7082), .Q (new_AGEMA_signal_7083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4566 ( .C (clk), .D (new_AGEMA_signal_7086), .Q (new_AGEMA_signal_7087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4570 ( .C (clk), .D (new_AGEMA_signal_7090), .Q (new_AGEMA_signal_7091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4574 ( .C (clk), .D (new_AGEMA_signal_7094), .Q (new_AGEMA_signal_7095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4578 ( .C (clk), .D (new_AGEMA_signal_7098), .Q (new_AGEMA_signal_7099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4582 ( .C (clk), .D (new_AGEMA_signal_7102), .Q (new_AGEMA_signal_7103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4586 ( .C (clk), .D (new_AGEMA_signal_7106), .Q (new_AGEMA_signal_7107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4590 ( .C (clk), .D (new_AGEMA_signal_7110), .Q (new_AGEMA_signal_7111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4594 ( .C (clk), .D (new_AGEMA_signal_7114), .Q (new_AGEMA_signal_7115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4598 ( .C (clk), .D (new_AGEMA_signal_7118), .Q (new_AGEMA_signal_7119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4602 ( .C (clk), .D (new_AGEMA_signal_7122), .Q (new_AGEMA_signal_7123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4606 ( .C (clk), .D (new_AGEMA_signal_7126), .Q (new_AGEMA_signal_7127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4610 ( .C (clk), .D (new_AGEMA_signal_7130), .Q (new_AGEMA_signal_7131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4614 ( .C (clk), .D (new_AGEMA_signal_7134), .Q (new_AGEMA_signal_7135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4618 ( .C (clk), .D (new_AGEMA_signal_7138), .Q (new_AGEMA_signal_7139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4622 ( .C (clk), .D (new_AGEMA_signal_7142), .Q (new_AGEMA_signal_7143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4626 ( .C (clk), .D (new_AGEMA_signal_7146), .Q (new_AGEMA_signal_7147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4630 ( .C (clk), .D (new_AGEMA_signal_7150), .Q (new_AGEMA_signal_7151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4634 ( .C (clk), .D (new_AGEMA_signal_7154), .Q (new_AGEMA_signal_7155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4638 ( .C (clk), .D (new_AGEMA_signal_7158), .Q (new_AGEMA_signal_7159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4642 ( .C (clk), .D (new_AGEMA_signal_7162), .Q (new_AGEMA_signal_7163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4646 ( .C (clk), .D (new_AGEMA_signal_7166), .Q (new_AGEMA_signal_7167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4650 ( .C (clk), .D (new_AGEMA_signal_7170), .Q (new_AGEMA_signal_7171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4654 ( .C (clk), .D (new_AGEMA_signal_7174), .Q (new_AGEMA_signal_7175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4658 ( .C (clk), .D (new_AGEMA_signal_7178), .Q (new_AGEMA_signal_7179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4662 ( .C (clk), .D (new_AGEMA_signal_7182), .Q (new_AGEMA_signal_7183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4666 ( .C (clk), .D (new_AGEMA_signal_7186), .Q (new_AGEMA_signal_7187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4670 ( .C (clk), .D (new_AGEMA_signal_7190), .Q (new_AGEMA_signal_7191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4674 ( .C (clk), .D (new_AGEMA_signal_7194), .Q (new_AGEMA_signal_7195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4678 ( .C (clk), .D (new_AGEMA_signal_7198), .Q (new_AGEMA_signal_7199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4682 ( .C (clk), .D (new_AGEMA_signal_7202), .Q (new_AGEMA_signal_7203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4686 ( .C (clk), .D (new_AGEMA_signal_7206), .Q (new_AGEMA_signal_7207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4690 ( .C (clk), .D (new_AGEMA_signal_7210), .Q (new_AGEMA_signal_7211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4694 ( .C (clk), .D (new_AGEMA_signal_7214), .Q (new_AGEMA_signal_7215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4698 ( .C (clk), .D (new_AGEMA_signal_7218), .Q (new_AGEMA_signal_7219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4702 ( .C (clk), .D (new_AGEMA_signal_7222), .Q (new_AGEMA_signal_7223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4706 ( .C (clk), .D (new_AGEMA_signal_7226), .Q (new_AGEMA_signal_7227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4710 ( .C (clk), .D (new_AGEMA_signal_7230), .Q (new_AGEMA_signal_7231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4714 ( .C (clk), .D (new_AGEMA_signal_7234), .Q (new_AGEMA_signal_7235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4718 ( .C (clk), .D (new_AGEMA_signal_7238), .Q (new_AGEMA_signal_7239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4722 ( .C (clk), .D (new_AGEMA_signal_7242), .Q (new_AGEMA_signal_7243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4726 ( .C (clk), .D (new_AGEMA_signal_7246), .Q (new_AGEMA_signal_7247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4730 ( .C (clk), .D (new_AGEMA_signal_7250), .Q (new_AGEMA_signal_7251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4734 ( .C (clk), .D (new_AGEMA_signal_7254), .Q (new_AGEMA_signal_7255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4738 ( .C (clk), .D (new_AGEMA_signal_7258), .Q (new_AGEMA_signal_7259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4742 ( .C (clk), .D (new_AGEMA_signal_7262), .Q (new_AGEMA_signal_7263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4746 ( .C (clk), .D (new_AGEMA_signal_7266), .Q (new_AGEMA_signal_7267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4750 ( .C (clk), .D (new_AGEMA_signal_7270), .Q (new_AGEMA_signal_7271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4754 ( .C (clk), .D (new_AGEMA_signal_7274), .Q (new_AGEMA_signal_7275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4758 ( .C (clk), .D (new_AGEMA_signal_7278), .Q (new_AGEMA_signal_7279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4762 ( .C (clk), .D (new_AGEMA_signal_7282), .Q (new_AGEMA_signal_7283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4766 ( .C (clk), .D (new_AGEMA_signal_7286), .Q (new_AGEMA_signal_7287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4770 ( .C (clk), .D (new_AGEMA_signal_7290), .Q (new_AGEMA_signal_7291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4774 ( .C (clk), .D (new_AGEMA_signal_7294), .Q (new_AGEMA_signal_7295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4778 ( .C (clk), .D (new_AGEMA_signal_7298), .Q (new_AGEMA_signal_7299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4782 ( .C (clk), .D (new_AGEMA_signal_7302), .Q (new_AGEMA_signal_7303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4786 ( .C (clk), .D (new_AGEMA_signal_7306), .Q (new_AGEMA_signal_7307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4790 ( .C (clk), .D (new_AGEMA_signal_7310), .Q (new_AGEMA_signal_7311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4794 ( .C (clk), .D (new_AGEMA_signal_7314), .Q (new_AGEMA_signal_7315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4798 ( .C (clk), .D (new_AGEMA_signal_7318), .Q (new_AGEMA_signal_7319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4802 ( .C (clk), .D (new_AGEMA_signal_7322), .Q (new_AGEMA_signal_7323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4806 ( .C (clk), .D (new_AGEMA_signal_7326), .Q (new_AGEMA_signal_7327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4810 ( .C (clk), .D (new_AGEMA_signal_7330), .Q (new_AGEMA_signal_7331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4814 ( .C (clk), .D (new_AGEMA_signal_7334), .Q (new_AGEMA_signal_7335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4818 ( .C (clk), .D (new_AGEMA_signal_7338), .Q (new_AGEMA_signal_7339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4822 ( .C (clk), .D (new_AGEMA_signal_7342), .Q (new_AGEMA_signal_7343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4826 ( .C (clk), .D (new_AGEMA_signal_7346), .Q (new_AGEMA_signal_7347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4830 ( .C (clk), .D (new_AGEMA_signal_7350), .Q (new_AGEMA_signal_7351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4834 ( .C (clk), .D (new_AGEMA_signal_7354), .Q (new_AGEMA_signal_7355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4838 ( .C (clk), .D (new_AGEMA_signal_7358), .Q (new_AGEMA_signal_7359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4842 ( .C (clk), .D (new_AGEMA_signal_7362), .Q (new_AGEMA_signal_7363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4846 ( .C (clk), .D (new_AGEMA_signal_7366), .Q (new_AGEMA_signal_7367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4850 ( .C (clk), .D (new_AGEMA_signal_7370), .Q (new_AGEMA_signal_7371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4854 ( .C (clk), .D (new_AGEMA_signal_7374), .Q (new_AGEMA_signal_7375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4858 ( .C (clk), .D (new_AGEMA_signal_7378), .Q (new_AGEMA_signal_7379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4862 ( .C (clk), .D (new_AGEMA_signal_7382), .Q (new_AGEMA_signal_7383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4866 ( .C (clk), .D (new_AGEMA_signal_7386), .Q (new_AGEMA_signal_7387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4870 ( .C (clk), .D (new_AGEMA_signal_7390), .Q (new_AGEMA_signal_7391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4874 ( .C (clk), .D (new_AGEMA_signal_7394), .Q (new_AGEMA_signal_7395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4878 ( .C (clk), .D (new_AGEMA_signal_7398), .Q (new_AGEMA_signal_7399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4882 ( .C (clk), .D (new_AGEMA_signal_7402), .Q (new_AGEMA_signal_7403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4886 ( .C (clk), .D (new_AGEMA_signal_7406), .Q (new_AGEMA_signal_7407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4890 ( .C (clk), .D (new_AGEMA_signal_7410), .Q (new_AGEMA_signal_7411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4894 ( .C (clk), .D (new_AGEMA_signal_7414), .Q (new_AGEMA_signal_7415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4898 ( .C (clk), .D (new_AGEMA_signal_7418), .Q (new_AGEMA_signal_7419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4902 ( .C (clk), .D (new_AGEMA_signal_7422), .Q (new_AGEMA_signal_7423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4906 ( .C (clk), .D (new_AGEMA_signal_7426), .Q (new_AGEMA_signal_7427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4910 ( .C (clk), .D (new_AGEMA_signal_7430), .Q (new_AGEMA_signal_7431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4914 ( .C (clk), .D (new_AGEMA_signal_7434), .Q (new_AGEMA_signal_7435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4918 ( .C (clk), .D (new_AGEMA_signal_7438), .Q (new_AGEMA_signal_7439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4922 ( .C (clk), .D (new_AGEMA_signal_7442), .Q (new_AGEMA_signal_7443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4926 ( .C (clk), .D (new_AGEMA_signal_7446), .Q (new_AGEMA_signal_7447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4930 ( .C (clk), .D (new_AGEMA_signal_7450), .Q (new_AGEMA_signal_7451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4934 ( .C (clk), .D (new_AGEMA_signal_7454), .Q (new_AGEMA_signal_7455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4938 ( .C (clk), .D (new_AGEMA_signal_7458), .Q (new_AGEMA_signal_7459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4942 ( .C (clk), .D (new_AGEMA_signal_7462), .Q (new_AGEMA_signal_7463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4946 ( .C (clk), .D (new_AGEMA_signal_7466), .Q (new_AGEMA_signal_7467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4950 ( .C (clk), .D (new_AGEMA_signal_7470), .Q (new_AGEMA_signal_7471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4954 ( .C (clk), .D (new_AGEMA_signal_7474), .Q (new_AGEMA_signal_7475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4958 ( .C (clk), .D (new_AGEMA_signal_7478), .Q (new_AGEMA_signal_7479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4962 ( .C (clk), .D (new_AGEMA_signal_7482), .Q (new_AGEMA_signal_7483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4966 ( .C (clk), .D (new_AGEMA_signal_7486), .Q (new_AGEMA_signal_7487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4970 ( .C (clk), .D (new_AGEMA_signal_7490), .Q (new_AGEMA_signal_7491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4974 ( .C (clk), .D (new_AGEMA_signal_7494), .Q (new_AGEMA_signal_7495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4978 ( .C (clk), .D (new_AGEMA_signal_7498), .Q (new_AGEMA_signal_7499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4982 ( .C (clk), .D (new_AGEMA_signal_7502), .Q (new_AGEMA_signal_7503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4986 ( .C (clk), .D (new_AGEMA_signal_7506), .Q (new_AGEMA_signal_7507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4990 ( .C (clk), .D (new_AGEMA_signal_7510), .Q (new_AGEMA_signal_7511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4994 ( .C (clk), .D (new_AGEMA_signal_7514), .Q (new_AGEMA_signal_7515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4998 ( .C (clk), .D (new_AGEMA_signal_7518), .Q (new_AGEMA_signal_7519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5002 ( .C (clk), .D (new_AGEMA_signal_7522), .Q (new_AGEMA_signal_7523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5006 ( .C (clk), .D (new_AGEMA_signal_7526), .Q (new_AGEMA_signal_7527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5010 ( .C (clk), .D (new_AGEMA_signal_7530), .Q (new_AGEMA_signal_7531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5014 ( .C (clk), .D (new_AGEMA_signal_7534), .Q (new_AGEMA_signal_7535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5018 ( .C (clk), .D (new_AGEMA_signal_7538), .Q (new_AGEMA_signal_7539) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5022 ( .C (clk), .D (new_AGEMA_signal_7542), .Q (new_AGEMA_signal_7543) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5026 ( .C (clk), .D (new_AGEMA_signal_7546), .Q (new_AGEMA_signal_7547) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5030 ( .C (clk), .D (new_AGEMA_signal_7550), .Q (new_AGEMA_signal_7551) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5034 ( .C (clk), .D (new_AGEMA_signal_7554), .Q (new_AGEMA_signal_7555) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5038 ( .C (clk), .D (new_AGEMA_signal_7558), .Q (new_AGEMA_signal_7559) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5042 ( .C (clk), .D (new_AGEMA_signal_7562), .Q (new_AGEMA_signal_7563) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5046 ( .C (clk), .D (new_AGEMA_signal_7566), .Q (new_AGEMA_signal_7567) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5050 ( .C (clk), .D (new_AGEMA_signal_7570), .Q (new_AGEMA_signal_7571) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5054 ( .C (clk), .D (new_AGEMA_signal_7574), .Q (new_AGEMA_signal_7575) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5058 ( .C (clk), .D (new_AGEMA_signal_7578), .Q (new_AGEMA_signal_7579) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5062 ( .C (clk), .D (new_AGEMA_signal_7582), .Q (new_AGEMA_signal_7583) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5066 ( .C (clk), .D (new_AGEMA_signal_7586), .Q (new_AGEMA_signal_7587) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5070 ( .C (clk), .D (new_AGEMA_signal_7590), .Q (new_AGEMA_signal_7591) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5074 ( .C (clk), .D (new_AGEMA_signal_7594), .Q (new_AGEMA_signal_7595) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5078 ( .C (clk), .D (new_AGEMA_signal_7598), .Q (new_AGEMA_signal_7599) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5082 ( .C (clk), .D (new_AGEMA_signal_7602), .Q (new_AGEMA_signal_7603) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5086 ( .C (clk), .D (new_AGEMA_signal_7606), .Q (new_AGEMA_signal_7607) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5090 ( .C (clk), .D (new_AGEMA_signal_7610), .Q (new_AGEMA_signal_7611) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5094 ( .C (clk), .D (new_AGEMA_signal_7614), .Q (new_AGEMA_signal_7615) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5098 ( .C (clk), .D (new_AGEMA_signal_7618), .Q (new_AGEMA_signal_7619) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5102 ( .C (clk), .D (new_AGEMA_signal_7622), .Q (new_AGEMA_signal_7623) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5106 ( .C (clk), .D (new_AGEMA_signal_7626), .Q (new_AGEMA_signal_7627) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5110 ( .C (clk), .D (new_AGEMA_signal_7630), .Q (new_AGEMA_signal_7631) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5114 ( .C (clk), .D (new_AGEMA_signal_7634), .Q (new_AGEMA_signal_7635) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5118 ( .C (clk), .D (new_AGEMA_signal_7638), .Q (new_AGEMA_signal_7639) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5122 ( .C (clk), .D (new_AGEMA_signal_7642), .Q (new_AGEMA_signal_7643) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5126 ( .C (clk), .D (new_AGEMA_signal_7646), .Q (new_AGEMA_signal_7647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5130 ( .C (clk), .D (new_AGEMA_signal_7650), .Q (new_AGEMA_signal_7651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5134 ( .C (clk), .D (new_AGEMA_signal_7654), .Q (new_AGEMA_signal_7655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5138 ( .C (clk), .D (new_AGEMA_signal_7658), .Q (new_AGEMA_signal_7659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5142 ( .C (clk), .D (new_AGEMA_signal_7662), .Q (new_AGEMA_signal_7663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5146 ( .C (clk), .D (new_AGEMA_signal_7666), .Q (new_AGEMA_signal_7667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5150 ( .C (clk), .D (new_AGEMA_signal_7670), .Q (new_AGEMA_signal_7671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5154 ( .C (clk), .D (new_AGEMA_signal_7674), .Q (new_AGEMA_signal_7675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5158 ( .C (clk), .D (new_AGEMA_signal_7678), .Q (new_AGEMA_signal_7679) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5162 ( .C (clk), .D (new_AGEMA_signal_7682), .Q (new_AGEMA_signal_7683) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5166 ( .C (clk), .D (new_AGEMA_signal_7686), .Q (new_AGEMA_signal_7687) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5170 ( .C (clk), .D (new_AGEMA_signal_7690), .Q (new_AGEMA_signal_7691) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5174 ( .C (clk), .D (new_AGEMA_signal_7694), .Q (new_AGEMA_signal_7695) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5178 ( .C (clk), .D (new_AGEMA_signal_7698), .Q (new_AGEMA_signal_7699) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5182 ( .C (clk), .D (new_AGEMA_signal_7702), .Q (new_AGEMA_signal_7703) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5186 ( .C (clk), .D (new_AGEMA_signal_7706), .Q (new_AGEMA_signal_7707) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5190 ( .C (clk), .D (new_AGEMA_signal_7710), .Q (new_AGEMA_signal_7711) ) ;
    buf_clk new_AGEMA_reg_buffer_5194 ( .C (clk), .D (new_AGEMA_signal_7714), .Q (new_AGEMA_signal_7715) ) ;
    buf_clk new_AGEMA_reg_buffer_5198 ( .C (clk), .D (new_AGEMA_signal_7718), .Q (new_AGEMA_signal_7719) ) ;
    buf_clk new_AGEMA_reg_buffer_5202 ( .C (clk), .D (new_AGEMA_signal_7722), .Q (new_AGEMA_signal_7723) ) ;
    buf_clk new_AGEMA_reg_buffer_5206 ( .C (clk), .D (new_AGEMA_signal_7726), .Q (new_AGEMA_signal_7727) ) ;
    buf_clk new_AGEMA_reg_buffer_5210 ( .C (clk), .D (new_AGEMA_signal_7730), .Q (new_AGEMA_signal_7731) ) ;
    buf_clk new_AGEMA_reg_buffer_5214 ( .C (clk), .D (new_AGEMA_signal_7734), .Q (new_AGEMA_signal_7735) ) ;
    buf_clk new_AGEMA_reg_buffer_5218 ( .C (clk), .D (new_AGEMA_signal_7738), .Q (new_AGEMA_signal_7739) ) ;
    buf_clk new_AGEMA_reg_buffer_5222 ( .C (clk), .D (new_AGEMA_signal_7742), .Q (new_AGEMA_signal_7743) ) ;
    buf_clk new_AGEMA_reg_buffer_5226 ( .C (clk), .D (new_AGEMA_signal_7746), .Q (new_AGEMA_signal_7747) ) ;
    buf_clk new_AGEMA_reg_buffer_5230 ( .C (clk), .D (new_AGEMA_signal_7750), .Q (new_AGEMA_signal_7751) ) ;
    buf_clk new_AGEMA_reg_buffer_5234 ( .C (clk), .D (new_AGEMA_signal_7754), .Q (new_AGEMA_signal_7755) ) ;
    buf_clk new_AGEMA_reg_buffer_5238 ( .C (clk), .D (new_AGEMA_signal_7758), .Q (new_AGEMA_signal_7759) ) ;
    buf_clk new_AGEMA_reg_buffer_5242 ( .C (clk), .D (new_AGEMA_signal_7762), .Q (new_AGEMA_signal_7763) ) ;
    buf_clk new_AGEMA_reg_buffer_5246 ( .C (clk), .D (new_AGEMA_signal_7766), .Q (new_AGEMA_signal_7767) ) ;
    buf_clk new_AGEMA_reg_buffer_5250 ( .C (clk), .D (new_AGEMA_signal_7770), .Q (new_AGEMA_signal_7771) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5254 ( .C (clk), .D (new_AGEMA_signal_7774), .Q (new_AGEMA_signal_7775) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5258 ( .C (clk), .D (new_AGEMA_signal_7778), .Q (new_AGEMA_signal_7779) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5262 ( .C (clk), .D (new_AGEMA_signal_7782), .Q (new_AGEMA_signal_7783) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5266 ( .C (clk), .D (new_AGEMA_signal_7786), .Q (new_AGEMA_signal_7787) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5270 ( .C (clk), .D (new_AGEMA_signal_7790), .Q (new_AGEMA_signal_7791) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5274 ( .C (clk), .D (new_AGEMA_signal_7794), .Q (new_AGEMA_signal_7795) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5278 ( .C (clk), .D (new_AGEMA_signal_7798), .Q (new_AGEMA_signal_7799) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5282 ( .C (clk), .D (new_AGEMA_signal_7802), .Q (new_AGEMA_signal_7803) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5286 ( .C (clk), .D (new_AGEMA_signal_7806), .Q (new_AGEMA_signal_7807) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5290 ( .C (clk), .D (new_AGEMA_signal_7810), .Q (new_AGEMA_signal_7811) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5294 ( .C (clk), .D (new_AGEMA_signal_7814), .Q (new_AGEMA_signal_7815) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5298 ( .C (clk), .D (new_AGEMA_signal_7818), .Q (new_AGEMA_signal_7819) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5302 ( .C (clk), .D (new_AGEMA_signal_7822), .Q (new_AGEMA_signal_7823) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5306 ( .C (clk), .D (new_AGEMA_signal_7826), .Q (new_AGEMA_signal_7827) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5310 ( .C (clk), .D (new_AGEMA_signal_7830), .Q (new_AGEMA_signal_7831) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5314 ( .C (clk), .D (new_AGEMA_signal_7834), .Q (new_AGEMA_signal_7835) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5318 ( .C (clk), .D (new_AGEMA_signal_7838), .Q (new_AGEMA_signal_7839) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5322 ( .C (clk), .D (new_AGEMA_signal_7842), .Q (new_AGEMA_signal_7843) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5326 ( .C (clk), .D (new_AGEMA_signal_7846), .Q (new_AGEMA_signal_7847) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5330 ( .C (clk), .D (new_AGEMA_signal_7850), .Q (new_AGEMA_signal_7851) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5334 ( .C (clk), .D (new_AGEMA_signal_7854), .Q (new_AGEMA_signal_7855) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5338 ( .C (clk), .D (new_AGEMA_signal_7858), .Q (new_AGEMA_signal_7859) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5342 ( .C (clk), .D (new_AGEMA_signal_7862), .Q (new_AGEMA_signal_7863) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5346 ( .C (clk), .D (new_AGEMA_signal_7866), .Q (new_AGEMA_signal_7867) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5350 ( .C (clk), .D (new_AGEMA_signal_7870), .Q (new_AGEMA_signal_7871) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5354 ( .C (clk), .D (new_AGEMA_signal_7874), .Q (new_AGEMA_signal_7875) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5358 ( .C (clk), .D (new_AGEMA_signal_7878), .Q (new_AGEMA_signal_7879) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5362 ( .C (clk), .D (new_AGEMA_signal_7882), .Q (new_AGEMA_signal_7883) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5366 ( .C (clk), .D (new_AGEMA_signal_7886), .Q (new_AGEMA_signal_7887) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5370 ( .C (clk), .D (new_AGEMA_signal_7890), .Q (new_AGEMA_signal_7891) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5374 ( .C (clk), .D (new_AGEMA_signal_7894), .Q (new_AGEMA_signal_7895) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5378 ( .C (clk), .D (new_AGEMA_signal_7898), .Q (new_AGEMA_signal_7899) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5382 ( .C (clk), .D (new_AGEMA_signal_7902), .Q (new_AGEMA_signal_7903) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5386 ( .C (clk), .D (new_AGEMA_signal_7906), .Q (new_AGEMA_signal_7907) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5390 ( .C (clk), .D (new_AGEMA_signal_7910), .Q (new_AGEMA_signal_7911) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5394 ( .C (clk), .D (new_AGEMA_signal_7914), .Q (new_AGEMA_signal_7915) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5398 ( .C (clk), .D (new_AGEMA_signal_7918), .Q (new_AGEMA_signal_7919) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5402 ( .C (clk), .D (new_AGEMA_signal_7922), .Q (new_AGEMA_signal_7923) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5406 ( .C (clk), .D (new_AGEMA_signal_7926), .Q (new_AGEMA_signal_7927) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5410 ( .C (clk), .D (new_AGEMA_signal_7930), .Q (new_AGEMA_signal_7931) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5414 ( .C (clk), .D (new_AGEMA_signal_7934), .Q (new_AGEMA_signal_7935) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5418 ( .C (clk), .D (new_AGEMA_signal_7938), .Q (new_AGEMA_signal_7939) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5422 ( .C (clk), .D (new_AGEMA_signal_7942), .Q (new_AGEMA_signal_7943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5426 ( .C (clk), .D (new_AGEMA_signal_7946), .Q (new_AGEMA_signal_7947) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5430 ( .C (clk), .D (new_AGEMA_signal_7950), .Q (new_AGEMA_signal_7951) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5434 ( .C (clk), .D (new_AGEMA_signal_7954), .Q (new_AGEMA_signal_7955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5438 ( .C (clk), .D (new_AGEMA_signal_7958), .Q (new_AGEMA_signal_7959) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5442 ( .C (clk), .D (new_AGEMA_signal_7962), .Q (new_AGEMA_signal_7963) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5446 ( .C (clk), .D (new_AGEMA_signal_7966), .Q (new_AGEMA_signal_7967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5450 ( .C (clk), .D (new_AGEMA_signal_7970), .Q (new_AGEMA_signal_7971) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5454 ( .C (clk), .D (new_AGEMA_signal_7974), .Q (new_AGEMA_signal_7975) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5458 ( .C (clk), .D (new_AGEMA_signal_7978), .Q (new_AGEMA_signal_7979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5462 ( .C (clk), .D (new_AGEMA_signal_7982), .Q (new_AGEMA_signal_7983) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5466 ( .C (clk), .D (new_AGEMA_signal_7986), .Q (new_AGEMA_signal_7987) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5470 ( .C (clk), .D (new_AGEMA_signal_7990), .Q (new_AGEMA_signal_7991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5474 ( .C (clk), .D (new_AGEMA_signal_7994), .Q (new_AGEMA_signal_7995) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5478 ( .C (clk), .D (new_AGEMA_signal_7998), .Q (new_AGEMA_signal_7999) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5482 ( .C (clk), .D (new_AGEMA_signal_8002), .Q (new_AGEMA_signal_8003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5486 ( .C (clk), .D (new_AGEMA_signal_8006), .Q (new_AGEMA_signal_8007) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5490 ( .C (clk), .D (new_AGEMA_signal_8010), .Q (new_AGEMA_signal_8011) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5494 ( .C (clk), .D (new_AGEMA_signal_8014), .Q (new_AGEMA_signal_8015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5498 ( .C (clk), .D (new_AGEMA_signal_8018), .Q (new_AGEMA_signal_8019) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5502 ( .C (clk), .D (new_AGEMA_signal_8022), .Q (new_AGEMA_signal_8023) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5506 ( .C (clk), .D (new_AGEMA_signal_8026), .Q (new_AGEMA_signal_8027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5510 ( .C (clk), .D (new_AGEMA_signal_8030), .Q (new_AGEMA_signal_8031) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5514 ( .C (clk), .D (new_AGEMA_signal_8034), .Q (new_AGEMA_signal_8035) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5518 ( .C (clk), .D (new_AGEMA_signal_8038), .Q (new_AGEMA_signal_8039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5522 ( .C (clk), .D (new_AGEMA_signal_8042), .Q (new_AGEMA_signal_8043) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5526 ( .C (clk), .D (new_AGEMA_signal_8046), .Q (new_AGEMA_signal_8047) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5530 ( .C (clk), .D (new_AGEMA_signal_8050), .Q (new_AGEMA_signal_8051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5534 ( .C (clk), .D (new_AGEMA_signal_8054), .Q (new_AGEMA_signal_8055) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5538 ( .C (clk), .D (new_AGEMA_signal_8058), .Q (new_AGEMA_signal_8059) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5542 ( .C (clk), .D (new_AGEMA_signal_8062), .Q (new_AGEMA_signal_8063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5546 ( .C (clk), .D (new_AGEMA_signal_8066), .Q (new_AGEMA_signal_8067) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5550 ( .C (clk), .D (new_AGEMA_signal_8070), .Q (new_AGEMA_signal_8071) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5554 ( .C (clk), .D (new_AGEMA_signal_8074), .Q (new_AGEMA_signal_8075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5558 ( .C (clk), .D (new_AGEMA_signal_8078), .Q (new_AGEMA_signal_8079) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5562 ( .C (clk), .D (new_AGEMA_signal_8082), .Q (new_AGEMA_signal_8083) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5566 ( .C (clk), .D (new_AGEMA_signal_8086), .Q (new_AGEMA_signal_8087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5570 ( .C (clk), .D (new_AGEMA_signal_8090), .Q (new_AGEMA_signal_8091) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5574 ( .C (clk), .D (new_AGEMA_signal_8094), .Q (new_AGEMA_signal_8095) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5578 ( .C (clk), .D (new_AGEMA_signal_8098), .Q (new_AGEMA_signal_8099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5582 ( .C (clk), .D (new_AGEMA_signal_8102), .Q (new_AGEMA_signal_8103) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5586 ( .C (clk), .D (new_AGEMA_signal_8106), .Q (new_AGEMA_signal_8107) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5590 ( .C (clk), .D (new_AGEMA_signal_8110), .Q (new_AGEMA_signal_8111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5594 ( .C (clk), .D (new_AGEMA_signal_8114), .Q (new_AGEMA_signal_8115) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5598 ( .C (clk), .D (new_AGEMA_signal_8118), .Q (new_AGEMA_signal_8119) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5602 ( .C (clk), .D (new_AGEMA_signal_8122), .Q (new_AGEMA_signal_8123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5606 ( .C (clk), .D (new_AGEMA_signal_8126), .Q (new_AGEMA_signal_8127) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5610 ( .C (clk), .D (new_AGEMA_signal_8130), .Q (new_AGEMA_signal_8131) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5614 ( .C (clk), .D (new_AGEMA_signal_8134), .Q (new_AGEMA_signal_8135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5618 ( .C (clk), .D (new_AGEMA_signal_8138), .Q (new_AGEMA_signal_8139) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5622 ( .C (clk), .D (new_AGEMA_signal_8142), .Q (new_AGEMA_signal_8143) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5626 ( .C (clk), .D (new_AGEMA_signal_8146), .Q (new_AGEMA_signal_8147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5630 ( .C (clk), .D (new_AGEMA_signal_8150), .Q (new_AGEMA_signal_8151) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5634 ( .C (clk), .D (new_AGEMA_signal_8154), .Q (new_AGEMA_signal_8155) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5638 ( .C (clk), .D (new_AGEMA_signal_8158), .Q (new_AGEMA_signal_8159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5642 ( .C (clk), .D (new_AGEMA_signal_8162), .Q (new_AGEMA_signal_8163) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5646 ( .C (clk), .D (new_AGEMA_signal_8166), .Q (new_AGEMA_signal_8167) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5650 ( .C (clk), .D (new_AGEMA_signal_8170), .Q (new_AGEMA_signal_8171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5654 ( .C (clk), .D (new_AGEMA_signal_8174), .Q (new_AGEMA_signal_8175) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5658 ( .C (clk), .D (new_AGEMA_signal_8178), .Q (new_AGEMA_signal_8179) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5662 ( .C (clk), .D (new_AGEMA_signal_8182), .Q (new_AGEMA_signal_8183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5666 ( .C (clk), .D (new_AGEMA_signal_8186), .Q (new_AGEMA_signal_8187) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5670 ( .C (clk), .D (new_AGEMA_signal_8190), .Q (new_AGEMA_signal_8191) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5674 ( .C (clk), .D (new_AGEMA_signal_8194), .Q (new_AGEMA_signal_8195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5678 ( .C (clk), .D (new_AGEMA_signal_8198), .Q (new_AGEMA_signal_8199) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5682 ( .C (clk), .D (new_AGEMA_signal_8202), .Q (new_AGEMA_signal_8203) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5686 ( .C (clk), .D (new_AGEMA_signal_8206), .Q (new_AGEMA_signal_8207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5690 ( .C (clk), .D (new_AGEMA_signal_8210), .Q (new_AGEMA_signal_8211) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5694 ( .C (clk), .D (new_AGEMA_signal_8214), .Q (new_AGEMA_signal_8215) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5698 ( .C (clk), .D (new_AGEMA_signal_8218), .Q (new_AGEMA_signal_8219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5702 ( .C (clk), .D (new_AGEMA_signal_8222), .Q (new_AGEMA_signal_8223) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5706 ( .C (clk), .D (new_AGEMA_signal_8226), .Q (new_AGEMA_signal_8227) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5710 ( .C (clk), .D (new_AGEMA_signal_8230), .Q (new_AGEMA_signal_8231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5714 ( .C (clk), .D (new_AGEMA_signal_8234), .Q (new_AGEMA_signal_8235) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5718 ( .C (clk), .D (new_AGEMA_signal_8238), .Q (new_AGEMA_signal_8239) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5722 ( .C (clk), .D (new_AGEMA_signal_8242), .Q (new_AGEMA_signal_8243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5726 ( .C (clk), .D (new_AGEMA_signal_8246), .Q (new_AGEMA_signal_8247) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5730 ( .C (clk), .D (new_AGEMA_signal_8250), .Q (new_AGEMA_signal_8251) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5734 ( .C (clk), .D (new_AGEMA_signal_8254), .Q (new_AGEMA_signal_8255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5738 ( .C (clk), .D (new_AGEMA_signal_8258), .Q (new_AGEMA_signal_8259) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5742 ( .C (clk), .D (new_AGEMA_signal_8262), .Q (new_AGEMA_signal_8263) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5746 ( .C (clk), .D (new_AGEMA_signal_8266), .Q (new_AGEMA_signal_8267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5750 ( .C (clk), .D (new_AGEMA_signal_8270), .Q (new_AGEMA_signal_8271) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5754 ( .C (clk), .D (new_AGEMA_signal_8274), .Q (new_AGEMA_signal_8275) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5758 ( .C (clk), .D (new_AGEMA_signal_8278), .Q (new_AGEMA_signal_8279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5762 ( .C (clk), .D (new_AGEMA_signal_8282), .Q (new_AGEMA_signal_8283) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5766 ( .C (clk), .D (new_AGEMA_signal_8286), .Q (new_AGEMA_signal_8287) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5770 ( .C (clk), .D (new_AGEMA_signal_8290), .Q (new_AGEMA_signal_8291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5774 ( .C (clk), .D (new_AGEMA_signal_8294), .Q (new_AGEMA_signal_8295) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5778 ( .C (clk), .D (new_AGEMA_signal_8298), .Q (new_AGEMA_signal_8299) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5782 ( .C (clk), .D (new_AGEMA_signal_8302), .Q (new_AGEMA_signal_8303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5786 ( .C (clk), .D (new_AGEMA_signal_8306), .Q (new_AGEMA_signal_8307) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5790 ( .C (clk), .D (new_AGEMA_signal_8310), .Q (new_AGEMA_signal_8311) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5794 ( .C (clk), .D (new_AGEMA_signal_8314), .Q (new_AGEMA_signal_8315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5798 ( .C (clk), .D (new_AGEMA_signal_8318), .Q (new_AGEMA_signal_8319) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5802 ( .C (clk), .D (new_AGEMA_signal_8322), .Q (new_AGEMA_signal_8323) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5806 ( .C (clk), .D (new_AGEMA_signal_8326), .Q (new_AGEMA_signal_8327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5810 ( .C (clk), .D (new_AGEMA_signal_8330), .Q (new_AGEMA_signal_8331) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5814 ( .C (clk), .D (new_AGEMA_signal_8334), .Q (new_AGEMA_signal_8335) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5818 ( .C (clk), .D (new_AGEMA_signal_8338), .Q (new_AGEMA_signal_8339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5822 ( .C (clk), .D (new_AGEMA_signal_8342), .Q (new_AGEMA_signal_8343) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5826 ( .C (clk), .D (new_AGEMA_signal_8346), .Q (new_AGEMA_signal_8347) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5830 ( .C (clk), .D (new_AGEMA_signal_8350), .Q (new_AGEMA_signal_8351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5834 ( .C (clk), .D (new_AGEMA_signal_8354), .Q (new_AGEMA_signal_8355) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5838 ( .C (clk), .D (new_AGEMA_signal_8358), .Q (new_AGEMA_signal_8359) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5842 ( .C (clk), .D (new_AGEMA_signal_8362), .Q (new_AGEMA_signal_8363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5846 ( .C (clk), .D (new_AGEMA_signal_8366), .Q (new_AGEMA_signal_8367) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5850 ( .C (clk), .D (new_AGEMA_signal_8370), .Q (new_AGEMA_signal_8371) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5854 ( .C (clk), .D (new_AGEMA_signal_8374), .Q (new_AGEMA_signal_8375) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5858 ( .C (clk), .D (new_AGEMA_signal_8378), .Q (new_AGEMA_signal_8379) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5862 ( .C (clk), .D (new_AGEMA_signal_8382), .Q (new_AGEMA_signal_8383) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5866 ( .C (clk), .D (new_AGEMA_signal_8386), .Q (new_AGEMA_signal_8387) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5870 ( .C (clk), .D (new_AGEMA_signal_8390), .Q (new_AGEMA_signal_8391) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5874 ( .C (clk), .D (new_AGEMA_signal_8394), .Q (new_AGEMA_signal_8395) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5878 ( .C (clk), .D (new_AGEMA_signal_8398), .Q (new_AGEMA_signal_8399) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5882 ( .C (clk), .D (new_AGEMA_signal_8402), .Q (new_AGEMA_signal_8403) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5886 ( .C (clk), .D (new_AGEMA_signal_8406), .Q (new_AGEMA_signal_8407) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5890 ( .C (clk), .D (new_AGEMA_signal_8410), .Q (new_AGEMA_signal_8411) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5894 ( .C (clk), .D (new_AGEMA_signal_8414), .Q (new_AGEMA_signal_8415) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5898 ( .C (clk), .D (new_AGEMA_signal_8418), .Q (new_AGEMA_signal_8419) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5902 ( .C (clk), .D (new_AGEMA_signal_8422), .Q (new_AGEMA_signal_8423) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5906 ( .C (clk), .D (new_AGEMA_signal_8426), .Q (new_AGEMA_signal_8427) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5910 ( .C (clk), .D (new_AGEMA_signal_8430), .Q (new_AGEMA_signal_8431) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5914 ( .C (clk), .D (new_AGEMA_signal_8434), .Q (new_AGEMA_signal_8435) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5918 ( .C (clk), .D (new_AGEMA_signal_8438), .Q (new_AGEMA_signal_8439) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5922 ( .C (clk), .D (new_AGEMA_signal_8442), .Q (new_AGEMA_signal_8443) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5926 ( .C (clk), .D (new_AGEMA_signal_8446), .Q (new_AGEMA_signal_8447) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5930 ( .C (clk), .D (new_AGEMA_signal_8450), .Q (new_AGEMA_signal_8451) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5934 ( .C (clk), .D (new_AGEMA_signal_8454), .Q (new_AGEMA_signal_8455) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5938 ( .C (clk), .D (new_AGEMA_signal_8458), .Q (new_AGEMA_signal_8459) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5942 ( .C (clk), .D (new_AGEMA_signal_8462), .Q (new_AGEMA_signal_8463) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5946 ( .C (clk), .D (new_AGEMA_signal_8466), .Q (new_AGEMA_signal_8467) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5950 ( .C (clk), .D (new_AGEMA_signal_8470), .Q (new_AGEMA_signal_8471) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5954 ( .C (clk), .D (new_AGEMA_signal_8474), .Q (new_AGEMA_signal_8475) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5958 ( .C (clk), .D (new_AGEMA_signal_8478), .Q (new_AGEMA_signal_8479) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5962 ( .C (clk), .D (new_AGEMA_signal_8482), .Q (new_AGEMA_signal_8483) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5966 ( .C (clk), .D (new_AGEMA_signal_8486), .Q (new_AGEMA_signal_8487) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5970 ( .C (clk), .D (new_AGEMA_signal_8490), .Q (new_AGEMA_signal_8491) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5974 ( .C (clk), .D (new_AGEMA_signal_8494), .Q (new_AGEMA_signal_8495) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5978 ( .C (clk), .D (new_AGEMA_signal_8498), .Q (new_AGEMA_signal_8499) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5982 ( .C (clk), .D (new_AGEMA_signal_8502), .Q (new_AGEMA_signal_8503) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5986 ( .C (clk), .D (new_AGEMA_signal_8506), .Q (new_AGEMA_signal_8507) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5990 ( .C (clk), .D (new_AGEMA_signal_8510), .Q (new_AGEMA_signal_8511) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5994 ( .C (clk), .D (new_AGEMA_signal_8514), .Q (new_AGEMA_signal_8515) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5998 ( .C (clk), .D (new_AGEMA_signal_8518), .Q (new_AGEMA_signal_8519) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6002 ( .C (clk), .D (new_AGEMA_signal_8522), .Q (new_AGEMA_signal_8523) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6006 ( .C (clk), .D (new_AGEMA_signal_8526), .Q (new_AGEMA_signal_8527) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6010 ( .C (clk), .D (new_AGEMA_signal_8530), .Q (new_AGEMA_signal_8531) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6014 ( .C (clk), .D (new_AGEMA_signal_8534), .Q (new_AGEMA_signal_8535) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6018 ( .C (clk), .D (new_AGEMA_signal_8538), .Q (new_AGEMA_signal_8539) ) ;
    buf_clk new_AGEMA_reg_buffer_6022 ( .C (clk), .D (new_AGEMA_signal_8542), .Q (new_AGEMA_signal_8543) ) ;
    buf_clk new_AGEMA_reg_buffer_6026 ( .C (clk), .D (new_AGEMA_signal_8546), .Q (new_AGEMA_signal_8547) ) ;
    buf_clk new_AGEMA_reg_buffer_6030 ( .C (clk), .D (new_AGEMA_signal_8550), .Q (new_AGEMA_signal_8551) ) ;
    buf_clk new_AGEMA_reg_buffer_6034 ( .C (clk), .D (new_AGEMA_signal_8554), .Q (new_AGEMA_signal_8555) ) ;
    buf_clk new_AGEMA_reg_buffer_6038 ( .C (clk), .D (new_AGEMA_signal_8558), .Q (new_AGEMA_signal_8559) ) ;
    buf_clk new_AGEMA_reg_buffer_6042 ( .C (clk), .D (new_AGEMA_signal_8562), .Q (new_AGEMA_signal_8563) ) ;
    buf_clk new_AGEMA_reg_buffer_6046 ( .C (clk), .D (new_AGEMA_signal_8566), .Q (new_AGEMA_signal_8567) ) ;

    /* cells in depth 3 */
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_3256, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_4619, new_AGEMA_signal_4618}), .clk (clk), .r ({Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_3274, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_3255, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_4621, new_AGEMA_signal_4620}), .clk (clk), .r ({Fresh[99], Fresh[98]}), .c ({new_AGEMA_signal_3275, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_4619, new_AGEMA_signal_4618}), .b ({new_AGEMA_signal_3257, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_3276, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_4621, new_AGEMA_signal_4620}), .b ({new_AGEMA_signal_3241, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_3277, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_4647, new_AGEMA_signal_4646}), .b ({new_AGEMA_signal_3274, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_3276, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_4649, new_AGEMA_signal_4648}), .c ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_4651, new_AGEMA_signal_4650}), .b ({new_AGEMA_signal_3275, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_3277, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652}), .c ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_3312, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_3313, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_3358, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_3261, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_4627, new_AGEMA_signal_4626}), .clk (clk), .r ({Fresh[105], Fresh[104]}), .c ({new_AGEMA_signal_3279, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_3260, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_4629, new_AGEMA_signal_4628}), .clk (clk), .r ({Fresh[107], Fresh[106]}), .c ({new_AGEMA_signal_3280, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4626}), .b ({new_AGEMA_signal_3262, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_3281, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_4629, new_AGEMA_signal_4628}), .b ({new_AGEMA_signal_3245, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[111], Fresh[110]}), .c ({new_AGEMA_signal_3282, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_4655, new_AGEMA_signal_4654}), .b ({new_AGEMA_signal_3279, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_3281, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_4657, new_AGEMA_signal_4656}), .c ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_4659, new_AGEMA_signal_4658}), .b ({new_AGEMA_signal_3280, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_3282, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_4661, new_AGEMA_signal_4660}), .c ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_3324, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_3325, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_3370, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_3266, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634}), .clk (clk), .r ({Fresh[113], Fresh[112]}), .c ({new_AGEMA_signal_3284, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_3265, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_4637, new_AGEMA_signal_4636}), .clk (clk), .r ({Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_3285, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_4635, new_AGEMA_signal_4634}), .b ({new_AGEMA_signal_3267, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[117], Fresh[116]}), .c ({new_AGEMA_signal_3286, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_4637, new_AGEMA_signal_4636}), .b ({new_AGEMA_signal_3249, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[119], Fresh[118]}), .c ({new_AGEMA_signal_3287, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_4663, new_AGEMA_signal_4662}), .b ({new_AGEMA_signal_3284, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_3286, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_4665, new_AGEMA_signal_4664}), .c ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_4667, new_AGEMA_signal_4666}), .b ({new_AGEMA_signal_3285, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_3287, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_4669, new_AGEMA_signal_4668}), .c ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_3336, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_3337, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_3382, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_3271, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_4643, new_AGEMA_signal_4642}), .clk (clk), .r ({Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_3289, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_3270, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_4645, new_AGEMA_signal_4644}), .clk (clk), .r ({Fresh[123], Fresh[122]}), .c ({new_AGEMA_signal_3290, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_4643, new_AGEMA_signal_4642}), .b ({new_AGEMA_signal_3272, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[125], Fresh[124]}), .c ({new_AGEMA_signal_3291, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_4645, new_AGEMA_signal_4644}), .b ({new_AGEMA_signal_3253, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_3292, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_4671, new_AGEMA_signal_4670}), .b ({new_AGEMA_signal_3289, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_3291, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_4673, new_AGEMA_signal_4672}), .c ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_4675, new_AGEMA_signal_4674}), .b ({new_AGEMA_signal_3290, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_3292, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_4677, new_AGEMA_signal_4676}), .c ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_3348, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_3349, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_3394, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2125 ( .C (clk), .D (new_AGEMA_signal_4614), .Q (new_AGEMA_signal_4646) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2126 ( .C (clk), .D (new_AGEMA_signal_4615), .Q (new_AGEMA_signal_4647) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2127 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M33), .Q (new_AGEMA_signal_4648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2128 ( .C (clk), .D (new_AGEMA_signal_3258), .Q (new_AGEMA_signal_4649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2129 ( .C (clk), .D (new_AGEMA_signal_4616), .Q (new_AGEMA_signal_4650) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2130 ( .C (clk), .D (new_AGEMA_signal_4617), .Q (new_AGEMA_signal_4651) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2131 ( .C (clk), .D (SubBytesIns_Inst_Sbox_0_M36), .Q (new_AGEMA_signal_4652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2132 ( .C (clk), .D (new_AGEMA_signal_3278), .Q (new_AGEMA_signal_4653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2133 ( .C (clk), .D (new_AGEMA_signal_4622), .Q (new_AGEMA_signal_4654) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2134 ( .C (clk), .D (new_AGEMA_signal_4623), .Q (new_AGEMA_signal_4655) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2135 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M33), .Q (new_AGEMA_signal_4656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2136 ( .C (clk), .D (new_AGEMA_signal_3263), .Q (new_AGEMA_signal_4657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2137 ( .C (clk), .D (new_AGEMA_signal_4624), .Q (new_AGEMA_signal_4658) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2138 ( .C (clk), .D (new_AGEMA_signal_4625), .Q (new_AGEMA_signal_4659) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2139 ( .C (clk), .D (SubBytesIns_Inst_Sbox_1_M36), .Q (new_AGEMA_signal_4660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2140 ( .C (clk), .D (new_AGEMA_signal_3283), .Q (new_AGEMA_signal_4661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2141 ( .C (clk), .D (new_AGEMA_signal_4630), .Q (new_AGEMA_signal_4662) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2142 ( .C (clk), .D (new_AGEMA_signal_4631), .Q (new_AGEMA_signal_4663) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2143 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M33), .Q (new_AGEMA_signal_4664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2144 ( .C (clk), .D (new_AGEMA_signal_3268), .Q (new_AGEMA_signal_4665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2145 ( .C (clk), .D (new_AGEMA_signal_4632), .Q (new_AGEMA_signal_4666) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2146 ( .C (clk), .D (new_AGEMA_signal_4633), .Q (new_AGEMA_signal_4667) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2147 ( .C (clk), .D (SubBytesIns_Inst_Sbox_2_M36), .Q (new_AGEMA_signal_4668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2148 ( .C (clk), .D (new_AGEMA_signal_3288), .Q (new_AGEMA_signal_4669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2149 ( .C (clk), .D (new_AGEMA_signal_4638), .Q (new_AGEMA_signal_4670) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2150 ( .C (clk), .D (new_AGEMA_signal_4639), .Q (new_AGEMA_signal_4671) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2151 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M33), .Q (new_AGEMA_signal_4672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2152 ( .C (clk), .D (new_AGEMA_signal_3273), .Q (new_AGEMA_signal_4673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2153 ( .C (clk), .D (new_AGEMA_signal_4640), .Q (new_AGEMA_signal_4674) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2154 ( .C (clk), .D (new_AGEMA_signal_4641), .Q (new_AGEMA_signal_4675) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2155 ( .C (clk), .D (SubBytesIns_Inst_Sbox_3_M36), .Q (new_AGEMA_signal_4676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2156 ( .C (clk), .D (new_AGEMA_signal_3293), .Q (new_AGEMA_signal_4677) ) ;
    buf_clk new_AGEMA_reg_buffer_2159 ( .C (clk), .D (new_AGEMA_signal_4679), .Q (new_AGEMA_signal_4680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2163 ( .C (clk), .D (new_AGEMA_signal_4683), .Q (new_AGEMA_signal_4684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2167 ( .C (clk), .D (new_AGEMA_signal_4687), .Q (new_AGEMA_signal_4688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2171 ( .C (clk), .D (new_AGEMA_signal_4691), .Q (new_AGEMA_signal_4692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2175 ( .C (clk), .D (new_AGEMA_signal_4695), .Q (new_AGEMA_signal_4696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2179 ( .C (clk), .D (new_AGEMA_signal_4699), .Q (new_AGEMA_signal_4700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2183 ( .C (clk), .D (new_AGEMA_signal_4703), .Q (new_AGEMA_signal_4704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2187 ( .C (clk), .D (new_AGEMA_signal_4707), .Q (new_AGEMA_signal_4708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2191 ( .C (clk), .D (new_AGEMA_signal_4711), .Q (new_AGEMA_signal_4712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2195 ( .C (clk), .D (new_AGEMA_signal_4715), .Q (new_AGEMA_signal_4716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2199 ( .C (clk), .D (new_AGEMA_signal_4719), .Q (new_AGEMA_signal_4720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2203 ( .C (clk), .D (new_AGEMA_signal_4723), .Q (new_AGEMA_signal_4724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2207 ( .C (clk), .D (new_AGEMA_signal_4727), .Q (new_AGEMA_signal_4728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2211 ( .C (clk), .D (new_AGEMA_signal_4731), .Q (new_AGEMA_signal_4732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2215 ( .C (clk), .D (new_AGEMA_signal_4735), .Q (new_AGEMA_signal_4736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2219 ( .C (clk), .D (new_AGEMA_signal_4739), .Q (new_AGEMA_signal_4740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2223 ( .C (clk), .D (new_AGEMA_signal_4743), .Q (new_AGEMA_signal_4744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2227 ( .C (clk), .D (new_AGEMA_signal_4747), .Q (new_AGEMA_signal_4748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2231 ( .C (clk), .D (new_AGEMA_signal_4751), .Q (new_AGEMA_signal_4752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2235 ( .C (clk), .D (new_AGEMA_signal_4755), .Q (new_AGEMA_signal_4756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2239 ( .C (clk), .D (new_AGEMA_signal_4759), .Q (new_AGEMA_signal_4760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2243 ( .C (clk), .D (new_AGEMA_signal_4763), .Q (new_AGEMA_signal_4764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2247 ( .C (clk), .D (new_AGEMA_signal_4767), .Q (new_AGEMA_signal_4768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2251 ( .C (clk), .D (new_AGEMA_signal_4771), .Q (new_AGEMA_signal_4772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2255 ( .C (clk), .D (new_AGEMA_signal_4775), .Q (new_AGEMA_signal_4776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2259 ( .C (clk), .D (new_AGEMA_signal_4779), .Q (new_AGEMA_signal_4780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2263 ( .C (clk), .D (new_AGEMA_signal_4783), .Q (new_AGEMA_signal_4784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2267 ( .C (clk), .D (new_AGEMA_signal_4787), .Q (new_AGEMA_signal_4788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2271 ( .C (clk), .D (new_AGEMA_signal_4791), .Q (new_AGEMA_signal_4792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2275 ( .C (clk), .D (new_AGEMA_signal_4795), .Q (new_AGEMA_signal_4796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2279 ( .C (clk), .D (new_AGEMA_signal_4799), .Q (new_AGEMA_signal_4800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2283 ( .C (clk), .D (new_AGEMA_signal_4803), .Q (new_AGEMA_signal_4804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2287 ( .C (clk), .D (new_AGEMA_signal_4807), .Q (new_AGEMA_signal_4808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2291 ( .C (clk), .D (new_AGEMA_signal_4811), .Q (new_AGEMA_signal_4812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2295 ( .C (clk), .D (new_AGEMA_signal_4815), .Q (new_AGEMA_signal_4816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2299 ( .C (clk), .D (new_AGEMA_signal_4819), .Q (new_AGEMA_signal_4820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2303 ( .C (clk), .D (new_AGEMA_signal_4823), .Q (new_AGEMA_signal_4824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2307 ( .C (clk), .D (new_AGEMA_signal_4827), .Q (new_AGEMA_signal_4828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2311 ( .C (clk), .D (new_AGEMA_signal_4831), .Q (new_AGEMA_signal_4832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2315 ( .C (clk), .D (new_AGEMA_signal_4835), .Q (new_AGEMA_signal_4836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2319 ( .C (clk), .D (new_AGEMA_signal_4839), .Q (new_AGEMA_signal_4840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2323 ( .C (clk), .D (new_AGEMA_signal_4843), .Q (new_AGEMA_signal_4844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2327 ( .C (clk), .D (new_AGEMA_signal_4847), .Q (new_AGEMA_signal_4848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2331 ( .C (clk), .D (new_AGEMA_signal_4851), .Q (new_AGEMA_signal_4852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2335 ( .C (clk), .D (new_AGEMA_signal_4855), .Q (new_AGEMA_signal_4856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2339 ( .C (clk), .D (new_AGEMA_signal_4859), .Q (new_AGEMA_signal_4860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2343 ( .C (clk), .D (new_AGEMA_signal_4863), .Q (new_AGEMA_signal_4864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2347 ( .C (clk), .D (new_AGEMA_signal_4867), .Q (new_AGEMA_signal_4868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2351 ( .C (clk), .D (new_AGEMA_signal_4871), .Q (new_AGEMA_signal_4872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2355 ( .C (clk), .D (new_AGEMA_signal_4875), .Q (new_AGEMA_signal_4876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2359 ( .C (clk), .D (new_AGEMA_signal_4879), .Q (new_AGEMA_signal_4880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2363 ( .C (clk), .D (new_AGEMA_signal_4883), .Q (new_AGEMA_signal_4884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2367 ( .C (clk), .D (new_AGEMA_signal_4887), .Q (new_AGEMA_signal_4888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2371 ( .C (clk), .D (new_AGEMA_signal_4891), .Q (new_AGEMA_signal_4892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2375 ( .C (clk), .D (new_AGEMA_signal_4895), .Q (new_AGEMA_signal_4896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2379 ( .C (clk), .D (new_AGEMA_signal_4899), .Q (new_AGEMA_signal_4900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2383 ( .C (clk), .D (new_AGEMA_signal_4903), .Q (new_AGEMA_signal_4904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2387 ( .C (clk), .D (new_AGEMA_signal_4907), .Q (new_AGEMA_signal_4908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2391 ( .C (clk), .D (new_AGEMA_signal_4911), .Q (new_AGEMA_signal_4912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2395 ( .C (clk), .D (new_AGEMA_signal_4915), .Q (new_AGEMA_signal_4916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2399 ( .C (clk), .D (new_AGEMA_signal_4919), .Q (new_AGEMA_signal_4920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2403 ( .C (clk), .D (new_AGEMA_signal_4923), .Q (new_AGEMA_signal_4924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2407 ( .C (clk), .D (new_AGEMA_signal_4927), .Q (new_AGEMA_signal_4928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2411 ( .C (clk), .D (new_AGEMA_signal_4931), .Q (new_AGEMA_signal_4932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2415 ( .C (clk), .D (new_AGEMA_signal_4935), .Q (new_AGEMA_signal_4936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2419 ( .C (clk), .D (new_AGEMA_signal_4939), .Q (new_AGEMA_signal_4940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2422 ( .C (clk), .D (new_AGEMA_signal_4942), .Q (new_AGEMA_signal_4943) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2425 ( .C (clk), .D (new_AGEMA_signal_4945), .Q (new_AGEMA_signal_4946) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2428 ( .C (clk), .D (new_AGEMA_signal_4948), .Q (new_AGEMA_signal_4949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2431 ( .C (clk), .D (new_AGEMA_signal_4951), .Q (new_AGEMA_signal_4952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2434 ( .C (clk), .D (new_AGEMA_signal_4954), .Q (new_AGEMA_signal_4955) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2437 ( .C (clk), .D (new_AGEMA_signal_4957), .Q (new_AGEMA_signal_4958) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2440 ( .C (clk), .D (new_AGEMA_signal_4960), .Q (new_AGEMA_signal_4961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2443 ( .C (clk), .D (new_AGEMA_signal_4963), .Q (new_AGEMA_signal_4964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2446 ( .C (clk), .D (new_AGEMA_signal_4966), .Q (new_AGEMA_signal_4967) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2449 ( .C (clk), .D (new_AGEMA_signal_4969), .Q (new_AGEMA_signal_4970) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2452 ( .C (clk), .D (new_AGEMA_signal_4972), .Q (new_AGEMA_signal_4973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2455 ( .C (clk), .D (new_AGEMA_signal_4975), .Q (new_AGEMA_signal_4976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2458 ( .C (clk), .D (new_AGEMA_signal_4978), .Q (new_AGEMA_signal_4979) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2461 ( .C (clk), .D (new_AGEMA_signal_4981), .Q (new_AGEMA_signal_4982) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2464 ( .C (clk), .D (new_AGEMA_signal_4984), .Q (new_AGEMA_signal_4985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2467 ( .C (clk), .D (new_AGEMA_signal_4987), .Q (new_AGEMA_signal_4988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2470 ( .C (clk), .D (new_AGEMA_signal_4990), .Q (new_AGEMA_signal_4991) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2473 ( .C (clk), .D (new_AGEMA_signal_4993), .Q (new_AGEMA_signal_4994) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2476 ( .C (clk), .D (new_AGEMA_signal_4996), .Q (new_AGEMA_signal_4997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2479 ( .C (clk), .D (new_AGEMA_signal_4999), .Q (new_AGEMA_signal_5000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2482 ( .C (clk), .D (new_AGEMA_signal_5002), .Q (new_AGEMA_signal_5003) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2485 ( .C (clk), .D (new_AGEMA_signal_5005), .Q (new_AGEMA_signal_5006) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2488 ( .C (clk), .D (new_AGEMA_signal_5008), .Q (new_AGEMA_signal_5009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2491 ( .C (clk), .D (new_AGEMA_signal_5011), .Q (new_AGEMA_signal_5012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2494 ( .C (clk), .D (new_AGEMA_signal_5014), .Q (new_AGEMA_signal_5015) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2497 ( .C (clk), .D (new_AGEMA_signal_5017), .Q (new_AGEMA_signal_5018) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2500 ( .C (clk), .D (new_AGEMA_signal_5020), .Q (new_AGEMA_signal_5021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2503 ( .C (clk), .D (new_AGEMA_signal_5023), .Q (new_AGEMA_signal_5024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2506 ( .C (clk), .D (new_AGEMA_signal_5026), .Q (new_AGEMA_signal_5027) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2509 ( .C (clk), .D (new_AGEMA_signal_5029), .Q (new_AGEMA_signal_5030) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2512 ( .C (clk), .D (new_AGEMA_signal_5032), .Q (new_AGEMA_signal_5033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2515 ( .C (clk), .D (new_AGEMA_signal_5035), .Q (new_AGEMA_signal_5036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2518 ( .C (clk), .D (new_AGEMA_signal_5038), .Q (new_AGEMA_signal_5039) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2521 ( .C (clk), .D (new_AGEMA_signal_5041), .Q (new_AGEMA_signal_5042) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2524 ( .C (clk), .D (new_AGEMA_signal_5044), .Q (new_AGEMA_signal_5045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2527 ( .C (clk), .D (new_AGEMA_signal_5047), .Q (new_AGEMA_signal_5048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2530 ( .C (clk), .D (new_AGEMA_signal_5050), .Q (new_AGEMA_signal_5051) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2533 ( .C (clk), .D (new_AGEMA_signal_5053), .Q (new_AGEMA_signal_5054) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2536 ( .C (clk), .D (new_AGEMA_signal_5056), .Q (new_AGEMA_signal_5057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2539 ( .C (clk), .D (new_AGEMA_signal_5059), .Q (new_AGEMA_signal_5060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2542 ( .C (clk), .D (new_AGEMA_signal_5062), .Q (new_AGEMA_signal_5063) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2545 ( .C (clk), .D (new_AGEMA_signal_5065), .Q (new_AGEMA_signal_5066) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2548 ( .C (clk), .D (new_AGEMA_signal_5068), .Q (new_AGEMA_signal_5069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2551 ( .C (clk), .D (new_AGEMA_signal_5071), .Q (new_AGEMA_signal_5072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2554 ( .C (clk), .D (new_AGEMA_signal_5074), .Q (new_AGEMA_signal_5075) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2557 ( .C (clk), .D (new_AGEMA_signal_5077), .Q (new_AGEMA_signal_5078) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2560 ( .C (clk), .D (new_AGEMA_signal_5080), .Q (new_AGEMA_signal_5081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2563 ( .C (clk), .D (new_AGEMA_signal_5083), .Q (new_AGEMA_signal_5084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2566 ( .C (clk), .D (new_AGEMA_signal_5086), .Q (new_AGEMA_signal_5087) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2569 ( .C (clk), .D (new_AGEMA_signal_5089), .Q (new_AGEMA_signal_5090) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2572 ( .C (clk), .D (new_AGEMA_signal_5092), .Q (new_AGEMA_signal_5093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2575 ( .C (clk), .D (new_AGEMA_signal_5095), .Q (new_AGEMA_signal_5096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2578 ( .C (clk), .D (new_AGEMA_signal_5098), .Q (new_AGEMA_signal_5099) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2581 ( .C (clk), .D (new_AGEMA_signal_5101), .Q (new_AGEMA_signal_5102) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2584 ( .C (clk), .D (new_AGEMA_signal_5104), .Q (new_AGEMA_signal_5105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2587 ( .C (clk), .D (new_AGEMA_signal_5107), .Q (new_AGEMA_signal_5108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2590 ( .C (clk), .D (new_AGEMA_signal_5110), .Q (new_AGEMA_signal_5111) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2593 ( .C (clk), .D (new_AGEMA_signal_5113), .Q (new_AGEMA_signal_5114) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2596 ( .C (clk), .D (new_AGEMA_signal_5116), .Q (new_AGEMA_signal_5117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2599 ( .C (clk), .D (new_AGEMA_signal_5119), .Q (new_AGEMA_signal_5120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2602 ( .C (clk), .D (new_AGEMA_signal_5122), .Q (new_AGEMA_signal_5123) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2605 ( .C (clk), .D (new_AGEMA_signal_5125), .Q (new_AGEMA_signal_5126) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2608 ( .C (clk), .D (new_AGEMA_signal_5128), .Q (new_AGEMA_signal_5129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2611 ( .C (clk), .D (new_AGEMA_signal_5131), .Q (new_AGEMA_signal_5132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2614 ( .C (clk), .D (new_AGEMA_signal_5134), .Q (new_AGEMA_signal_5135) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2617 ( .C (clk), .D (new_AGEMA_signal_5137), .Q (new_AGEMA_signal_5138) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2620 ( .C (clk), .D (new_AGEMA_signal_5140), .Q (new_AGEMA_signal_5141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2623 ( .C (clk), .D (new_AGEMA_signal_5143), .Q (new_AGEMA_signal_5144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2626 ( .C (clk), .D (new_AGEMA_signal_5146), .Q (new_AGEMA_signal_5147) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2629 ( .C (clk), .D (new_AGEMA_signal_5149), .Q (new_AGEMA_signal_5150) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2632 ( .C (clk), .D (new_AGEMA_signal_5152), .Q (new_AGEMA_signal_5153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2635 ( .C (clk), .D (new_AGEMA_signal_5155), .Q (new_AGEMA_signal_5156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2638 ( .C (clk), .D (new_AGEMA_signal_5158), .Q (new_AGEMA_signal_5159) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2641 ( .C (clk), .D (new_AGEMA_signal_5161), .Q (new_AGEMA_signal_5162) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2644 ( .C (clk), .D (new_AGEMA_signal_5164), .Q (new_AGEMA_signal_5165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2647 ( .C (clk), .D (new_AGEMA_signal_5167), .Q (new_AGEMA_signal_5168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2650 ( .C (clk), .D (new_AGEMA_signal_5170), .Q (new_AGEMA_signal_5171) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2653 ( .C (clk), .D (new_AGEMA_signal_5173), .Q (new_AGEMA_signal_5174) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2656 ( .C (clk), .D (new_AGEMA_signal_5176), .Q (new_AGEMA_signal_5177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2659 ( .C (clk), .D (new_AGEMA_signal_5179), .Q (new_AGEMA_signal_5180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2662 ( .C (clk), .D (new_AGEMA_signal_5182), .Q (new_AGEMA_signal_5183) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2665 ( .C (clk), .D (new_AGEMA_signal_5185), .Q (new_AGEMA_signal_5186) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2668 ( .C (clk), .D (new_AGEMA_signal_5188), .Q (new_AGEMA_signal_5189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2671 ( .C (clk), .D (new_AGEMA_signal_5191), .Q (new_AGEMA_signal_5192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2674 ( .C (clk), .D (new_AGEMA_signal_5194), .Q (new_AGEMA_signal_5195) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2677 ( .C (clk), .D (new_AGEMA_signal_5197), .Q (new_AGEMA_signal_5198) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2680 ( .C (clk), .D (new_AGEMA_signal_5200), .Q (new_AGEMA_signal_5201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2683 ( .C (clk), .D (new_AGEMA_signal_5203), .Q (new_AGEMA_signal_5204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2686 ( .C (clk), .D (new_AGEMA_signal_5206), .Q (new_AGEMA_signal_5207) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2689 ( .C (clk), .D (new_AGEMA_signal_5209), .Q (new_AGEMA_signal_5210) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2692 ( .C (clk), .D (new_AGEMA_signal_5212), .Q (new_AGEMA_signal_5213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2695 ( .C (clk), .D (new_AGEMA_signal_5215), .Q (new_AGEMA_signal_5216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2698 ( .C (clk), .D (new_AGEMA_signal_5218), .Q (new_AGEMA_signal_5219) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2701 ( .C (clk), .D (new_AGEMA_signal_5221), .Q (new_AGEMA_signal_5222) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2704 ( .C (clk), .D (new_AGEMA_signal_5224), .Q (new_AGEMA_signal_5225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2707 ( .C (clk), .D (new_AGEMA_signal_5227), .Q (new_AGEMA_signal_5228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2710 ( .C (clk), .D (new_AGEMA_signal_5230), .Q (new_AGEMA_signal_5231) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2713 ( .C (clk), .D (new_AGEMA_signal_5233), .Q (new_AGEMA_signal_5234) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2716 ( .C (clk), .D (new_AGEMA_signal_5236), .Q (new_AGEMA_signal_5237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2719 ( .C (clk), .D (new_AGEMA_signal_5239), .Q (new_AGEMA_signal_5240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2722 ( .C (clk), .D (new_AGEMA_signal_5242), .Q (new_AGEMA_signal_5243) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2725 ( .C (clk), .D (new_AGEMA_signal_5245), .Q (new_AGEMA_signal_5246) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2728 ( .C (clk), .D (new_AGEMA_signal_5248), .Q (new_AGEMA_signal_5249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2731 ( .C (clk), .D (new_AGEMA_signal_5251), .Q (new_AGEMA_signal_5252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2734 ( .C (clk), .D (new_AGEMA_signal_5254), .Q (new_AGEMA_signal_5255) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2737 ( .C (clk), .D (new_AGEMA_signal_5257), .Q (new_AGEMA_signal_5258) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2740 ( .C (clk), .D (new_AGEMA_signal_5260), .Q (new_AGEMA_signal_5261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2743 ( .C (clk), .D (new_AGEMA_signal_5263), .Q (new_AGEMA_signal_5264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2746 ( .C (clk), .D (new_AGEMA_signal_5266), .Q (new_AGEMA_signal_5267) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2749 ( .C (clk), .D (new_AGEMA_signal_5269), .Q (new_AGEMA_signal_5270) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2752 ( .C (clk), .D (new_AGEMA_signal_5272), .Q (new_AGEMA_signal_5273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2755 ( .C (clk), .D (new_AGEMA_signal_5275), .Q (new_AGEMA_signal_5276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2758 ( .C (clk), .D (new_AGEMA_signal_5278), .Q (new_AGEMA_signal_5279) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2761 ( .C (clk), .D (new_AGEMA_signal_5281), .Q (new_AGEMA_signal_5282) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2764 ( .C (clk), .D (new_AGEMA_signal_5284), .Q (new_AGEMA_signal_5285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2767 ( .C (clk), .D (new_AGEMA_signal_5287), .Q (new_AGEMA_signal_5288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2770 ( .C (clk), .D (new_AGEMA_signal_5290), .Q (new_AGEMA_signal_5291) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2773 ( .C (clk), .D (new_AGEMA_signal_5293), .Q (new_AGEMA_signal_5294) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2776 ( .C (clk), .D (new_AGEMA_signal_5296), .Q (new_AGEMA_signal_5297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2779 ( .C (clk), .D (new_AGEMA_signal_5299), .Q (new_AGEMA_signal_5300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2782 ( .C (clk), .D (new_AGEMA_signal_5302), .Q (new_AGEMA_signal_5303) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2785 ( .C (clk), .D (new_AGEMA_signal_5305), .Q (new_AGEMA_signal_5306) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2788 ( .C (clk), .D (new_AGEMA_signal_5308), .Q (new_AGEMA_signal_5309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2791 ( .C (clk), .D (new_AGEMA_signal_5311), .Q (new_AGEMA_signal_5312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2794 ( .C (clk), .D (new_AGEMA_signal_5314), .Q (new_AGEMA_signal_5315) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2797 ( .C (clk), .D (new_AGEMA_signal_5317), .Q (new_AGEMA_signal_5318) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2800 ( .C (clk), .D (new_AGEMA_signal_5320), .Q (new_AGEMA_signal_5321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2803 ( .C (clk), .D (new_AGEMA_signal_5323), .Q (new_AGEMA_signal_5324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2806 ( .C (clk), .D (new_AGEMA_signal_5326), .Q (new_AGEMA_signal_5327) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2809 ( .C (clk), .D (new_AGEMA_signal_5329), .Q (new_AGEMA_signal_5330) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2812 ( .C (clk), .D (new_AGEMA_signal_5332), .Q (new_AGEMA_signal_5333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2815 ( .C (clk), .D (new_AGEMA_signal_5335), .Q (new_AGEMA_signal_5336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2818 ( .C (clk), .D (new_AGEMA_signal_5338), .Q (new_AGEMA_signal_5339) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2821 ( .C (clk), .D (new_AGEMA_signal_5341), .Q (new_AGEMA_signal_5342) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2824 ( .C (clk), .D (new_AGEMA_signal_5344), .Q (new_AGEMA_signal_5345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2827 ( .C (clk), .D (new_AGEMA_signal_5347), .Q (new_AGEMA_signal_5348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2830 ( .C (clk), .D (new_AGEMA_signal_5350), .Q (new_AGEMA_signal_5351) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2833 ( .C (clk), .D (new_AGEMA_signal_5353), .Q (new_AGEMA_signal_5354) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2836 ( .C (clk), .D (new_AGEMA_signal_5356), .Q (new_AGEMA_signal_5357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2839 ( .C (clk), .D (new_AGEMA_signal_5359), .Q (new_AGEMA_signal_5360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2842 ( .C (clk), .D (new_AGEMA_signal_5362), .Q (new_AGEMA_signal_5363) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2845 ( .C (clk), .D (new_AGEMA_signal_5365), .Q (new_AGEMA_signal_5366) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2848 ( .C (clk), .D (new_AGEMA_signal_5368), .Q (new_AGEMA_signal_5369) ) ;
    buf_clk new_AGEMA_reg_buffer_2851 ( .C (clk), .D (new_AGEMA_signal_5371), .Q (new_AGEMA_signal_5372) ) ;
    buf_clk new_AGEMA_reg_buffer_2855 ( .C (clk), .D (new_AGEMA_signal_5375), .Q (new_AGEMA_signal_5376) ) ;
    buf_clk new_AGEMA_reg_buffer_2859 ( .C (clk), .D (new_AGEMA_signal_5379), .Q (new_AGEMA_signal_5380) ) ;
    buf_clk new_AGEMA_reg_buffer_2863 ( .C (clk), .D (new_AGEMA_signal_5383), .Q (new_AGEMA_signal_5384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2867 ( .C (clk), .D (new_AGEMA_signal_5387), .Q (new_AGEMA_signal_5388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2871 ( .C (clk), .D (new_AGEMA_signal_5391), .Q (new_AGEMA_signal_5392) ) ;
    buf_clk new_AGEMA_reg_buffer_2875 ( .C (clk), .D (new_AGEMA_signal_5395), .Q (new_AGEMA_signal_5396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2879 ( .C (clk), .D (new_AGEMA_signal_5399), .Q (new_AGEMA_signal_5400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2883 ( .C (clk), .D (new_AGEMA_signal_5403), .Q (new_AGEMA_signal_5404) ) ;
    buf_clk new_AGEMA_reg_buffer_2887 ( .C (clk), .D (new_AGEMA_signal_5407), .Q (new_AGEMA_signal_5408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2891 ( .C (clk), .D (new_AGEMA_signal_5411), .Q (new_AGEMA_signal_5412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2895 ( .C (clk), .D (new_AGEMA_signal_5415), .Q (new_AGEMA_signal_5416) ) ;
    buf_clk new_AGEMA_reg_buffer_2899 ( .C (clk), .D (new_AGEMA_signal_5419), .Q (new_AGEMA_signal_5420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2903 ( .C (clk), .D (new_AGEMA_signal_5423), .Q (new_AGEMA_signal_5424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2907 ( .C (clk), .D (new_AGEMA_signal_5427), .Q (new_AGEMA_signal_5428) ) ;
    buf_clk new_AGEMA_reg_buffer_2911 ( .C (clk), .D (new_AGEMA_signal_5431), .Q (new_AGEMA_signal_5432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2915 ( .C (clk), .D (new_AGEMA_signal_5435), .Q (new_AGEMA_signal_5436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2919 ( .C (clk), .D (new_AGEMA_signal_5439), .Q (new_AGEMA_signal_5440) ) ;
    buf_clk new_AGEMA_reg_buffer_2923 ( .C (clk), .D (new_AGEMA_signal_5443), .Q (new_AGEMA_signal_5444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2927 ( .C (clk), .D (new_AGEMA_signal_5447), .Q (new_AGEMA_signal_5448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2931 ( .C (clk), .D (new_AGEMA_signal_5451), .Q (new_AGEMA_signal_5452) ) ;
    buf_clk new_AGEMA_reg_buffer_2935 ( .C (clk), .D (new_AGEMA_signal_5455), .Q (new_AGEMA_signal_5456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2939 ( .C (clk), .D (new_AGEMA_signal_5459), .Q (new_AGEMA_signal_5460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2943 ( .C (clk), .D (new_AGEMA_signal_5463), .Q (new_AGEMA_signal_5464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2947 ( .C (clk), .D (new_AGEMA_signal_5467), .Q (new_AGEMA_signal_5468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2951 ( .C (clk), .D (new_AGEMA_signal_5471), .Q (new_AGEMA_signal_5472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2955 ( .C (clk), .D (new_AGEMA_signal_5475), .Q (new_AGEMA_signal_5476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2959 ( .C (clk), .D (new_AGEMA_signal_5479), .Q (new_AGEMA_signal_5480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2963 ( .C (clk), .D (new_AGEMA_signal_5483), .Q (new_AGEMA_signal_5484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2967 ( .C (clk), .D (new_AGEMA_signal_5487), .Q (new_AGEMA_signal_5488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2971 ( .C (clk), .D (new_AGEMA_signal_5491), .Q (new_AGEMA_signal_5492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2975 ( .C (clk), .D (new_AGEMA_signal_5495), .Q (new_AGEMA_signal_5496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2979 ( .C (clk), .D (new_AGEMA_signal_5499), .Q (new_AGEMA_signal_5500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2983 ( .C (clk), .D (new_AGEMA_signal_5503), .Q (new_AGEMA_signal_5504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2987 ( .C (clk), .D (new_AGEMA_signal_5507), .Q (new_AGEMA_signal_5508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2991 ( .C (clk), .D (new_AGEMA_signal_5511), .Q (new_AGEMA_signal_5512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2995 ( .C (clk), .D (new_AGEMA_signal_5515), .Q (new_AGEMA_signal_5516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2999 ( .C (clk), .D (new_AGEMA_signal_5519), .Q (new_AGEMA_signal_5520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3003 ( .C (clk), .D (new_AGEMA_signal_5523), .Q (new_AGEMA_signal_5524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3007 ( .C (clk), .D (new_AGEMA_signal_5527), .Q (new_AGEMA_signal_5528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3011 ( .C (clk), .D (new_AGEMA_signal_5531), .Q (new_AGEMA_signal_5532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3015 ( .C (clk), .D (new_AGEMA_signal_5535), .Q (new_AGEMA_signal_5536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3019 ( .C (clk), .D (new_AGEMA_signal_5539), .Q (new_AGEMA_signal_5540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3023 ( .C (clk), .D (new_AGEMA_signal_5543), .Q (new_AGEMA_signal_5544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3027 ( .C (clk), .D (new_AGEMA_signal_5547), .Q (new_AGEMA_signal_5548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3031 ( .C (clk), .D (new_AGEMA_signal_5551), .Q (new_AGEMA_signal_5552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3035 ( .C (clk), .D (new_AGEMA_signal_5555), .Q (new_AGEMA_signal_5556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3039 ( .C (clk), .D (new_AGEMA_signal_5559), .Q (new_AGEMA_signal_5560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3043 ( .C (clk), .D (new_AGEMA_signal_5563), .Q (new_AGEMA_signal_5564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3047 ( .C (clk), .D (new_AGEMA_signal_5567), .Q (new_AGEMA_signal_5568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3051 ( .C (clk), .D (new_AGEMA_signal_5571), .Q (new_AGEMA_signal_5572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3055 ( .C (clk), .D (new_AGEMA_signal_5575), .Q (new_AGEMA_signal_5576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3059 ( .C (clk), .D (new_AGEMA_signal_5579), .Q (new_AGEMA_signal_5580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3063 ( .C (clk), .D (new_AGEMA_signal_5583), .Q (new_AGEMA_signal_5584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3067 ( .C (clk), .D (new_AGEMA_signal_5587), .Q (new_AGEMA_signal_5588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3071 ( .C (clk), .D (new_AGEMA_signal_5591), .Q (new_AGEMA_signal_5592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3075 ( .C (clk), .D (new_AGEMA_signal_5595), .Q (new_AGEMA_signal_5596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3079 ( .C (clk), .D (new_AGEMA_signal_5599), .Q (new_AGEMA_signal_5600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3083 ( .C (clk), .D (new_AGEMA_signal_5603), .Q (new_AGEMA_signal_5604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3087 ( .C (clk), .D (new_AGEMA_signal_5607), .Q (new_AGEMA_signal_5608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3091 ( .C (clk), .D (new_AGEMA_signal_5611), .Q (new_AGEMA_signal_5612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3095 ( .C (clk), .D (new_AGEMA_signal_5615), .Q (new_AGEMA_signal_5616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3099 ( .C (clk), .D (new_AGEMA_signal_5619), .Q (new_AGEMA_signal_5620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3103 ( .C (clk), .D (new_AGEMA_signal_5623), .Q (new_AGEMA_signal_5624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3107 ( .C (clk), .D (new_AGEMA_signal_5627), .Q (new_AGEMA_signal_5628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3111 ( .C (clk), .D (new_AGEMA_signal_5631), .Q (new_AGEMA_signal_5632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3115 ( .C (clk), .D (new_AGEMA_signal_5635), .Q (new_AGEMA_signal_5636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3119 ( .C (clk), .D (new_AGEMA_signal_5639), .Q (new_AGEMA_signal_5640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3123 ( .C (clk), .D (new_AGEMA_signal_5643), .Q (new_AGEMA_signal_5644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3127 ( .C (clk), .D (new_AGEMA_signal_5647), .Q (new_AGEMA_signal_5648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3131 ( .C (clk), .D (new_AGEMA_signal_5651), .Q (new_AGEMA_signal_5652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3135 ( .C (clk), .D (new_AGEMA_signal_5655), .Q (new_AGEMA_signal_5656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3139 ( .C (clk), .D (new_AGEMA_signal_5659), .Q (new_AGEMA_signal_5660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3143 ( .C (clk), .D (new_AGEMA_signal_5663), .Q (new_AGEMA_signal_5664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3147 ( .C (clk), .D (new_AGEMA_signal_5667), .Q (new_AGEMA_signal_5668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3151 ( .C (clk), .D (new_AGEMA_signal_5671), .Q (new_AGEMA_signal_5672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3155 ( .C (clk), .D (new_AGEMA_signal_5675), .Q (new_AGEMA_signal_5676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3159 ( .C (clk), .D (new_AGEMA_signal_5679), .Q (new_AGEMA_signal_5680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3163 ( .C (clk), .D (new_AGEMA_signal_5683), .Q (new_AGEMA_signal_5684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3167 ( .C (clk), .D (new_AGEMA_signal_5687), .Q (new_AGEMA_signal_5688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3171 ( .C (clk), .D (new_AGEMA_signal_5691), .Q (new_AGEMA_signal_5692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3175 ( .C (clk), .D (new_AGEMA_signal_5695), .Q (new_AGEMA_signal_5696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3179 ( .C (clk), .D (new_AGEMA_signal_5699), .Q (new_AGEMA_signal_5700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3183 ( .C (clk), .D (new_AGEMA_signal_5703), .Q (new_AGEMA_signal_5704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3187 ( .C (clk), .D (new_AGEMA_signal_5707), .Q (new_AGEMA_signal_5708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3191 ( .C (clk), .D (new_AGEMA_signal_5711), .Q (new_AGEMA_signal_5712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3195 ( .C (clk), .D (new_AGEMA_signal_5715), .Q (new_AGEMA_signal_5716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3199 ( .C (clk), .D (new_AGEMA_signal_5719), .Q (new_AGEMA_signal_5720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3203 ( .C (clk), .D (new_AGEMA_signal_5723), .Q (new_AGEMA_signal_5724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3207 ( .C (clk), .D (new_AGEMA_signal_5727), .Q (new_AGEMA_signal_5728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3211 ( .C (clk), .D (new_AGEMA_signal_5731), .Q (new_AGEMA_signal_5732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3215 ( .C (clk), .D (new_AGEMA_signal_5735), .Q (new_AGEMA_signal_5736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3219 ( .C (clk), .D (new_AGEMA_signal_5739), .Q (new_AGEMA_signal_5740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3223 ( .C (clk), .D (new_AGEMA_signal_5743), .Q (new_AGEMA_signal_5744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3227 ( .C (clk), .D (new_AGEMA_signal_5747), .Q (new_AGEMA_signal_5748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3231 ( .C (clk), .D (new_AGEMA_signal_5751), .Q (new_AGEMA_signal_5752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3235 ( .C (clk), .D (new_AGEMA_signal_5755), .Q (new_AGEMA_signal_5756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3239 ( .C (clk), .D (new_AGEMA_signal_5759), .Q (new_AGEMA_signal_5760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3243 ( .C (clk), .D (new_AGEMA_signal_5763), .Q (new_AGEMA_signal_5764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3247 ( .C (clk), .D (new_AGEMA_signal_5767), .Q (new_AGEMA_signal_5768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3251 ( .C (clk), .D (new_AGEMA_signal_5771), .Q (new_AGEMA_signal_5772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3255 ( .C (clk), .D (new_AGEMA_signal_5775), .Q (new_AGEMA_signal_5776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3259 ( .C (clk), .D (new_AGEMA_signal_5779), .Q (new_AGEMA_signal_5780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3263 ( .C (clk), .D (new_AGEMA_signal_5783), .Q (new_AGEMA_signal_5784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3267 ( .C (clk), .D (new_AGEMA_signal_5787), .Q (new_AGEMA_signal_5788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3271 ( .C (clk), .D (new_AGEMA_signal_5791), .Q (new_AGEMA_signal_5792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3275 ( .C (clk), .D (new_AGEMA_signal_5795), .Q (new_AGEMA_signal_5796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3279 ( .C (clk), .D (new_AGEMA_signal_5799), .Q (new_AGEMA_signal_5800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3283 ( .C (clk), .D (new_AGEMA_signal_5803), .Q (new_AGEMA_signal_5804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3287 ( .C (clk), .D (new_AGEMA_signal_5807), .Q (new_AGEMA_signal_5808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3291 ( .C (clk), .D (new_AGEMA_signal_5811), .Q (new_AGEMA_signal_5812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3295 ( .C (clk), .D (new_AGEMA_signal_5815), .Q (new_AGEMA_signal_5816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3299 ( .C (clk), .D (new_AGEMA_signal_5819), .Q (new_AGEMA_signal_5820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3303 ( .C (clk), .D (new_AGEMA_signal_5823), .Q (new_AGEMA_signal_5824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3307 ( .C (clk), .D (new_AGEMA_signal_5827), .Q (new_AGEMA_signal_5828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3311 ( .C (clk), .D (new_AGEMA_signal_5831), .Q (new_AGEMA_signal_5832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3315 ( .C (clk), .D (new_AGEMA_signal_5835), .Q (new_AGEMA_signal_5836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3319 ( .C (clk), .D (new_AGEMA_signal_5839), .Q (new_AGEMA_signal_5840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3323 ( .C (clk), .D (new_AGEMA_signal_5843), .Q (new_AGEMA_signal_5844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3327 ( .C (clk), .D (new_AGEMA_signal_5847), .Q (new_AGEMA_signal_5848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3331 ( .C (clk), .D (new_AGEMA_signal_5851), .Q (new_AGEMA_signal_5852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3335 ( .C (clk), .D (new_AGEMA_signal_5855), .Q (new_AGEMA_signal_5856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3339 ( .C (clk), .D (new_AGEMA_signal_5859), .Q (new_AGEMA_signal_5860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3343 ( .C (clk), .D (new_AGEMA_signal_5863), .Q (new_AGEMA_signal_5864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3347 ( .C (clk), .D (new_AGEMA_signal_5867), .Q (new_AGEMA_signal_5868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3351 ( .C (clk), .D (new_AGEMA_signal_5871), .Q (new_AGEMA_signal_5872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3355 ( .C (clk), .D (new_AGEMA_signal_5875), .Q (new_AGEMA_signal_5876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3359 ( .C (clk), .D (new_AGEMA_signal_5879), .Q (new_AGEMA_signal_5880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3363 ( .C (clk), .D (new_AGEMA_signal_5883), .Q (new_AGEMA_signal_5884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3367 ( .C (clk), .D (new_AGEMA_signal_5887), .Q (new_AGEMA_signal_5888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3371 ( .C (clk), .D (new_AGEMA_signal_5891), .Q (new_AGEMA_signal_5892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3375 ( .C (clk), .D (new_AGEMA_signal_5895), .Q (new_AGEMA_signal_5896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3379 ( .C (clk), .D (new_AGEMA_signal_5899), .Q (new_AGEMA_signal_5900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3383 ( .C (clk), .D (new_AGEMA_signal_5903), .Q (new_AGEMA_signal_5904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3387 ( .C (clk), .D (new_AGEMA_signal_5907), .Q (new_AGEMA_signal_5908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3391 ( .C (clk), .D (new_AGEMA_signal_5911), .Q (new_AGEMA_signal_5912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3395 ( .C (clk), .D (new_AGEMA_signal_5915), .Q (new_AGEMA_signal_5916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3399 ( .C (clk), .D (new_AGEMA_signal_5919), .Q (new_AGEMA_signal_5920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3403 ( .C (clk), .D (new_AGEMA_signal_5923), .Q (new_AGEMA_signal_5924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3407 ( .C (clk), .D (new_AGEMA_signal_5927), .Q (new_AGEMA_signal_5928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3411 ( .C (clk), .D (new_AGEMA_signal_5931), .Q (new_AGEMA_signal_5932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3415 ( .C (clk), .D (new_AGEMA_signal_5935), .Q (new_AGEMA_signal_5936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3419 ( .C (clk), .D (new_AGEMA_signal_5939), .Q (new_AGEMA_signal_5940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3423 ( .C (clk), .D (new_AGEMA_signal_5943), .Q (new_AGEMA_signal_5944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3427 ( .C (clk), .D (new_AGEMA_signal_5947), .Q (new_AGEMA_signal_5948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3431 ( .C (clk), .D (new_AGEMA_signal_5951), .Q (new_AGEMA_signal_5952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3435 ( .C (clk), .D (new_AGEMA_signal_5955), .Q (new_AGEMA_signal_5956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3439 ( .C (clk), .D (new_AGEMA_signal_5959), .Q (new_AGEMA_signal_5960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3443 ( .C (clk), .D (new_AGEMA_signal_5963), .Q (new_AGEMA_signal_5964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3447 ( .C (clk), .D (new_AGEMA_signal_5967), .Q (new_AGEMA_signal_5968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3451 ( .C (clk), .D (new_AGEMA_signal_5971), .Q (new_AGEMA_signal_5972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3455 ( .C (clk), .D (new_AGEMA_signal_5975), .Q (new_AGEMA_signal_5976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3459 ( .C (clk), .D (new_AGEMA_signal_5979), .Q (new_AGEMA_signal_5980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3463 ( .C (clk), .D (new_AGEMA_signal_5983), .Q (new_AGEMA_signal_5984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3467 ( .C (clk), .D (new_AGEMA_signal_5987), .Q (new_AGEMA_signal_5988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3471 ( .C (clk), .D (new_AGEMA_signal_5991), .Q (new_AGEMA_signal_5992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3475 ( .C (clk), .D (new_AGEMA_signal_5995), .Q (new_AGEMA_signal_5996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3479 ( .C (clk), .D (new_AGEMA_signal_5999), .Q (new_AGEMA_signal_6000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3483 ( .C (clk), .D (new_AGEMA_signal_6003), .Q (new_AGEMA_signal_6004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3487 ( .C (clk), .D (new_AGEMA_signal_6007), .Q (new_AGEMA_signal_6008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3491 ( .C (clk), .D (new_AGEMA_signal_6011), .Q (new_AGEMA_signal_6012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3495 ( .C (clk), .D (new_AGEMA_signal_6015), .Q (new_AGEMA_signal_6016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3499 ( .C (clk), .D (new_AGEMA_signal_6019), .Q (new_AGEMA_signal_6020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3503 ( .C (clk), .D (new_AGEMA_signal_6023), .Q (new_AGEMA_signal_6024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3507 ( .C (clk), .D (new_AGEMA_signal_6027), .Q (new_AGEMA_signal_6028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3511 ( .C (clk), .D (new_AGEMA_signal_6031), .Q (new_AGEMA_signal_6032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3515 ( .C (clk), .D (new_AGEMA_signal_6035), .Q (new_AGEMA_signal_6036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3519 ( .C (clk), .D (new_AGEMA_signal_6039), .Q (new_AGEMA_signal_6040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3523 ( .C (clk), .D (new_AGEMA_signal_6043), .Q (new_AGEMA_signal_6044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3527 ( .C (clk), .D (new_AGEMA_signal_6047), .Q (new_AGEMA_signal_6048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3531 ( .C (clk), .D (new_AGEMA_signal_6051), .Q (new_AGEMA_signal_6052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3535 ( .C (clk), .D (new_AGEMA_signal_6055), .Q (new_AGEMA_signal_6056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3539 ( .C (clk), .D (new_AGEMA_signal_6059), .Q (new_AGEMA_signal_6060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3543 ( .C (clk), .D (new_AGEMA_signal_6063), .Q (new_AGEMA_signal_6064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3547 ( .C (clk), .D (new_AGEMA_signal_6067), .Q (new_AGEMA_signal_6068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3551 ( .C (clk), .D (new_AGEMA_signal_6071), .Q (new_AGEMA_signal_6072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3555 ( .C (clk), .D (new_AGEMA_signal_6075), .Q (new_AGEMA_signal_6076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3559 ( .C (clk), .D (new_AGEMA_signal_6079), .Q (new_AGEMA_signal_6080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3563 ( .C (clk), .D (new_AGEMA_signal_6083), .Q (new_AGEMA_signal_6084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3567 ( .C (clk), .D (new_AGEMA_signal_6087), .Q (new_AGEMA_signal_6088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3571 ( .C (clk), .D (new_AGEMA_signal_6091), .Q (new_AGEMA_signal_6092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3575 ( .C (clk), .D (new_AGEMA_signal_6095), .Q (new_AGEMA_signal_6096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3579 ( .C (clk), .D (new_AGEMA_signal_6099), .Q (new_AGEMA_signal_6100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3583 ( .C (clk), .D (new_AGEMA_signal_6103), .Q (new_AGEMA_signal_6104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3587 ( .C (clk), .D (new_AGEMA_signal_6107), .Q (new_AGEMA_signal_6108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3591 ( .C (clk), .D (new_AGEMA_signal_6111), .Q (new_AGEMA_signal_6112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3595 ( .C (clk), .D (new_AGEMA_signal_6115), .Q (new_AGEMA_signal_6116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3599 ( .C (clk), .D (new_AGEMA_signal_6119), .Q (new_AGEMA_signal_6120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3603 ( .C (clk), .D (new_AGEMA_signal_6123), .Q (new_AGEMA_signal_6124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3607 ( .C (clk), .D (new_AGEMA_signal_6127), .Q (new_AGEMA_signal_6128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3611 ( .C (clk), .D (new_AGEMA_signal_6131), .Q (new_AGEMA_signal_6132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3615 ( .C (clk), .D (new_AGEMA_signal_6135), .Q (new_AGEMA_signal_6136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3619 ( .C (clk), .D (new_AGEMA_signal_6139), .Q (new_AGEMA_signal_6140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3623 ( .C (clk), .D (new_AGEMA_signal_6143), .Q (new_AGEMA_signal_6144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3627 ( .C (clk), .D (new_AGEMA_signal_6147), .Q (new_AGEMA_signal_6148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3631 ( .C (clk), .D (new_AGEMA_signal_6151), .Q (new_AGEMA_signal_6152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3635 ( .C (clk), .D (new_AGEMA_signal_6155), .Q (new_AGEMA_signal_6156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3639 ( .C (clk), .D (new_AGEMA_signal_6159), .Q (new_AGEMA_signal_6160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3643 ( .C (clk), .D (new_AGEMA_signal_6163), .Q (new_AGEMA_signal_6164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3647 ( .C (clk), .D (new_AGEMA_signal_6167), .Q (new_AGEMA_signal_6168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3651 ( .C (clk), .D (new_AGEMA_signal_6171), .Q (new_AGEMA_signal_6172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3655 ( .C (clk), .D (new_AGEMA_signal_6175), .Q (new_AGEMA_signal_6176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3659 ( .C (clk), .D (new_AGEMA_signal_6179), .Q (new_AGEMA_signal_6180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3663 ( .C (clk), .D (new_AGEMA_signal_6183), .Q (new_AGEMA_signal_6184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3667 ( .C (clk), .D (new_AGEMA_signal_6187), .Q (new_AGEMA_signal_6188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3671 ( .C (clk), .D (new_AGEMA_signal_6191), .Q (new_AGEMA_signal_6192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3675 ( .C (clk), .D (new_AGEMA_signal_6195), .Q (new_AGEMA_signal_6196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3679 ( .C (clk), .D (new_AGEMA_signal_6199), .Q (new_AGEMA_signal_6200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3683 ( .C (clk), .D (new_AGEMA_signal_6203), .Q (new_AGEMA_signal_6204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3687 ( .C (clk), .D (new_AGEMA_signal_6207), .Q (new_AGEMA_signal_6208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3691 ( .C (clk), .D (new_AGEMA_signal_6211), .Q (new_AGEMA_signal_6212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3695 ( .C (clk), .D (new_AGEMA_signal_6215), .Q (new_AGEMA_signal_6216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3699 ( .C (clk), .D (new_AGEMA_signal_6219), .Q (new_AGEMA_signal_6220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3703 ( .C (clk), .D (new_AGEMA_signal_6223), .Q (new_AGEMA_signal_6224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3707 ( .C (clk), .D (new_AGEMA_signal_6227), .Q (new_AGEMA_signal_6228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3711 ( .C (clk), .D (new_AGEMA_signal_6231), .Q (new_AGEMA_signal_6232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3715 ( .C (clk), .D (new_AGEMA_signal_6235), .Q (new_AGEMA_signal_6236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3719 ( .C (clk), .D (new_AGEMA_signal_6239), .Q (new_AGEMA_signal_6240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3723 ( .C (clk), .D (new_AGEMA_signal_6243), .Q (new_AGEMA_signal_6244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3727 ( .C (clk), .D (new_AGEMA_signal_6247), .Q (new_AGEMA_signal_6248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3731 ( .C (clk), .D (new_AGEMA_signal_6251), .Q (new_AGEMA_signal_6252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3735 ( .C (clk), .D (new_AGEMA_signal_6255), .Q (new_AGEMA_signal_6256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3739 ( .C (clk), .D (new_AGEMA_signal_6259), .Q (new_AGEMA_signal_6260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3743 ( .C (clk), .D (new_AGEMA_signal_6263), .Q (new_AGEMA_signal_6264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3747 ( .C (clk), .D (new_AGEMA_signal_6267), .Q (new_AGEMA_signal_6268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3751 ( .C (clk), .D (new_AGEMA_signal_6271), .Q (new_AGEMA_signal_6272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3755 ( .C (clk), .D (new_AGEMA_signal_6275), .Q (new_AGEMA_signal_6276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3759 ( .C (clk), .D (new_AGEMA_signal_6279), .Q (new_AGEMA_signal_6280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3763 ( .C (clk), .D (new_AGEMA_signal_6283), .Q (new_AGEMA_signal_6284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3767 ( .C (clk), .D (new_AGEMA_signal_6287), .Q (new_AGEMA_signal_6288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3771 ( .C (clk), .D (new_AGEMA_signal_6291), .Q (new_AGEMA_signal_6292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3775 ( .C (clk), .D (new_AGEMA_signal_6295), .Q (new_AGEMA_signal_6296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3779 ( .C (clk), .D (new_AGEMA_signal_6299), .Q (new_AGEMA_signal_6300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3783 ( .C (clk), .D (new_AGEMA_signal_6303), .Q (new_AGEMA_signal_6304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3787 ( .C (clk), .D (new_AGEMA_signal_6307), .Q (new_AGEMA_signal_6308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3791 ( .C (clk), .D (new_AGEMA_signal_6311), .Q (new_AGEMA_signal_6312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3795 ( .C (clk), .D (new_AGEMA_signal_6315), .Q (new_AGEMA_signal_6316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3799 ( .C (clk), .D (new_AGEMA_signal_6319), .Q (new_AGEMA_signal_6320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3803 ( .C (clk), .D (new_AGEMA_signal_6323), .Q (new_AGEMA_signal_6324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3807 ( .C (clk), .D (new_AGEMA_signal_6327), .Q (new_AGEMA_signal_6328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3811 ( .C (clk), .D (new_AGEMA_signal_6331), .Q (new_AGEMA_signal_6332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3815 ( .C (clk), .D (new_AGEMA_signal_6335), .Q (new_AGEMA_signal_6336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3819 ( .C (clk), .D (new_AGEMA_signal_6339), .Q (new_AGEMA_signal_6340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3823 ( .C (clk), .D (new_AGEMA_signal_6343), .Q (new_AGEMA_signal_6344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3827 ( .C (clk), .D (new_AGEMA_signal_6347), .Q (new_AGEMA_signal_6348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3831 ( .C (clk), .D (new_AGEMA_signal_6351), .Q (new_AGEMA_signal_6352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3835 ( .C (clk), .D (new_AGEMA_signal_6355), .Q (new_AGEMA_signal_6356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3839 ( .C (clk), .D (new_AGEMA_signal_6359), .Q (new_AGEMA_signal_6360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3843 ( .C (clk), .D (new_AGEMA_signal_6363), .Q (new_AGEMA_signal_6364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3847 ( .C (clk), .D (new_AGEMA_signal_6367), .Q (new_AGEMA_signal_6368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3851 ( .C (clk), .D (new_AGEMA_signal_6371), .Q (new_AGEMA_signal_6372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3855 ( .C (clk), .D (new_AGEMA_signal_6375), .Q (new_AGEMA_signal_6376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3859 ( .C (clk), .D (new_AGEMA_signal_6379), .Q (new_AGEMA_signal_6380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3863 ( .C (clk), .D (new_AGEMA_signal_6383), .Q (new_AGEMA_signal_6384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3867 ( .C (clk), .D (new_AGEMA_signal_6387), .Q (new_AGEMA_signal_6388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3871 ( .C (clk), .D (new_AGEMA_signal_6391), .Q (new_AGEMA_signal_6392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3875 ( .C (clk), .D (new_AGEMA_signal_6395), .Q (new_AGEMA_signal_6396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3879 ( .C (clk), .D (new_AGEMA_signal_6399), .Q (new_AGEMA_signal_6400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3883 ( .C (clk), .D (new_AGEMA_signal_6403), .Q (new_AGEMA_signal_6404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3887 ( .C (clk), .D (new_AGEMA_signal_6407), .Q (new_AGEMA_signal_6408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3891 ( .C (clk), .D (new_AGEMA_signal_6411), .Q (new_AGEMA_signal_6412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3895 ( .C (clk), .D (new_AGEMA_signal_6415), .Q (new_AGEMA_signal_6416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3899 ( .C (clk), .D (new_AGEMA_signal_6419), .Q (new_AGEMA_signal_6420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3903 ( .C (clk), .D (new_AGEMA_signal_6423), .Q (new_AGEMA_signal_6424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3907 ( .C (clk), .D (new_AGEMA_signal_6427), .Q (new_AGEMA_signal_6428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3911 ( .C (clk), .D (new_AGEMA_signal_6431), .Q (new_AGEMA_signal_6432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3915 ( .C (clk), .D (new_AGEMA_signal_6435), .Q (new_AGEMA_signal_6436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3919 ( .C (clk), .D (new_AGEMA_signal_6439), .Q (new_AGEMA_signal_6440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3923 ( .C (clk), .D (new_AGEMA_signal_6443), .Q (new_AGEMA_signal_6444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3927 ( .C (clk), .D (new_AGEMA_signal_6447), .Q (new_AGEMA_signal_6448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3931 ( .C (clk), .D (new_AGEMA_signal_6451), .Q (new_AGEMA_signal_6452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3935 ( .C (clk), .D (new_AGEMA_signal_6455), .Q (new_AGEMA_signal_6456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3939 ( .C (clk), .D (new_AGEMA_signal_6459), .Q (new_AGEMA_signal_6460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3943 ( .C (clk), .D (new_AGEMA_signal_6463), .Q (new_AGEMA_signal_6464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3947 ( .C (clk), .D (new_AGEMA_signal_6467), .Q (new_AGEMA_signal_6468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3951 ( .C (clk), .D (new_AGEMA_signal_6471), .Q (new_AGEMA_signal_6472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3955 ( .C (clk), .D (new_AGEMA_signal_6475), .Q (new_AGEMA_signal_6476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3959 ( .C (clk), .D (new_AGEMA_signal_6479), .Q (new_AGEMA_signal_6480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3963 ( .C (clk), .D (new_AGEMA_signal_6483), .Q (new_AGEMA_signal_6484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3967 ( .C (clk), .D (new_AGEMA_signal_6487), .Q (new_AGEMA_signal_6488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3971 ( .C (clk), .D (new_AGEMA_signal_6491), .Q (new_AGEMA_signal_6492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3975 ( .C (clk), .D (new_AGEMA_signal_6495), .Q (new_AGEMA_signal_6496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3979 ( .C (clk), .D (new_AGEMA_signal_6499), .Q (new_AGEMA_signal_6500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3983 ( .C (clk), .D (new_AGEMA_signal_6503), .Q (new_AGEMA_signal_6504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3987 ( .C (clk), .D (new_AGEMA_signal_6507), .Q (new_AGEMA_signal_6508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3991 ( .C (clk), .D (new_AGEMA_signal_6511), .Q (new_AGEMA_signal_6512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3995 ( .C (clk), .D (new_AGEMA_signal_6515), .Q (new_AGEMA_signal_6516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3999 ( .C (clk), .D (new_AGEMA_signal_6519), .Q (new_AGEMA_signal_6520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4003 ( .C (clk), .D (new_AGEMA_signal_6523), .Q (new_AGEMA_signal_6524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4007 ( .C (clk), .D (new_AGEMA_signal_6527), .Q (new_AGEMA_signal_6528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4011 ( .C (clk), .D (new_AGEMA_signal_6531), .Q (new_AGEMA_signal_6532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4015 ( .C (clk), .D (new_AGEMA_signal_6535), .Q (new_AGEMA_signal_6536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4019 ( .C (clk), .D (new_AGEMA_signal_6539), .Q (new_AGEMA_signal_6540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4023 ( .C (clk), .D (new_AGEMA_signal_6543), .Q (new_AGEMA_signal_6544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4027 ( .C (clk), .D (new_AGEMA_signal_6547), .Q (new_AGEMA_signal_6548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4031 ( .C (clk), .D (new_AGEMA_signal_6551), .Q (new_AGEMA_signal_6552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4035 ( .C (clk), .D (new_AGEMA_signal_6555), .Q (new_AGEMA_signal_6556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4039 ( .C (clk), .D (new_AGEMA_signal_6559), .Q (new_AGEMA_signal_6560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4043 ( .C (clk), .D (new_AGEMA_signal_6563), .Q (new_AGEMA_signal_6564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4047 ( .C (clk), .D (new_AGEMA_signal_6567), .Q (new_AGEMA_signal_6568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4051 ( .C (clk), .D (new_AGEMA_signal_6571), .Q (new_AGEMA_signal_6572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4055 ( .C (clk), .D (new_AGEMA_signal_6575), .Q (new_AGEMA_signal_6576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4059 ( .C (clk), .D (new_AGEMA_signal_6579), .Q (new_AGEMA_signal_6580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4063 ( .C (clk), .D (new_AGEMA_signal_6583), .Q (new_AGEMA_signal_6584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4067 ( .C (clk), .D (new_AGEMA_signal_6587), .Q (new_AGEMA_signal_6588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4071 ( .C (clk), .D (new_AGEMA_signal_6591), .Q (new_AGEMA_signal_6592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4075 ( .C (clk), .D (new_AGEMA_signal_6595), .Q (new_AGEMA_signal_6596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4079 ( .C (clk), .D (new_AGEMA_signal_6599), .Q (new_AGEMA_signal_6600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4083 ( .C (clk), .D (new_AGEMA_signal_6603), .Q (new_AGEMA_signal_6604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4087 ( .C (clk), .D (new_AGEMA_signal_6607), .Q (new_AGEMA_signal_6608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4091 ( .C (clk), .D (new_AGEMA_signal_6611), .Q (new_AGEMA_signal_6612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4095 ( .C (clk), .D (new_AGEMA_signal_6615), .Q (new_AGEMA_signal_6616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4099 ( .C (clk), .D (new_AGEMA_signal_6619), .Q (new_AGEMA_signal_6620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4103 ( .C (clk), .D (new_AGEMA_signal_6623), .Q (new_AGEMA_signal_6624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4107 ( .C (clk), .D (new_AGEMA_signal_6627), .Q (new_AGEMA_signal_6628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4111 ( .C (clk), .D (new_AGEMA_signal_6631), .Q (new_AGEMA_signal_6632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4115 ( .C (clk), .D (new_AGEMA_signal_6635), .Q (new_AGEMA_signal_6636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4119 ( .C (clk), .D (new_AGEMA_signal_6639), .Q (new_AGEMA_signal_6640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4123 ( .C (clk), .D (new_AGEMA_signal_6643), .Q (new_AGEMA_signal_6644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4127 ( .C (clk), .D (new_AGEMA_signal_6647), .Q (new_AGEMA_signal_6648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4131 ( .C (clk), .D (new_AGEMA_signal_6651), .Q (new_AGEMA_signal_6652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4135 ( .C (clk), .D (new_AGEMA_signal_6655), .Q (new_AGEMA_signal_6656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4139 ( .C (clk), .D (new_AGEMA_signal_6659), .Q (new_AGEMA_signal_6660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4143 ( .C (clk), .D (new_AGEMA_signal_6663), .Q (new_AGEMA_signal_6664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4147 ( .C (clk), .D (new_AGEMA_signal_6667), .Q (new_AGEMA_signal_6668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4151 ( .C (clk), .D (new_AGEMA_signal_6671), .Q (new_AGEMA_signal_6672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4155 ( .C (clk), .D (new_AGEMA_signal_6675), .Q (new_AGEMA_signal_6676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4159 ( .C (clk), .D (new_AGEMA_signal_6679), .Q (new_AGEMA_signal_6680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4163 ( .C (clk), .D (new_AGEMA_signal_6683), .Q (new_AGEMA_signal_6684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4167 ( .C (clk), .D (new_AGEMA_signal_6687), .Q (new_AGEMA_signal_6688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4171 ( .C (clk), .D (new_AGEMA_signal_6691), .Q (new_AGEMA_signal_6692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4175 ( .C (clk), .D (new_AGEMA_signal_6695), .Q (new_AGEMA_signal_6696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4179 ( .C (clk), .D (new_AGEMA_signal_6699), .Q (new_AGEMA_signal_6700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4183 ( .C (clk), .D (new_AGEMA_signal_6703), .Q (new_AGEMA_signal_6704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4187 ( .C (clk), .D (new_AGEMA_signal_6707), .Q (new_AGEMA_signal_6708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4191 ( .C (clk), .D (new_AGEMA_signal_6711), .Q (new_AGEMA_signal_6712) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4195 ( .C (clk), .D (new_AGEMA_signal_6715), .Q (new_AGEMA_signal_6716) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4199 ( .C (clk), .D (new_AGEMA_signal_6719), .Q (new_AGEMA_signal_6720) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4203 ( .C (clk), .D (new_AGEMA_signal_6723), .Q (new_AGEMA_signal_6724) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4207 ( .C (clk), .D (new_AGEMA_signal_6727), .Q (new_AGEMA_signal_6728) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4211 ( .C (clk), .D (new_AGEMA_signal_6731), .Q (new_AGEMA_signal_6732) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4215 ( .C (clk), .D (new_AGEMA_signal_6735), .Q (new_AGEMA_signal_6736) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4219 ( .C (clk), .D (new_AGEMA_signal_6739), .Q (new_AGEMA_signal_6740) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4223 ( .C (clk), .D (new_AGEMA_signal_6743), .Q (new_AGEMA_signal_6744) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4227 ( .C (clk), .D (new_AGEMA_signal_6747), .Q (new_AGEMA_signal_6748) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4231 ( .C (clk), .D (new_AGEMA_signal_6751), .Q (new_AGEMA_signal_6752) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4235 ( .C (clk), .D (new_AGEMA_signal_6755), .Q (new_AGEMA_signal_6756) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4239 ( .C (clk), .D (new_AGEMA_signal_6759), .Q (new_AGEMA_signal_6760) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4243 ( .C (clk), .D (new_AGEMA_signal_6763), .Q (new_AGEMA_signal_6764) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4247 ( .C (clk), .D (new_AGEMA_signal_6767), .Q (new_AGEMA_signal_6768) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4251 ( .C (clk), .D (new_AGEMA_signal_6771), .Q (new_AGEMA_signal_6772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4255 ( .C (clk), .D (new_AGEMA_signal_6775), .Q (new_AGEMA_signal_6776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4259 ( .C (clk), .D (new_AGEMA_signal_6779), .Q (new_AGEMA_signal_6780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4263 ( .C (clk), .D (new_AGEMA_signal_6783), .Q (new_AGEMA_signal_6784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4267 ( .C (clk), .D (new_AGEMA_signal_6787), .Q (new_AGEMA_signal_6788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4271 ( .C (clk), .D (new_AGEMA_signal_6791), .Q (new_AGEMA_signal_6792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4275 ( .C (clk), .D (new_AGEMA_signal_6795), .Q (new_AGEMA_signal_6796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4279 ( .C (clk), .D (new_AGEMA_signal_6799), .Q (new_AGEMA_signal_6800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4283 ( .C (clk), .D (new_AGEMA_signal_6803), .Q (new_AGEMA_signal_6804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4287 ( .C (clk), .D (new_AGEMA_signal_6807), .Q (new_AGEMA_signal_6808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4291 ( .C (clk), .D (new_AGEMA_signal_6811), .Q (new_AGEMA_signal_6812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4295 ( .C (clk), .D (new_AGEMA_signal_6815), .Q (new_AGEMA_signal_6816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4299 ( .C (clk), .D (new_AGEMA_signal_6819), .Q (new_AGEMA_signal_6820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4303 ( .C (clk), .D (new_AGEMA_signal_6823), .Q (new_AGEMA_signal_6824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4307 ( .C (clk), .D (new_AGEMA_signal_6827), .Q (new_AGEMA_signal_6828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4311 ( .C (clk), .D (new_AGEMA_signal_6831), .Q (new_AGEMA_signal_6832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4315 ( .C (clk), .D (new_AGEMA_signal_6835), .Q (new_AGEMA_signal_6836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4319 ( .C (clk), .D (new_AGEMA_signal_6839), .Q (new_AGEMA_signal_6840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4323 ( .C (clk), .D (new_AGEMA_signal_6843), .Q (new_AGEMA_signal_6844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4327 ( .C (clk), .D (new_AGEMA_signal_6847), .Q (new_AGEMA_signal_6848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4331 ( .C (clk), .D (new_AGEMA_signal_6851), .Q (new_AGEMA_signal_6852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4335 ( .C (clk), .D (new_AGEMA_signal_6855), .Q (new_AGEMA_signal_6856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4339 ( .C (clk), .D (new_AGEMA_signal_6859), .Q (new_AGEMA_signal_6860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4343 ( .C (clk), .D (new_AGEMA_signal_6863), .Q (new_AGEMA_signal_6864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4347 ( .C (clk), .D (new_AGEMA_signal_6867), .Q (new_AGEMA_signal_6868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4351 ( .C (clk), .D (new_AGEMA_signal_6871), .Q (new_AGEMA_signal_6872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4355 ( .C (clk), .D (new_AGEMA_signal_6875), .Q (new_AGEMA_signal_6876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4359 ( .C (clk), .D (new_AGEMA_signal_6879), .Q (new_AGEMA_signal_6880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4363 ( .C (clk), .D (new_AGEMA_signal_6883), .Q (new_AGEMA_signal_6884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4367 ( .C (clk), .D (new_AGEMA_signal_6887), .Q (new_AGEMA_signal_6888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4371 ( .C (clk), .D (new_AGEMA_signal_6891), .Q (new_AGEMA_signal_6892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4375 ( .C (clk), .D (new_AGEMA_signal_6895), .Q (new_AGEMA_signal_6896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4379 ( .C (clk), .D (new_AGEMA_signal_6899), .Q (new_AGEMA_signal_6900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4383 ( .C (clk), .D (new_AGEMA_signal_6903), .Q (new_AGEMA_signal_6904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4387 ( .C (clk), .D (new_AGEMA_signal_6907), .Q (new_AGEMA_signal_6908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4391 ( .C (clk), .D (new_AGEMA_signal_6911), .Q (new_AGEMA_signal_6912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4395 ( .C (clk), .D (new_AGEMA_signal_6915), .Q (new_AGEMA_signal_6916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4399 ( .C (clk), .D (new_AGEMA_signal_6919), .Q (new_AGEMA_signal_6920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4403 ( .C (clk), .D (new_AGEMA_signal_6923), .Q (new_AGEMA_signal_6924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4407 ( .C (clk), .D (new_AGEMA_signal_6927), .Q (new_AGEMA_signal_6928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4411 ( .C (clk), .D (new_AGEMA_signal_6931), .Q (new_AGEMA_signal_6932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4415 ( .C (clk), .D (new_AGEMA_signal_6935), .Q (new_AGEMA_signal_6936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4419 ( .C (clk), .D (new_AGEMA_signal_6939), .Q (new_AGEMA_signal_6940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4423 ( .C (clk), .D (new_AGEMA_signal_6943), .Q (new_AGEMA_signal_6944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4427 ( .C (clk), .D (new_AGEMA_signal_6947), .Q (new_AGEMA_signal_6948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4431 ( .C (clk), .D (new_AGEMA_signal_6951), .Q (new_AGEMA_signal_6952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4435 ( .C (clk), .D (new_AGEMA_signal_6955), .Q (new_AGEMA_signal_6956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4439 ( .C (clk), .D (new_AGEMA_signal_6959), .Q (new_AGEMA_signal_6960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4443 ( .C (clk), .D (new_AGEMA_signal_6963), .Q (new_AGEMA_signal_6964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4447 ( .C (clk), .D (new_AGEMA_signal_6967), .Q (new_AGEMA_signal_6968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4451 ( .C (clk), .D (new_AGEMA_signal_6971), .Q (new_AGEMA_signal_6972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4455 ( .C (clk), .D (new_AGEMA_signal_6975), .Q (new_AGEMA_signal_6976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4459 ( .C (clk), .D (new_AGEMA_signal_6979), .Q (new_AGEMA_signal_6980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4463 ( .C (clk), .D (new_AGEMA_signal_6983), .Q (new_AGEMA_signal_6984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4467 ( .C (clk), .D (new_AGEMA_signal_6987), .Q (new_AGEMA_signal_6988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4471 ( .C (clk), .D (new_AGEMA_signal_6991), .Q (new_AGEMA_signal_6992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4475 ( .C (clk), .D (new_AGEMA_signal_6995), .Q (new_AGEMA_signal_6996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4479 ( .C (clk), .D (new_AGEMA_signal_6999), .Q (new_AGEMA_signal_7000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4483 ( .C (clk), .D (new_AGEMA_signal_7003), .Q (new_AGEMA_signal_7004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4487 ( .C (clk), .D (new_AGEMA_signal_7007), .Q (new_AGEMA_signal_7008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4491 ( .C (clk), .D (new_AGEMA_signal_7011), .Q (new_AGEMA_signal_7012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4495 ( .C (clk), .D (new_AGEMA_signal_7015), .Q (new_AGEMA_signal_7016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4499 ( .C (clk), .D (new_AGEMA_signal_7019), .Q (new_AGEMA_signal_7020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4503 ( .C (clk), .D (new_AGEMA_signal_7023), .Q (new_AGEMA_signal_7024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4507 ( .C (clk), .D (new_AGEMA_signal_7027), .Q (new_AGEMA_signal_7028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4511 ( .C (clk), .D (new_AGEMA_signal_7031), .Q (new_AGEMA_signal_7032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4515 ( .C (clk), .D (new_AGEMA_signal_7035), .Q (new_AGEMA_signal_7036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4519 ( .C (clk), .D (new_AGEMA_signal_7039), .Q (new_AGEMA_signal_7040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4523 ( .C (clk), .D (new_AGEMA_signal_7043), .Q (new_AGEMA_signal_7044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4527 ( .C (clk), .D (new_AGEMA_signal_7047), .Q (new_AGEMA_signal_7048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4531 ( .C (clk), .D (new_AGEMA_signal_7051), .Q (new_AGEMA_signal_7052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4535 ( .C (clk), .D (new_AGEMA_signal_7055), .Q (new_AGEMA_signal_7056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4539 ( .C (clk), .D (new_AGEMA_signal_7059), .Q (new_AGEMA_signal_7060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4543 ( .C (clk), .D (new_AGEMA_signal_7063), .Q (new_AGEMA_signal_7064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4547 ( .C (clk), .D (new_AGEMA_signal_7067), .Q (new_AGEMA_signal_7068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4551 ( .C (clk), .D (new_AGEMA_signal_7071), .Q (new_AGEMA_signal_7072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4555 ( .C (clk), .D (new_AGEMA_signal_7075), .Q (new_AGEMA_signal_7076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4559 ( .C (clk), .D (new_AGEMA_signal_7079), .Q (new_AGEMA_signal_7080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4563 ( .C (clk), .D (new_AGEMA_signal_7083), .Q (new_AGEMA_signal_7084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4567 ( .C (clk), .D (new_AGEMA_signal_7087), .Q (new_AGEMA_signal_7088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4571 ( .C (clk), .D (new_AGEMA_signal_7091), .Q (new_AGEMA_signal_7092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4575 ( .C (clk), .D (new_AGEMA_signal_7095), .Q (new_AGEMA_signal_7096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4579 ( .C (clk), .D (new_AGEMA_signal_7099), .Q (new_AGEMA_signal_7100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4583 ( .C (clk), .D (new_AGEMA_signal_7103), .Q (new_AGEMA_signal_7104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4587 ( .C (clk), .D (new_AGEMA_signal_7107), .Q (new_AGEMA_signal_7108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4591 ( .C (clk), .D (new_AGEMA_signal_7111), .Q (new_AGEMA_signal_7112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4595 ( .C (clk), .D (new_AGEMA_signal_7115), .Q (new_AGEMA_signal_7116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4599 ( .C (clk), .D (new_AGEMA_signal_7119), .Q (new_AGEMA_signal_7120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4603 ( .C (clk), .D (new_AGEMA_signal_7123), .Q (new_AGEMA_signal_7124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4607 ( .C (clk), .D (new_AGEMA_signal_7127), .Q (new_AGEMA_signal_7128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4611 ( .C (clk), .D (new_AGEMA_signal_7131), .Q (new_AGEMA_signal_7132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4615 ( .C (clk), .D (new_AGEMA_signal_7135), .Q (new_AGEMA_signal_7136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4619 ( .C (clk), .D (new_AGEMA_signal_7139), .Q (new_AGEMA_signal_7140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4623 ( .C (clk), .D (new_AGEMA_signal_7143), .Q (new_AGEMA_signal_7144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4627 ( .C (clk), .D (new_AGEMA_signal_7147), .Q (new_AGEMA_signal_7148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4631 ( .C (clk), .D (new_AGEMA_signal_7151), .Q (new_AGEMA_signal_7152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4635 ( .C (clk), .D (new_AGEMA_signal_7155), .Q (new_AGEMA_signal_7156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4639 ( .C (clk), .D (new_AGEMA_signal_7159), .Q (new_AGEMA_signal_7160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4643 ( .C (clk), .D (new_AGEMA_signal_7163), .Q (new_AGEMA_signal_7164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4647 ( .C (clk), .D (new_AGEMA_signal_7167), .Q (new_AGEMA_signal_7168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4651 ( .C (clk), .D (new_AGEMA_signal_7171), .Q (new_AGEMA_signal_7172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4655 ( .C (clk), .D (new_AGEMA_signal_7175), .Q (new_AGEMA_signal_7176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4659 ( .C (clk), .D (new_AGEMA_signal_7179), .Q (new_AGEMA_signal_7180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4663 ( .C (clk), .D (new_AGEMA_signal_7183), .Q (new_AGEMA_signal_7184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4667 ( .C (clk), .D (new_AGEMA_signal_7187), .Q (new_AGEMA_signal_7188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4671 ( .C (clk), .D (new_AGEMA_signal_7191), .Q (new_AGEMA_signal_7192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4675 ( .C (clk), .D (new_AGEMA_signal_7195), .Q (new_AGEMA_signal_7196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4679 ( .C (clk), .D (new_AGEMA_signal_7199), .Q (new_AGEMA_signal_7200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4683 ( .C (clk), .D (new_AGEMA_signal_7203), .Q (new_AGEMA_signal_7204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4687 ( .C (clk), .D (new_AGEMA_signal_7207), .Q (new_AGEMA_signal_7208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4691 ( .C (clk), .D (new_AGEMA_signal_7211), .Q (new_AGEMA_signal_7212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4695 ( .C (clk), .D (new_AGEMA_signal_7215), .Q (new_AGEMA_signal_7216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4699 ( .C (clk), .D (new_AGEMA_signal_7219), .Q (new_AGEMA_signal_7220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4703 ( .C (clk), .D (new_AGEMA_signal_7223), .Q (new_AGEMA_signal_7224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4707 ( .C (clk), .D (new_AGEMA_signal_7227), .Q (new_AGEMA_signal_7228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4711 ( .C (clk), .D (new_AGEMA_signal_7231), .Q (new_AGEMA_signal_7232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4715 ( .C (clk), .D (new_AGEMA_signal_7235), .Q (new_AGEMA_signal_7236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4719 ( .C (clk), .D (new_AGEMA_signal_7239), .Q (new_AGEMA_signal_7240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4723 ( .C (clk), .D (new_AGEMA_signal_7243), .Q (new_AGEMA_signal_7244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4727 ( .C (clk), .D (new_AGEMA_signal_7247), .Q (new_AGEMA_signal_7248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4731 ( .C (clk), .D (new_AGEMA_signal_7251), .Q (new_AGEMA_signal_7252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4735 ( .C (clk), .D (new_AGEMA_signal_7255), .Q (new_AGEMA_signal_7256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4739 ( .C (clk), .D (new_AGEMA_signal_7259), .Q (new_AGEMA_signal_7260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4743 ( .C (clk), .D (new_AGEMA_signal_7263), .Q (new_AGEMA_signal_7264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4747 ( .C (clk), .D (new_AGEMA_signal_7267), .Q (new_AGEMA_signal_7268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4751 ( .C (clk), .D (new_AGEMA_signal_7271), .Q (new_AGEMA_signal_7272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4755 ( .C (clk), .D (new_AGEMA_signal_7275), .Q (new_AGEMA_signal_7276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4759 ( .C (clk), .D (new_AGEMA_signal_7279), .Q (new_AGEMA_signal_7280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4763 ( .C (clk), .D (new_AGEMA_signal_7283), .Q (new_AGEMA_signal_7284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4767 ( .C (clk), .D (new_AGEMA_signal_7287), .Q (new_AGEMA_signal_7288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4771 ( .C (clk), .D (new_AGEMA_signal_7291), .Q (new_AGEMA_signal_7292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4775 ( .C (clk), .D (new_AGEMA_signal_7295), .Q (new_AGEMA_signal_7296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4779 ( .C (clk), .D (new_AGEMA_signal_7299), .Q (new_AGEMA_signal_7300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4783 ( .C (clk), .D (new_AGEMA_signal_7303), .Q (new_AGEMA_signal_7304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4787 ( .C (clk), .D (new_AGEMA_signal_7307), .Q (new_AGEMA_signal_7308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4791 ( .C (clk), .D (new_AGEMA_signal_7311), .Q (new_AGEMA_signal_7312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4795 ( .C (clk), .D (new_AGEMA_signal_7315), .Q (new_AGEMA_signal_7316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4799 ( .C (clk), .D (new_AGEMA_signal_7319), .Q (new_AGEMA_signal_7320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4803 ( .C (clk), .D (new_AGEMA_signal_7323), .Q (new_AGEMA_signal_7324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4807 ( .C (clk), .D (new_AGEMA_signal_7327), .Q (new_AGEMA_signal_7328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4811 ( .C (clk), .D (new_AGEMA_signal_7331), .Q (new_AGEMA_signal_7332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4815 ( .C (clk), .D (new_AGEMA_signal_7335), .Q (new_AGEMA_signal_7336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4819 ( .C (clk), .D (new_AGEMA_signal_7339), .Q (new_AGEMA_signal_7340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4823 ( .C (clk), .D (new_AGEMA_signal_7343), .Q (new_AGEMA_signal_7344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4827 ( .C (clk), .D (new_AGEMA_signal_7347), .Q (new_AGEMA_signal_7348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4831 ( .C (clk), .D (new_AGEMA_signal_7351), .Q (new_AGEMA_signal_7352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4835 ( .C (clk), .D (new_AGEMA_signal_7355), .Q (new_AGEMA_signal_7356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4839 ( .C (clk), .D (new_AGEMA_signal_7359), .Q (new_AGEMA_signal_7360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4843 ( .C (clk), .D (new_AGEMA_signal_7363), .Q (new_AGEMA_signal_7364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4847 ( .C (clk), .D (new_AGEMA_signal_7367), .Q (new_AGEMA_signal_7368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4851 ( .C (clk), .D (new_AGEMA_signal_7371), .Q (new_AGEMA_signal_7372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4855 ( .C (clk), .D (new_AGEMA_signal_7375), .Q (new_AGEMA_signal_7376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4859 ( .C (clk), .D (new_AGEMA_signal_7379), .Q (new_AGEMA_signal_7380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4863 ( .C (clk), .D (new_AGEMA_signal_7383), .Q (new_AGEMA_signal_7384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4867 ( .C (clk), .D (new_AGEMA_signal_7387), .Q (new_AGEMA_signal_7388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4871 ( .C (clk), .D (new_AGEMA_signal_7391), .Q (new_AGEMA_signal_7392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4875 ( .C (clk), .D (new_AGEMA_signal_7395), .Q (new_AGEMA_signal_7396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4879 ( .C (clk), .D (new_AGEMA_signal_7399), .Q (new_AGEMA_signal_7400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4883 ( .C (clk), .D (new_AGEMA_signal_7403), .Q (new_AGEMA_signal_7404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4887 ( .C (clk), .D (new_AGEMA_signal_7407), .Q (new_AGEMA_signal_7408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4891 ( .C (clk), .D (new_AGEMA_signal_7411), .Q (new_AGEMA_signal_7412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4895 ( .C (clk), .D (new_AGEMA_signal_7415), .Q (new_AGEMA_signal_7416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4899 ( .C (clk), .D (new_AGEMA_signal_7419), .Q (new_AGEMA_signal_7420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4903 ( .C (clk), .D (new_AGEMA_signal_7423), .Q (new_AGEMA_signal_7424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4907 ( .C (clk), .D (new_AGEMA_signal_7427), .Q (new_AGEMA_signal_7428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4911 ( .C (clk), .D (new_AGEMA_signal_7431), .Q (new_AGEMA_signal_7432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4915 ( .C (clk), .D (new_AGEMA_signal_7435), .Q (new_AGEMA_signal_7436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4919 ( .C (clk), .D (new_AGEMA_signal_7439), .Q (new_AGEMA_signal_7440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4923 ( .C (clk), .D (new_AGEMA_signal_7443), .Q (new_AGEMA_signal_7444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4927 ( .C (clk), .D (new_AGEMA_signal_7447), .Q (new_AGEMA_signal_7448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4931 ( .C (clk), .D (new_AGEMA_signal_7451), .Q (new_AGEMA_signal_7452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4935 ( .C (clk), .D (new_AGEMA_signal_7455), .Q (new_AGEMA_signal_7456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4939 ( .C (clk), .D (new_AGEMA_signal_7459), .Q (new_AGEMA_signal_7460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4943 ( .C (clk), .D (new_AGEMA_signal_7463), .Q (new_AGEMA_signal_7464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4947 ( .C (clk), .D (new_AGEMA_signal_7467), .Q (new_AGEMA_signal_7468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4951 ( .C (clk), .D (new_AGEMA_signal_7471), .Q (new_AGEMA_signal_7472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4955 ( .C (clk), .D (new_AGEMA_signal_7475), .Q (new_AGEMA_signal_7476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4959 ( .C (clk), .D (new_AGEMA_signal_7479), .Q (new_AGEMA_signal_7480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4963 ( .C (clk), .D (new_AGEMA_signal_7483), .Q (new_AGEMA_signal_7484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4967 ( .C (clk), .D (new_AGEMA_signal_7487), .Q (new_AGEMA_signal_7488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4971 ( .C (clk), .D (new_AGEMA_signal_7491), .Q (new_AGEMA_signal_7492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4975 ( .C (clk), .D (new_AGEMA_signal_7495), .Q (new_AGEMA_signal_7496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4979 ( .C (clk), .D (new_AGEMA_signal_7499), .Q (new_AGEMA_signal_7500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4983 ( .C (clk), .D (new_AGEMA_signal_7503), .Q (new_AGEMA_signal_7504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4987 ( .C (clk), .D (new_AGEMA_signal_7507), .Q (new_AGEMA_signal_7508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4991 ( .C (clk), .D (new_AGEMA_signal_7511), .Q (new_AGEMA_signal_7512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4995 ( .C (clk), .D (new_AGEMA_signal_7515), .Q (new_AGEMA_signal_7516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4999 ( .C (clk), .D (new_AGEMA_signal_7519), .Q (new_AGEMA_signal_7520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5003 ( .C (clk), .D (new_AGEMA_signal_7523), .Q (new_AGEMA_signal_7524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5007 ( .C (clk), .D (new_AGEMA_signal_7527), .Q (new_AGEMA_signal_7528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5011 ( .C (clk), .D (new_AGEMA_signal_7531), .Q (new_AGEMA_signal_7532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5015 ( .C (clk), .D (new_AGEMA_signal_7535), .Q (new_AGEMA_signal_7536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5019 ( .C (clk), .D (new_AGEMA_signal_7539), .Q (new_AGEMA_signal_7540) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5023 ( .C (clk), .D (new_AGEMA_signal_7543), .Q (new_AGEMA_signal_7544) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5027 ( .C (clk), .D (new_AGEMA_signal_7547), .Q (new_AGEMA_signal_7548) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5031 ( .C (clk), .D (new_AGEMA_signal_7551), .Q (new_AGEMA_signal_7552) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5035 ( .C (clk), .D (new_AGEMA_signal_7555), .Q (new_AGEMA_signal_7556) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5039 ( .C (clk), .D (new_AGEMA_signal_7559), .Q (new_AGEMA_signal_7560) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5043 ( .C (clk), .D (new_AGEMA_signal_7563), .Q (new_AGEMA_signal_7564) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5047 ( .C (clk), .D (new_AGEMA_signal_7567), .Q (new_AGEMA_signal_7568) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5051 ( .C (clk), .D (new_AGEMA_signal_7571), .Q (new_AGEMA_signal_7572) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5055 ( .C (clk), .D (new_AGEMA_signal_7575), .Q (new_AGEMA_signal_7576) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5059 ( .C (clk), .D (new_AGEMA_signal_7579), .Q (new_AGEMA_signal_7580) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5063 ( .C (clk), .D (new_AGEMA_signal_7583), .Q (new_AGEMA_signal_7584) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5067 ( .C (clk), .D (new_AGEMA_signal_7587), .Q (new_AGEMA_signal_7588) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5071 ( .C (clk), .D (new_AGEMA_signal_7591), .Q (new_AGEMA_signal_7592) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5075 ( .C (clk), .D (new_AGEMA_signal_7595), .Q (new_AGEMA_signal_7596) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5079 ( .C (clk), .D (new_AGEMA_signal_7599), .Q (new_AGEMA_signal_7600) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5083 ( .C (clk), .D (new_AGEMA_signal_7603), .Q (new_AGEMA_signal_7604) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5087 ( .C (clk), .D (new_AGEMA_signal_7607), .Q (new_AGEMA_signal_7608) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5091 ( .C (clk), .D (new_AGEMA_signal_7611), .Q (new_AGEMA_signal_7612) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5095 ( .C (clk), .D (new_AGEMA_signal_7615), .Q (new_AGEMA_signal_7616) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5099 ( .C (clk), .D (new_AGEMA_signal_7619), .Q (new_AGEMA_signal_7620) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5103 ( .C (clk), .D (new_AGEMA_signal_7623), .Q (new_AGEMA_signal_7624) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5107 ( .C (clk), .D (new_AGEMA_signal_7627), .Q (new_AGEMA_signal_7628) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5111 ( .C (clk), .D (new_AGEMA_signal_7631), .Q (new_AGEMA_signal_7632) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5115 ( .C (clk), .D (new_AGEMA_signal_7635), .Q (new_AGEMA_signal_7636) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5119 ( .C (clk), .D (new_AGEMA_signal_7639), .Q (new_AGEMA_signal_7640) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5123 ( .C (clk), .D (new_AGEMA_signal_7643), .Q (new_AGEMA_signal_7644) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5127 ( .C (clk), .D (new_AGEMA_signal_7647), .Q (new_AGEMA_signal_7648) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5131 ( .C (clk), .D (new_AGEMA_signal_7651), .Q (new_AGEMA_signal_7652) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5135 ( .C (clk), .D (new_AGEMA_signal_7655), .Q (new_AGEMA_signal_7656) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5139 ( .C (clk), .D (new_AGEMA_signal_7659), .Q (new_AGEMA_signal_7660) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5143 ( .C (clk), .D (new_AGEMA_signal_7663), .Q (new_AGEMA_signal_7664) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5147 ( .C (clk), .D (new_AGEMA_signal_7667), .Q (new_AGEMA_signal_7668) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5151 ( .C (clk), .D (new_AGEMA_signal_7671), .Q (new_AGEMA_signal_7672) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5155 ( .C (clk), .D (new_AGEMA_signal_7675), .Q (new_AGEMA_signal_7676) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5159 ( .C (clk), .D (new_AGEMA_signal_7679), .Q (new_AGEMA_signal_7680) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5163 ( .C (clk), .D (new_AGEMA_signal_7683), .Q (new_AGEMA_signal_7684) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5167 ( .C (clk), .D (new_AGEMA_signal_7687), .Q (new_AGEMA_signal_7688) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5171 ( .C (clk), .D (new_AGEMA_signal_7691), .Q (new_AGEMA_signal_7692) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5175 ( .C (clk), .D (new_AGEMA_signal_7695), .Q (new_AGEMA_signal_7696) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5179 ( .C (clk), .D (new_AGEMA_signal_7699), .Q (new_AGEMA_signal_7700) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5183 ( .C (clk), .D (new_AGEMA_signal_7703), .Q (new_AGEMA_signal_7704) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5187 ( .C (clk), .D (new_AGEMA_signal_7707), .Q (new_AGEMA_signal_7708) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5191 ( .C (clk), .D (new_AGEMA_signal_7711), .Q (new_AGEMA_signal_7712) ) ;
    buf_clk new_AGEMA_reg_buffer_5195 ( .C (clk), .D (new_AGEMA_signal_7715), .Q (new_AGEMA_signal_7716) ) ;
    buf_clk new_AGEMA_reg_buffer_5199 ( .C (clk), .D (new_AGEMA_signal_7719), .Q (new_AGEMA_signal_7720) ) ;
    buf_clk new_AGEMA_reg_buffer_5203 ( .C (clk), .D (new_AGEMA_signal_7723), .Q (new_AGEMA_signal_7724) ) ;
    buf_clk new_AGEMA_reg_buffer_5207 ( .C (clk), .D (new_AGEMA_signal_7727), .Q (new_AGEMA_signal_7728) ) ;
    buf_clk new_AGEMA_reg_buffer_5211 ( .C (clk), .D (new_AGEMA_signal_7731), .Q (new_AGEMA_signal_7732) ) ;
    buf_clk new_AGEMA_reg_buffer_5215 ( .C (clk), .D (new_AGEMA_signal_7735), .Q (new_AGEMA_signal_7736) ) ;
    buf_clk new_AGEMA_reg_buffer_5219 ( .C (clk), .D (new_AGEMA_signal_7739), .Q (new_AGEMA_signal_7740) ) ;
    buf_clk new_AGEMA_reg_buffer_5223 ( .C (clk), .D (new_AGEMA_signal_7743), .Q (new_AGEMA_signal_7744) ) ;
    buf_clk new_AGEMA_reg_buffer_5227 ( .C (clk), .D (new_AGEMA_signal_7747), .Q (new_AGEMA_signal_7748) ) ;
    buf_clk new_AGEMA_reg_buffer_5231 ( .C (clk), .D (new_AGEMA_signal_7751), .Q (new_AGEMA_signal_7752) ) ;
    buf_clk new_AGEMA_reg_buffer_5235 ( .C (clk), .D (new_AGEMA_signal_7755), .Q (new_AGEMA_signal_7756) ) ;
    buf_clk new_AGEMA_reg_buffer_5239 ( .C (clk), .D (new_AGEMA_signal_7759), .Q (new_AGEMA_signal_7760) ) ;
    buf_clk new_AGEMA_reg_buffer_5243 ( .C (clk), .D (new_AGEMA_signal_7763), .Q (new_AGEMA_signal_7764) ) ;
    buf_clk new_AGEMA_reg_buffer_5247 ( .C (clk), .D (new_AGEMA_signal_7767), .Q (new_AGEMA_signal_7768) ) ;
    buf_clk new_AGEMA_reg_buffer_5251 ( .C (clk), .D (new_AGEMA_signal_7771), .Q (new_AGEMA_signal_7772) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5255 ( .C (clk), .D (new_AGEMA_signal_7775), .Q (new_AGEMA_signal_7776) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5259 ( .C (clk), .D (new_AGEMA_signal_7779), .Q (new_AGEMA_signal_7780) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5263 ( .C (clk), .D (new_AGEMA_signal_7783), .Q (new_AGEMA_signal_7784) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5267 ( .C (clk), .D (new_AGEMA_signal_7787), .Q (new_AGEMA_signal_7788) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5271 ( .C (clk), .D (new_AGEMA_signal_7791), .Q (new_AGEMA_signal_7792) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5275 ( .C (clk), .D (new_AGEMA_signal_7795), .Q (new_AGEMA_signal_7796) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5279 ( .C (clk), .D (new_AGEMA_signal_7799), .Q (new_AGEMA_signal_7800) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5283 ( .C (clk), .D (new_AGEMA_signal_7803), .Q (new_AGEMA_signal_7804) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5287 ( .C (clk), .D (new_AGEMA_signal_7807), .Q (new_AGEMA_signal_7808) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5291 ( .C (clk), .D (new_AGEMA_signal_7811), .Q (new_AGEMA_signal_7812) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5295 ( .C (clk), .D (new_AGEMA_signal_7815), .Q (new_AGEMA_signal_7816) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5299 ( .C (clk), .D (new_AGEMA_signal_7819), .Q (new_AGEMA_signal_7820) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5303 ( .C (clk), .D (new_AGEMA_signal_7823), .Q (new_AGEMA_signal_7824) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5307 ( .C (clk), .D (new_AGEMA_signal_7827), .Q (new_AGEMA_signal_7828) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5311 ( .C (clk), .D (new_AGEMA_signal_7831), .Q (new_AGEMA_signal_7832) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5315 ( .C (clk), .D (new_AGEMA_signal_7835), .Q (new_AGEMA_signal_7836) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5319 ( .C (clk), .D (new_AGEMA_signal_7839), .Q (new_AGEMA_signal_7840) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5323 ( .C (clk), .D (new_AGEMA_signal_7843), .Q (new_AGEMA_signal_7844) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5327 ( .C (clk), .D (new_AGEMA_signal_7847), .Q (new_AGEMA_signal_7848) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5331 ( .C (clk), .D (new_AGEMA_signal_7851), .Q (new_AGEMA_signal_7852) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5335 ( .C (clk), .D (new_AGEMA_signal_7855), .Q (new_AGEMA_signal_7856) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5339 ( .C (clk), .D (new_AGEMA_signal_7859), .Q (new_AGEMA_signal_7860) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5343 ( .C (clk), .D (new_AGEMA_signal_7863), .Q (new_AGEMA_signal_7864) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5347 ( .C (clk), .D (new_AGEMA_signal_7867), .Q (new_AGEMA_signal_7868) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5351 ( .C (clk), .D (new_AGEMA_signal_7871), .Q (new_AGEMA_signal_7872) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5355 ( .C (clk), .D (new_AGEMA_signal_7875), .Q (new_AGEMA_signal_7876) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5359 ( .C (clk), .D (new_AGEMA_signal_7879), .Q (new_AGEMA_signal_7880) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5363 ( .C (clk), .D (new_AGEMA_signal_7883), .Q (new_AGEMA_signal_7884) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5367 ( .C (clk), .D (new_AGEMA_signal_7887), .Q (new_AGEMA_signal_7888) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5371 ( .C (clk), .D (new_AGEMA_signal_7891), .Q (new_AGEMA_signal_7892) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5375 ( .C (clk), .D (new_AGEMA_signal_7895), .Q (new_AGEMA_signal_7896) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5379 ( .C (clk), .D (new_AGEMA_signal_7899), .Q (new_AGEMA_signal_7900) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5383 ( .C (clk), .D (new_AGEMA_signal_7903), .Q (new_AGEMA_signal_7904) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5387 ( .C (clk), .D (new_AGEMA_signal_7907), .Q (new_AGEMA_signal_7908) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5391 ( .C (clk), .D (new_AGEMA_signal_7911), .Q (new_AGEMA_signal_7912) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5395 ( .C (clk), .D (new_AGEMA_signal_7915), .Q (new_AGEMA_signal_7916) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5399 ( .C (clk), .D (new_AGEMA_signal_7919), .Q (new_AGEMA_signal_7920) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5403 ( .C (clk), .D (new_AGEMA_signal_7923), .Q (new_AGEMA_signal_7924) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5407 ( .C (clk), .D (new_AGEMA_signal_7927), .Q (new_AGEMA_signal_7928) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5411 ( .C (clk), .D (new_AGEMA_signal_7931), .Q (new_AGEMA_signal_7932) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5415 ( .C (clk), .D (new_AGEMA_signal_7935), .Q (new_AGEMA_signal_7936) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5419 ( .C (clk), .D (new_AGEMA_signal_7939), .Q (new_AGEMA_signal_7940) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5423 ( .C (clk), .D (new_AGEMA_signal_7943), .Q (new_AGEMA_signal_7944) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5427 ( .C (clk), .D (new_AGEMA_signal_7947), .Q (new_AGEMA_signal_7948) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5431 ( .C (clk), .D (new_AGEMA_signal_7951), .Q (new_AGEMA_signal_7952) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5435 ( .C (clk), .D (new_AGEMA_signal_7955), .Q (new_AGEMA_signal_7956) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5439 ( .C (clk), .D (new_AGEMA_signal_7959), .Q (new_AGEMA_signal_7960) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5443 ( .C (clk), .D (new_AGEMA_signal_7963), .Q (new_AGEMA_signal_7964) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5447 ( .C (clk), .D (new_AGEMA_signal_7967), .Q (new_AGEMA_signal_7968) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5451 ( .C (clk), .D (new_AGEMA_signal_7971), .Q (new_AGEMA_signal_7972) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5455 ( .C (clk), .D (new_AGEMA_signal_7975), .Q (new_AGEMA_signal_7976) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5459 ( .C (clk), .D (new_AGEMA_signal_7979), .Q (new_AGEMA_signal_7980) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5463 ( .C (clk), .D (new_AGEMA_signal_7983), .Q (new_AGEMA_signal_7984) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5467 ( .C (clk), .D (new_AGEMA_signal_7987), .Q (new_AGEMA_signal_7988) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5471 ( .C (clk), .D (new_AGEMA_signal_7991), .Q (new_AGEMA_signal_7992) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5475 ( .C (clk), .D (new_AGEMA_signal_7995), .Q (new_AGEMA_signal_7996) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5479 ( .C (clk), .D (new_AGEMA_signal_7999), .Q (new_AGEMA_signal_8000) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5483 ( .C (clk), .D (new_AGEMA_signal_8003), .Q (new_AGEMA_signal_8004) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5487 ( .C (clk), .D (new_AGEMA_signal_8007), .Q (new_AGEMA_signal_8008) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5491 ( .C (clk), .D (new_AGEMA_signal_8011), .Q (new_AGEMA_signal_8012) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5495 ( .C (clk), .D (new_AGEMA_signal_8015), .Q (new_AGEMA_signal_8016) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5499 ( .C (clk), .D (new_AGEMA_signal_8019), .Q (new_AGEMA_signal_8020) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5503 ( .C (clk), .D (new_AGEMA_signal_8023), .Q (new_AGEMA_signal_8024) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5507 ( .C (clk), .D (new_AGEMA_signal_8027), .Q (new_AGEMA_signal_8028) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5511 ( .C (clk), .D (new_AGEMA_signal_8031), .Q (new_AGEMA_signal_8032) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5515 ( .C (clk), .D (new_AGEMA_signal_8035), .Q (new_AGEMA_signal_8036) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5519 ( .C (clk), .D (new_AGEMA_signal_8039), .Q (new_AGEMA_signal_8040) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5523 ( .C (clk), .D (new_AGEMA_signal_8043), .Q (new_AGEMA_signal_8044) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5527 ( .C (clk), .D (new_AGEMA_signal_8047), .Q (new_AGEMA_signal_8048) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5531 ( .C (clk), .D (new_AGEMA_signal_8051), .Q (new_AGEMA_signal_8052) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5535 ( .C (clk), .D (new_AGEMA_signal_8055), .Q (new_AGEMA_signal_8056) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5539 ( .C (clk), .D (new_AGEMA_signal_8059), .Q (new_AGEMA_signal_8060) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5543 ( .C (clk), .D (new_AGEMA_signal_8063), .Q (new_AGEMA_signal_8064) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5547 ( .C (clk), .D (new_AGEMA_signal_8067), .Q (new_AGEMA_signal_8068) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5551 ( .C (clk), .D (new_AGEMA_signal_8071), .Q (new_AGEMA_signal_8072) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5555 ( .C (clk), .D (new_AGEMA_signal_8075), .Q (new_AGEMA_signal_8076) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5559 ( .C (clk), .D (new_AGEMA_signal_8079), .Q (new_AGEMA_signal_8080) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5563 ( .C (clk), .D (new_AGEMA_signal_8083), .Q (new_AGEMA_signal_8084) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5567 ( .C (clk), .D (new_AGEMA_signal_8087), .Q (new_AGEMA_signal_8088) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5571 ( .C (clk), .D (new_AGEMA_signal_8091), .Q (new_AGEMA_signal_8092) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5575 ( .C (clk), .D (new_AGEMA_signal_8095), .Q (new_AGEMA_signal_8096) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5579 ( .C (clk), .D (new_AGEMA_signal_8099), .Q (new_AGEMA_signal_8100) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5583 ( .C (clk), .D (new_AGEMA_signal_8103), .Q (new_AGEMA_signal_8104) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5587 ( .C (clk), .D (new_AGEMA_signal_8107), .Q (new_AGEMA_signal_8108) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5591 ( .C (clk), .D (new_AGEMA_signal_8111), .Q (new_AGEMA_signal_8112) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5595 ( .C (clk), .D (new_AGEMA_signal_8115), .Q (new_AGEMA_signal_8116) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5599 ( .C (clk), .D (new_AGEMA_signal_8119), .Q (new_AGEMA_signal_8120) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5603 ( .C (clk), .D (new_AGEMA_signal_8123), .Q (new_AGEMA_signal_8124) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5607 ( .C (clk), .D (new_AGEMA_signal_8127), .Q (new_AGEMA_signal_8128) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5611 ( .C (clk), .D (new_AGEMA_signal_8131), .Q (new_AGEMA_signal_8132) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5615 ( .C (clk), .D (new_AGEMA_signal_8135), .Q (new_AGEMA_signal_8136) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5619 ( .C (clk), .D (new_AGEMA_signal_8139), .Q (new_AGEMA_signal_8140) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5623 ( .C (clk), .D (new_AGEMA_signal_8143), .Q (new_AGEMA_signal_8144) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5627 ( .C (clk), .D (new_AGEMA_signal_8147), .Q (new_AGEMA_signal_8148) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5631 ( .C (clk), .D (new_AGEMA_signal_8151), .Q (new_AGEMA_signal_8152) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5635 ( .C (clk), .D (new_AGEMA_signal_8155), .Q (new_AGEMA_signal_8156) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5639 ( .C (clk), .D (new_AGEMA_signal_8159), .Q (new_AGEMA_signal_8160) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5643 ( .C (clk), .D (new_AGEMA_signal_8163), .Q (new_AGEMA_signal_8164) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5647 ( .C (clk), .D (new_AGEMA_signal_8167), .Q (new_AGEMA_signal_8168) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5651 ( .C (clk), .D (new_AGEMA_signal_8171), .Q (new_AGEMA_signal_8172) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5655 ( .C (clk), .D (new_AGEMA_signal_8175), .Q (new_AGEMA_signal_8176) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5659 ( .C (clk), .D (new_AGEMA_signal_8179), .Q (new_AGEMA_signal_8180) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5663 ( .C (clk), .D (new_AGEMA_signal_8183), .Q (new_AGEMA_signal_8184) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5667 ( .C (clk), .D (new_AGEMA_signal_8187), .Q (new_AGEMA_signal_8188) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5671 ( .C (clk), .D (new_AGEMA_signal_8191), .Q (new_AGEMA_signal_8192) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5675 ( .C (clk), .D (new_AGEMA_signal_8195), .Q (new_AGEMA_signal_8196) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5679 ( .C (clk), .D (new_AGEMA_signal_8199), .Q (new_AGEMA_signal_8200) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5683 ( .C (clk), .D (new_AGEMA_signal_8203), .Q (new_AGEMA_signal_8204) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5687 ( .C (clk), .D (new_AGEMA_signal_8207), .Q (new_AGEMA_signal_8208) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5691 ( .C (clk), .D (new_AGEMA_signal_8211), .Q (new_AGEMA_signal_8212) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5695 ( .C (clk), .D (new_AGEMA_signal_8215), .Q (new_AGEMA_signal_8216) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5699 ( .C (clk), .D (new_AGEMA_signal_8219), .Q (new_AGEMA_signal_8220) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5703 ( .C (clk), .D (new_AGEMA_signal_8223), .Q (new_AGEMA_signal_8224) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5707 ( .C (clk), .D (new_AGEMA_signal_8227), .Q (new_AGEMA_signal_8228) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5711 ( .C (clk), .D (new_AGEMA_signal_8231), .Q (new_AGEMA_signal_8232) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5715 ( .C (clk), .D (new_AGEMA_signal_8235), .Q (new_AGEMA_signal_8236) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5719 ( .C (clk), .D (new_AGEMA_signal_8239), .Q (new_AGEMA_signal_8240) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5723 ( .C (clk), .D (new_AGEMA_signal_8243), .Q (new_AGEMA_signal_8244) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5727 ( .C (clk), .D (new_AGEMA_signal_8247), .Q (new_AGEMA_signal_8248) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5731 ( .C (clk), .D (new_AGEMA_signal_8251), .Q (new_AGEMA_signal_8252) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5735 ( .C (clk), .D (new_AGEMA_signal_8255), .Q (new_AGEMA_signal_8256) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5739 ( .C (clk), .D (new_AGEMA_signal_8259), .Q (new_AGEMA_signal_8260) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5743 ( .C (clk), .D (new_AGEMA_signal_8263), .Q (new_AGEMA_signal_8264) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5747 ( .C (clk), .D (new_AGEMA_signal_8267), .Q (new_AGEMA_signal_8268) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5751 ( .C (clk), .D (new_AGEMA_signal_8271), .Q (new_AGEMA_signal_8272) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5755 ( .C (clk), .D (new_AGEMA_signal_8275), .Q (new_AGEMA_signal_8276) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5759 ( .C (clk), .D (new_AGEMA_signal_8279), .Q (new_AGEMA_signal_8280) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5763 ( .C (clk), .D (new_AGEMA_signal_8283), .Q (new_AGEMA_signal_8284) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5767 ( .C (clk), .D (new_AGEMA_signal_8287), .Q (new_AGEMA_signal_8288) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5771 ( .C (clk), .D (new_AGEMA_signal_8291), .Q (new_AGEMA_signal_8292) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5775 ( .C (clk), .D (new_AGEMA_signal_8295), .Q (new_AGEMA_signal_8296) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5779 ( .C (clk), .D (new_AGEMA_signal_8299), .Q (new_AGEMA_signal_8300) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5783 ( .C (clk), .D (new_AGEMA_signal_8303), .Q (new_AGEMA_signal_8304) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5787 ( .C (clk), .D (new_AGEMA_signal_8307), .Q (new_AGEMA_signal_8308) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5791 ( .C (clk), .D (new_AGEMA_signal_8311), .Q (new_AGEMA_signal_8312) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5795 ( .C (clk), .D (new_AGEMA_signal_8315), .Q (new_AGEMA_signal_8316) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5799 ( .C (clk), .D (new_AGEMA_signal_8319), .Q (new_AGEMA_signal_8320) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5803 ( .C (clk), .D (new_AGEMA_signal_8323), .Q (new_AGEMA_signal_8324) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5807 ( .C (clk), .D (new_AGEMA_signal_8327), .Q (new_AGEMA_signal_8328) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5811 ( .C (clk), .D (new_AGEMA_signal_8331), .Q (new_AGEMA_signal_8332) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5815 ( .C (clk), .D (new_AGEMA_signal_8335), .Q (new_AGEMA_signal_8336) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5819 ( .C (clk), .D (new_AGEMA_signal_8339), .Q (new_AGEMA_signal_8340) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5823 ( .C (clk), .D (new_AGEMA_signal_8343), .Q (new_AGEMA_signal_8344) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5827 ( .C (clk), .D (new_AGEMA_signal_8347), .Q (new_AGEMA_signal_8348) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5831 ( .C (clk), .D (new_AGEMA_signal_8351), .Q (new_AGEMA_signal_8352) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5835 ( .C (clk), .D (new_AGEMA_signal_8355), .Q (new_AGEMA_signal_8356) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5839 ( .C (clk), .D (new_AGEMA_signal_8359), .Q (new_AGEMA_signal_8360) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5843 ( .C (clk), .D (new_AGEMA_signal_8363), .Q (new_AGEMA_signal_8364) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5847 ( .C (clk), .D (new_AGEMA_signal_8367), .Q (new_AGEMA_signal_8368) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5851 ( .C (clk), .D (new_AGEMA_signal_8371), .Q (new_AGEMA_signal_8372) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5855 ( .C (clk), .D (new_AGEMA_signal_8375), .Q (new_AGEMA_signal_8376) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5859 ( .C (clk), .D (new_AGEMA_signal_8379), .Q (new_AGEMA_signal_8380) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5863 ( .C (clk), .D (new_AGEMA_signal_8383), .Q (new_AGEMA_signal_8384) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5867 ( .C (clk), .D (new_AGEMA_signal_8387), .Q (new_AGEMA_signal_8388) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5871 ( .C (clk), .D (new_AGEMA_signal_8391), .Q (new_AGEMA_signal_8392) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5875 ( .C (clk), .D (new_AGEMA_signal_8395), .Q (new_AGEMA_signal_8396) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5879 ( .C (clk), .D (new_AGEMA_signal_8399), .Q (new_AGEMA_signal_8400) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5883 ( .C (clk), .D (new_AGEMA_signal_8403), .Q (new_AGEMA_signal_8404) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5887 ( .C (clk), .D (new_AGEMA_signal_8407), .Q (new_AGEMA_signal_8408) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5891 ( .C (clk), .D (new_AGEMA_signal_8411), .Q (new_AGEMA_signal_8412) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5895 ( .C (clk), .D (new_AGEMA_signal_8415), .Q (new_AGEMA_signal_8416) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5899 ( .C (clk), .D (new_AGEMA_signal_8419), .Q (new_AGEMA_signal_8420) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5903 ( .C (clk), .D (new_AGEMA_signal_8423), .Q (new_AGEMA_signal_8424) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5907 ( .C (clk), .D (new_AGEMA_signal_8427), .Q (new_AGEMA_signal_8428) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5911 ( .C (clk), .D (new_AGEMA_signal_8431), .Q (new_AGEMA_signal_8432) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5915 ( .C (clk), .D (new_AGEMA_signal_8435), .Q (new_AGEMA_signal_8436) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5919 ( .C (clk), .D (new_AGEMA_signal_8439), .Q (new_AGEMA_signal_8440) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5923 ( .C (clk), .D (new_AGEMA_signal_8443), .Q (new_AGEMA_signal_8444) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5927 ( .C (clk), .D (new_AGEMA_signal_8447), .Q (new_AGEMA_signal_8448) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5931 ( .C (clk), .D (new_AGEMA_signal_8451), .Q (new_AGEMA_signal_8452) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5935 ( .C (clk), .D (new_AGEMA_signal_8455), .Q (new_AGEMA_signal_8456) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5939 ( .C (clk), .D (new_AGEMA_signal_8459), .Q (new_AGEMA_signal_8460) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5943 ( .C (clk), .D (new_AGEMA_signal_8463), .Q (new_AGEMA_signal_8464) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5947 ( .C (clk), .D (new_AGEMA_signal_8467), .Q (new_AGEMA_signal_8468) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5951 ( .C (clk), .D (new_AGEMA_signal_8471), .Q (new_AGEMA_signal_8472) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5955 ( .C (clk), .D (new_AGEMA_signal_8475), .Q (new_AGEMA_signal_8476) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5959 ( .C (clk), .D (new_AGEMA_signal_8479), .Q (new_AGEMA_signal_8480) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5963 ( .C (clk), .D (new_AGEMA_signal_8483), .Q (new_AGEMA_signal_8484) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5967 ( .C (clk), .D (new_AGEMA_signal_8487), .Q (new_AGEMA_signal_8488) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5971 ( .C (clk), .D (new_AGEMA_signal_8491), .Q (new_AGEMA_signal_8492) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5975 ( .C (clk), .D (new_AGEMA_signal_8495), .Q (new_AGEMA_signal_8496) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5979 ( .C (clk), .D (new_AGEMA_signal_8499), .Q (new_AGEMA_signal_8500) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5983 ( .C (clk), .D (new_AGEMA_signal_8503), .Q (new_AGEMA_signal_8504) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5987 ( .C (clk), .D (new_AGEMA_signal_8507), .Q (new_AGEMA_signal_8508) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5991 ( .C (clk), .D (new_AGEMA_signal_8511), .Q (new_AGEMA_signal_8512) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5995 ( .C (clk), .D (new_AGEMA_signal_8515), .Q (new_AGEMA_signal_8516) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5999 ( .C (clk), .D (new_AGEMA_signal_8519), .Q (new_AGEMA_signal_8520) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6003 ( .C (clk), .D (new_AGEMA_signal_8523), .Q (new_AGEMA_signal_8524) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6007 ( .C (clk), .D (new_AGEMA_signal_8527), .Q (new_AGEMA_signal_8528) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6011 ( .C (clk), .D (new_AGEMA_signal_8531), .Q (new_AGEMA_signal_8532) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6015 ( .C (clk), .D (new_AGEMA_signal_8535), .Q (new_AGEMA_signal_8536) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6019 ( .C (clk), .D (new_AGEMA_signal_8539), .Q (new_AGEMA_signal_8540) ) ;
    buf_clk new_AGEMA_reg_buffer_6023 ( .C (clk), .D (new_AGEMA_signal_8543), .Q (new_AGEMA_signal_8544) ) ;
    buf_clk new_AGEMA_reg_buffer_6027 ( .C (clk), .D (new_AGEMA_signal_8547), .Q (new_AGEMA_signal_8548) ) ;
    buf_clk new_AGEMA_reg_buffer_6031 ( .C (clk), .D (new_AGEMA_signal_8551), .Q (new_AGEMA_signal_8552) ) ;
    buf_clk new_AGEMA_reg_buffer_6035 ( .C (clk), .D (new_AGEMA_signal_8555), .Q (new_AGEMA_signal_8556) ) ;
    buf_clk new_AGEMA_reg_buffer_6039 ( .C (clk), .D (new_AGEMA_signal_8559), .Q (new_AGEMA_signal_8560) ) ;
    buf_clk new_AGEMA_reg_buffer_6043 ( .C (clk), .D (new_AGEMA_signal_8563), .Q (new_AGEMA_signal_8564) ) ;
    buf_clk new_AGEMA_reg_buffer_6047 ( .C (clk), .D (new_AGEMA_signal_8567), .Q (new_AGEMA_signal_8568) ) ;

    /* cells in depth 4 */
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4035, RoundOutput[0]}), .a ({new_AGEMA_signal_4689, new_AGEMA_signal_4685}), .c ({new_AGEMA_signal_4156, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4195, RoundOutput[1]}), .a ({new_AGEMA_signal_4697, new_AGEMA_signal_4693}), .c ({new_AGEMA_signal_4273, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4036, RoundOutput[2]}), .a ({new_AGEMA_signal_4705, new_AGEMA_signal_4701}), .c ({new_AGEMA_signal_4158, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4196, RoundOutput[3]}), .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4709}), .c ({new_AGEMA_signal_4275, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4197, RoundOutput[4]}), .a ({new_AGEMA_signal_4721, new_AGEMA_signal_4717}), .c ({new_AGEMA_signal_4277, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4037, RoundOutput[5]}), .a ({new_AGEMA_signal_4729, new_AGEMA_signal_4725}), .c ({new_AGEMA_signal_4160, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4038, RoundOutput[6]}), .a ({new_AGEMA_signal_4737, new_AGEMA_signal_4733}), .c ({new_AGEMA_signal_4162, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4039, RoundOutput[7]}), .a ({new_AGEMA_signal_4745, new_AGEMA_signal_4741}), .c ({new_AGEMA_signal_4164, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4040, RoundOutput[8]}), .a ({new_AGEMA_signal_4753, new_AGEMA_signal_4749}), .c ({new_AGEMA_signal_4166, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4198, RoundOutput[9]}), .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4757}), .c ({new_AGEMA_signal_4279, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4041, RoundOutput[10]}), .a ({new_AGEMA_signal_4769, new_AGEMA_signal_4765}), .c ({new_AGEMA_signal_4168, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4199, RoundOutput[11]}), .a ({new_AGEMA_signal_4777, new_AGEMA_signal_4773}), .c ({new_AGEMA_signal_4281, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4200, RoundOutput[12]}), .a ({new_AGEMA_signal_4785, new_AGEMA_signal_4781}), .c ({new_AGEMA_signal_4283, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4042, RoundOutput[13]}), .a ({new_AGEMA_signal_4793, new_AGEMA_signal_4789}), .c ({new_AGEMA_signal_4170, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4043, RoundOutput[14]}), .a ({new_AGEMA_signal_4801, new_AGEMA_signal_4797}), .c ({new_AGEMA_signal_4172, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4044, RoundOutput[15]}), .a ({new_AGEMA_signal_4809, new_AGEMA_signal_4805}), .c ({new_AGEMA_signal_4174, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4045, RoundOutput[16]}), .a ({new_AGEMA_signal_4817, new_AGEMA_signal_4813}), .c ({new_AGEMA_signal_4176, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4201, RoundOutput[17]}), .a ({new_AGEMA_signal_4825, new_AGEMA_signal_4821}), .c ({new_AGEMA_signal_4285, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4046, RoundOutput[18]}), .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4829}), .c ({new_AGEMA_signal_4178, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4202, RoundOutput[19]}), .a ({new_AGEMA_signal_4841, new_AGEMA_signal_4837}), .c ({new_AGEMA_signal_4287, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4203, RoundOutput[20]}), .a ({new_AGEMA_signal_4849, new_AGEMA_signal_4845}), .c ({new_AGEMA_signal_4289, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4047, RoundOutput[21]}), .a ({new_AGEMA_signal_4857, new_AGEMA_signal_4853}), .c ({new_AGEMA_signal_4180, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4048, RoundOutput[22]}), .a ({new_AGEMA_signal_4865, new_AGEMA_signal_4861}), .c ({new_AGEMA_signal_4182, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4049, RoundOutput[23]}), .a ({new_AGEMA_signal_4873, new_AGEMA_signal_4869}), .c ({new_AGEMA_signal_4184, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4050, RoundOutput[24]}), .a ({new_AGEMA_signal_4881, new_AGEMA_signal_4877}), .c ({new_AGEMA_signal_4186, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4204, RoundOutput[25]}), .a ({new_AGEMA_signal_4889, new_AGEMA_signal_4885}), .c ({new_AGEMA_signal_4291, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4051, RoundOutput[26]}), .a ({new_AGEMA_signal_4897, new_AGEMA_signal_4893}), .c ({new_AGEMA_signal_4188, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4205, RoundOutput[27]}), .a ({new_AGEMA_signal_4905, new_AGEMA_signal_4901}), .c ({new_AGEMA_signal_4293, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4206, RoundOutput[28]}), .a ({new_AGEMA_signal_4913, new_AGEMA_signal_4909}), .c ({new_AGEMA_signal_4295, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4052, RoundOutput[29]}), .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4917}), .c ({new_AGEMA_signal_4190, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4053, RoundOutput[30]}), .a ({new_AGEMA_signal_4929, new_AGEMA_signal_4925}), .c ({new_AGEMA_signal_4192, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4054, RoundOutput[31]}), .a ({new_AGEMA_signal_4937, new_AGEMA_signal_4933}), .c ({new_AGEMA_signal_4194, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_3313, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_4943, new_AGEMA_signal_4940}), .clk (clk), .r ({Fresh[129], Fresh[128]}), .c ({new_AGEMA_signal_3359, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_4949, new_AGEMA_signal_4946}), .clk (clk), .r ({Fresh[131], Fresh[130]}), .c ({new_AGEMA_signal_3314, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_4955, new_AGEMA_signal_4952}), .clk (clk), .r ({Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_3315, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_3312, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_4961, new_AGEMA_signal_4958}), .clk (clk), .r ({Fresh[135], Fresh[134]}), .c ({new_AGEMA_signal_3360, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_4967, new_AGEMA_signal_4964}), .clk (clk), .r ({Fresh[137], Fresh[136]}), .c ({new_AGEMA_signal_3316, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_4973, new_AGEMA_signal_4970}), .clk (clk), .r ({Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_3317, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_4979, new_AGEMA_signal_4976}), .clk (clk), .r ({Fresh[141], Fresh[140]}), .c ({new_AGEMA_signal_3361, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_3358, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_4985, new_AGEMA_signal_4982}), .clk (clk), .r ({Fresh[143], Fresh[142]}), .c ({new_AGEMA_signal_3406, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_4991, new_AGEMA_signal_4988}), .clk (clk), .r ({Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_3362, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_3313, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_4997, new_AGEMA_signal_4994}), .clk (clk), .r ({Fresh[147], Fresh[146]}), .c ({new_AGEMA_signal_3363, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_3297, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_5003, new_AGEMA_signal_5000}), .clk (clk), .r ({Fresh[149], Fresh[148]}), .c ({new_AGEMA_signal_3318, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_3296, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_5009, new_AGEMA_signal_5006}), .clk (clk), .r ({Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_3319, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_3312, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5015, new_AGEMA_signal_5012}), .clk (clk), .r ({Fresh[153], Fresh[152]}), .c ({new_AGEMA_signal_3364, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_3295, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_5021, new_AGEMA_signal_5018}), .clk (clk), .r ({Fresh[155], Fresh[154]}), .c ({new_AGEMA_signal_3320, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_3294, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_5027, new_AGEMA_signal_5024}), .clk (clk), .r ({Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_3321, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_3311, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5033, new_AGEMA_signal_5030}), .clk (clk), .r ({Fresh[159], Fresh[158]}), .c ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_3358, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5039, new_AGEMA_signal_5036}), .clk (clk), .r ({Fresh[161], Fresh[160]}), .c ({new_AGEMA_signal_3407, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_3310, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5045, new_AGEMA_signal_5042}), .clk (clk), .r ({Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_3366, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_3407, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_3316, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_3318, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_3359, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_3315, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_3408, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_3314, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_3363, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_3409, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_3362, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_3364, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_3410, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_3360, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_3411, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_3407, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_3411, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_3359, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_3409, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_3448, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_3317, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_3320, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_3368, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_3361, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_3406, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_3449, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_3406, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_3410, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_3450, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_3321, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_3408, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_3451, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_3315, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_3317, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_3369, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_3316, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_3482, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_3361, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_3365, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_3412, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_3363, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_3413, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_3318, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_3483, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_3319, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_3414, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_3364, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_3368, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_3415, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_3366, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_3410, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_3452, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_3446, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_3484, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_3367, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_3448, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_3485, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_3409, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_3369, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_3453, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_3415, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_3408, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_3454, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_3413, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_3449, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_3486, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3450, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_3487, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_3448, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_3449, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_3488, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_3368, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_3450, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_3489, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_3451, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_3412, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_3490, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_3451, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_3414, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_3491, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3486, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_3483, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_3488, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_3452, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_3490, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3485, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_3484, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_3453, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_3530, SubBytesOutput[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_3487, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_3491, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_3531, SubBytesOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_3482, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_3489, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_3447, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_3454, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_3492, SubBytesOutput[0]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_3325, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5051, new_AGEMA_signal_5048}), .clk (clk), .r ({Fresh[165], Fresh[164]}), .c ({new_AGEMA_signal_3371, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_5057, new_AGEMA_signal_5054}), .clk (clk), .r ({Fresh[167], Fresh[166]}), .c ({new_AGEMA_signal_3326, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5063, new_AGEMA_signal_5060}), .clk (clk), .r ({Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_3327, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_3324, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5069, new_AGEMA_signal_5066}), .clk (clk), .r ({Fresh[171], Fresh[170]}), .c ({new_AGEMA_signal_3372, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5075, new_AGEMA_signal_5072}), .clk (clk), .r ({Fresh[173], Fresh[172]}), .c ({new_AGEMA_signal_3328, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5081, new_AGEMA_signal_5078}), .clk (clk), .r ({Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_3329, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5087, new_AGEMA_signal_5084}), .clk (clk), .r ({Fresh[177], Fresh[176]}), .c ({new_AGEMA_signal_3373, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_3370, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5093, new_AGEMA_signal_5090}), .clk (clk), .r ({Fresh[179], Fresh[178]}), .c ({new_AGEMA_signal_3416, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5099, new_AGEMA_signal_5096}), .clk (clk), .r ({Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_3374, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_3325, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_5105, new_AGEMA_signal_5102}), .clk (clk), .r ({Fresh[183], Fresh[182]}), .c ({new_AGEMA_signal_3375, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_3301, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_5111, new_AGEMA_signal_5108}), .clk (clk), .r ({Fresh[185], Fresh[184]}), .c ({new_AGEMA_signal_3330, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_3300, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5117, new_AGEMA_signal_5114}), .clk (clk), .r ({Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_3331, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_3324, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5123, new_AGEMA_signal_5120}), .clk (clk), .r ({Fresh[189], Fresh[188]}), .c ({new_AGEMA_signal_3376, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_3299, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_5129, new_AGEMA_signal_5126}), .clk (clk), .r ({Fresh[191], Fresh[190]}), .c ({new_AGEMA_signal_3332, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_3298, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_5135, new_AGEMA_signal_5132}), .clk (clk), .r ({Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_3333, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_3323, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5141, new_AGEMA_signal_5138}), .clk (clk), .r ({Fresh[195], Fresh[194]}), .c ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_3370, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5147, new_AGEMA_signal_5144}), .clk (clk), .r ({Fresh[197], Fresh[196]}), .c ({new_AGEMA_signal_3417, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_3322, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5153, new_AGEMA_signal_5150}), .clk (clk), .r ({Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_3378, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_3417, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_3328, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_3330, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_3371, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_3327, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_3418, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_3326, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_3375, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_3419, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_3374, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_3376, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_3420, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_3372, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_3421, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_3417, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_3421, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_3371, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_3419, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_3457, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_3329, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_3332, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_3380, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_3373, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_3416, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_3458, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_3416, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_3420, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_3459, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_3333, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_3418, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_3460, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_3327, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_3329, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_3381, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_3328, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_3493, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_3373, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_3377, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_3422, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_3375, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_3423, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_3330, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_3494, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_3331, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_3424, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_3376, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_3380, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_3425, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_3378, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_3420, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_3461, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_3455, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_3495, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_3379, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_3457, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_3496, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_3419, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_3381, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_3462, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_3425, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_3418, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_3463, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_3423, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_3458, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_3497, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3459, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_3498, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_3457, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_3458, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_3499, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_3380, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_3459, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_3500, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_3460, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_3422, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_3501, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_3460, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_3424, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_3502, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3497, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_3494, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_3499, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_3461, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_3501, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3496, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_3495, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_3462, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_3498, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_3502, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_3493, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_3500, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_3456, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_3463, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_3337, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5159, new_AGEMA_signal_5156}), .clk (clk), .r ({Fresh[201], Fresh[200]}), .c ({new_AGEMA_signal_3383, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_5165, new_AGEMA_signal_5162}), .clk (clk), .r ({Fresh[203], Fresh[202]}), .c ({new_AGEMA_signal_3338, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5171, new_AGEMA_signal_5168}), .clk (clk), .r ({Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_3339, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_3336, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5177, new_AGEMA_signal_5174}), .clk (clk), .r ({Fresh[207], Fresh[206]}), .c ({new_AGEMA_signal_3384, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5183, new_AGEMA_signal_5180}), .clk (clk), .r ({Fresh[209], Fresh[208]}), .c ({new_AGEMA_signal_3340, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5189, new_AGEMA_signal_5186}), .clk (clk), .r ({Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_3341, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5195, new_AGEMA_signal_5192}), .clk (clk), .r ({Fresh[213], Fresh[212]}), .c ({new_AGEMA_signal_3385, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_3382, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5201, new_AGEMA_signal_5198}), .clk (clk), .r ({Fresh[215], Fresh[214]}), .c ({new_AGEMA_signal_3426, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5207, new_AGEMA_signal_5204}), .clk (clk), .r ({Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_3386, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_3337, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_5213, new_AGEMA_signal_5210}), .clk (clk), .r ({Fresh[219], Fresh[218]}), .c ({new_AGEMA_signal_3387, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_3305, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_5219, new_AGEMA_signal_5216}), .clk (clk), .r ({Fresh[221], Fresh[220]}), .c ({new_AGEMA_signal_3342, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_3304, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_5225, new_AGEMA_signal_5222}), .clk (clk), .r ({Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_3343, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_3336, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5231, new_AGEMA_signal_5228}), .clk (clk), .r ({Fresh[225], Fresh[224]}), .c ({new_AGEMA_signal_3388, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_3303, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_5237, new_AGEMA_signal_5234}), .clk (clk), .r ({Fresh[227], Fresh[226]}), .c ({new_AGEMA_signal_3344, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_3302, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_5243, new_AGEMA_signal_5240}), .clk (clk), .r ({Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_3345, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_3335, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5249, new_AGEMA_signal_5246}), .clk (clk), .r ({Fresh[231], Fresh[230]}), .c ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_3382, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5255, new_AGEMA_signal_5252}), .clk (clk), .r ({Fresh[233], Fresh[232]}), .c ({new_AGEMA_signal_3427, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_3334, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5261, new_AGEMA_signal_5258}), .clk (clk), .r ({Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_3390, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_3427, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_3340, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_3342, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_3383, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_3339, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_3428, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_3338, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_3387, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_3429, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_3386, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_3388, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_3430, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_3384, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_3431, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_3427, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_3431, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_3383, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_3429, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_3466, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_3341, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_3344, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_3392, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_3385, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_3426, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_3467, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_3426, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_3430, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_3468, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_3345, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_3428, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_3469, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_3339, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_3341, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_3393, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_3340, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_3504, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_3385, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_3389, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_3432, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_3387, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_3433, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_3342, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_3505, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_3343, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_3434, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_3388, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_3392, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_3435, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_3390, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_3430, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_3470, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_3464, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_3506, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_3391, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_3466, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_3507, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_3429, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_3393, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_3471, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_3435, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_3428, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_3472, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_3433, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_3467, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_3508, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3468, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_3509, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_3466, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_3467, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_3510, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_3392, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_3468, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_3511, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_3469, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_3432, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_3512, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_3469, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_3434, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_3513, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3508, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_3505, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_3510, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_3470, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_3512, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3507, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_3506, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_3471, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_3509, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_3513, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_3504, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_3511, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_3465, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_3472, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_3349, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5267, new_AGEMA_signal_5264}), .clk (clk), .r ({Fresh[237], Fresh[236]}), .c ({new_AGEMA_signal_3395, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_5273, new_AGEMA_signal_5270}), .clk (clk), .r ({Fresh[239], Fresh[238]}), .c ({new_AGEMA_signal_3350, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5279, new_AGEMA_signal_5276}), .clk (clk), .r ({Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_3351, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_3348, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5285, new_AGEMA_signal_5282}), .clk (clk), .r ({Fresh[243], Fresh[242]}), .c ({new_AGEMA_signal_3396, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5291, new_AGEMA_signal_5288}), .clk (clk), .r ({Fresh[245], Fresh[244]}), .c ({new_AGEMA_signal_3352, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5297, new_AGEMA_signal_5294}), .clk (clk), .r ({Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_3353, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5303, new_AGEMA_signal_5300}), .clk (clk), .r ({Fresh[249], Fresh[248]}), .c ({new_AGEMA_signal_3397, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_3394, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5309, new_AGEMA_signal_5306}), .clk (clk), .r ({Fresh[251], Fresh[250]}), .c ({new_AGEMA_signal_3436, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5315, new_AGEMA_signal_5312}), .clk (clk), .r ({Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_3398, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_3349, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_5321, new_AGEMA_signal_5318}), .clk (clk), .r ({Fresh[255], Fresh[254]}), .c ({new_AGEMA_signal_3399, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_3309, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_5327, new_AGEMA_signal_5324}), .clk (clk), .r ({Fresh[257], Fresh[256]}), .c ({new_AGEMA_signal_3354, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_3308, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_5333, new_AGEMA_signal_5330}), .clk (clk), .r ({Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_3355, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_3348, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5339, new_AGEMA_signal_5336}), .clk (clk), .r ({Fresh[261], Fresh[260]}), .c ({new_AGEMA_signal_3400, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_3307, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_5345, new_AGEMA_signal_5342}), .clk (clk), .r ({Fresh[263], Fresh[262]}), .c ({new_AGEMA_signal_3356, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_3306, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_5351, new_AGEMA_signal_5348}), .clk (clk), .r ({Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_3357, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_3347, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5357, new_AGEMA_signal_5354}), .clk (clk), .r ({Fresh[267], Fresh[266]}), .c ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_3394, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5363, new_AGEMA_signal_5360}), .clk (clk), .r ({Fresh[269], Fresh[268]}), .c ({new_AGEMA_signal_3437, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_3346, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5369, new_AGEMA_signal_5366}), .clk (clk), .r ({Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_3402, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_3437, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_3352, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_3354, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_3395, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_3351, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_3438, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_3350, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_3399, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_3439, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_3398, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_3400, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_3440, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_3396, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_3441, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_3437, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_3441, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_3395, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_3439, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_3475, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_3353, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_3356, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_3404, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_3397, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_3436, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_3476, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_3436, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_3440, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_3477, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_3357, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_3438, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_3478, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_3351, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_3353, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_3405, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_3352, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_3515, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_3397, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_3401, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_3442, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_3399, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_3443, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_3354, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_3516, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_3355, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_3444, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_3400, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_3404, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_3445, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_3402, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_3440, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_3479, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_3473, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_3517, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_3403, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_3475, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_3518, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_3439, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_3405, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_3480, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_3445, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_3438, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_3481, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_3443, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_3476, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_3519, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3477, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_3520, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_3475, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_3476, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_3521, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_3404, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_3477, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_3522, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_3478, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_3442, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_3523, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_3478, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_3444, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_3524, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3519, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_3516, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_3521, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_3479, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_3523, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3518, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_3517, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_3480, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_3520, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_3524, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_3515, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_3522, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_3474, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_3481, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U96 ( .a ({new_AGEMA_signal_3720, MixColumnsIns_n64}), .b ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_3866, MixColumnsOutput[9]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U95 ( .a ({new_AGEMA_signal_3646, MixColumnsIns_n63}), .b ({new_AGEMA_signal_3642, MixColumnsIns_n62}), .c ({new_AGEMA_signal_3720, MixColumnsIns_n64}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U94 ( .a ({new_AGEMA_signal_3625, MixColumnsIns_n61}), .b ({new_AGEMA_signal_3567, MixColumnsIns_n60}), .c ({new_AGEMA_signal_3721, MixColumnsOutput[8]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U93 ( .a ({new_AGEMA_signal_3577, MixColumnsIns_n59}), .b ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3625, MixColumnsIns_n61}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U92 ( .a ({new_AGEMA_signal_3626, MixColumnsIns_n58}), .b ({new_AGEMA_signal_3558, MixColumnsIns_n57}), .c ({new_AGEMA_signal_3722, MixColumnsOutput[7]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U91 ( .a ({new_AGEMA_signal_3569, MixColumnsIns_n56}), .b ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_3626, MixColumnsIns_n58}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U90 ( .a ({new_AGEMA_signal_3627, MixColumnsIns_n55}), .b ({new_AGEMA_signal_3559, MixColumnsIns_n54}), .c ({new_AGEMA_signal_3723, MixColumnsOutput[6]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U89 ( .a ({new_AGEMA_signal_3571, MixColumnsIns_n53}), .b ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3627, MixColumnsIns_n55}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U88 ( .a ({new_AGEMA_signal_3628, MixColumnsIns_n52}), .b ({new_AGEMA_signal_3560, MixColumnsIns_n51}), .c ({new_AGEMA_signal_3724, MixColumnsOutput[5]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U87 ( .a ({new_AGEMA_signal_3573, MixColumnsIns_n50}), .b ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3628, MixColumnsIns_n52}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U86 ( .a ({new_AGEMA_signal_3725, MixColumnsIns_n49}), .b ({new_AGEMA_signal_3633, MixColumnsIns_n48}), .c ({new_AGEMA_signal_3867, MixColumnsOutput[4]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U85 ( .a ({new_AGEMA_signal_3652, MixColumnsIns_n47}), .b ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_3725, MixColumnsIns_n49}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U84 ( .a ({new_AGEMA_signal_3726, MixColumnsIns_n46}), .b ({new_AGEMA_signal_3634, MixColumnsIns_n45}), .c ({new_AGEMA_signal_3868, MixColumnsOutput[3]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U83 ( .a ({new_AGEMA_signal_3654, MixColumnsIns_n44}), .b ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_3726, MixColumnsIns_n46}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U82 ( .a ({new_AGEMA_signal_3629, MixColumnsIns_n43}), .b ({new_AGEMA_signal_3558, MixColumnsIns_n57}), .c ({new_AGEMA_signal_3727, MixColumnsOutput[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U81 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3558, MixColumnsIns_n57}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U80 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3562, MixColumnsIns_n42}), .c ({new_AGEMA_signal_3629, MixColumnsIns_n43}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U79 ( .a ({new_AGEMA_signal_3630, MixColumnsIns_n41}), .b ({new_AGEMA_signal_3559, MixColumnsIns_n54}), .c ({new_AGEMA_signal_3728, MixColumnsOutput[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U78 ( .a ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .b ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3559, MixColumnsIns_n54}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U77 ( .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_3563, MixColumnsIns_n40}), .c ({new_AGEMA_signal_3630, MixColumnsIns_n41}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U76 ( .a ({new_AGEMA_signal_3631, MixColumnsIns_n39}), .b ({new_AGEMA_signal_3561, MixColumnsIns_n38}), .c ({new_AGEMA_signal_3729, MixColumnsOutput[2]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U75 ( .a ({new_AGEMA_signal_3575, MixColumnsIns_n37}), .b ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3631, MixColumnsIns_n39}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U74 ( .a ({new_AGEMA_signal_3632, MixColumnsIns_n36}), .b ({new_AGEMA_signal_3560, MixColumnsIns_n51}), .c ({new_AGEMA_signal_3730, MixColumnsOutput[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U73 ( .a ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .b ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_3560, MixColumnsIns_n51}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U72 ( .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_3564, MixColumnsIns_n35}), .c ({new_AGEMA_signal_3632, MixColumnsIns_n36}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U71 ( .a ({new_AGEMA_signal_3731, MixColumnsIns_n34}), .b ({new_AGEMA_signal_3633, MixColumnsIns_n48}), .c ({new_AGEMA_signal_3869, MixColumnsOutput[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U70 ( .a ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .b ({new_AGEMA_signal_3578, MixColumnsIns_DoubleBytes[28]}), .c ({new_AGEMA_signal_3633, MixColumnsIns_n48}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U69 ( .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_3640, MixColumnsIns_n33}), .c ({new_AGEMA_signal_3731, MixColumnsIns_n34}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U68 ( .a ({new_AGEMA_signal_3732, MixColumnsIns_n32}), .b ({new_AGEMA_signal_3634, MixColumnsIns_n45}), .c ({new_AGEMA_signal_3870, MixColumnsOutput[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U67 ( .a ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .b ({new_AGEMA_signal_3579, MixColumnsIns_DoubleBytes[27]}), .c ({new_AGEMA_signal_3634, MixColumnsIns_n45}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U66 ( .a ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .b ({new_AGEMA_signal_3643, MixColumnsIns_n31}), .c ({new_AGEMA_signal_3732, MixColumnsIns_n32}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U65 ( .a ({new_AGEMA_signal_3635, MixColumnsIns_n30}), .b ({new_AGEMA_signal_3561, MixColumnsIns_n38}), .c ({new_AGEMA_signal_3733, MixColumnsOutput[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U64 ( .a ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .b ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_3561, MixColumnsIns_n38}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U63 ( .a ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .b ({new_AGEMA_signal_3565, MixColumnsIns_n29}), .c ({new_AGEMA_signal_3635, MixColumnsIns_n30}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U62 ( .a ({new_AGEMA_signal_3734, MixColumnsIns_n28}), .b ({new_AGEMA_signal_3641, MixColumnsIns_n27}), .c ({new_AGEMA_signal_3871, MixColumnsOutput[25]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U61 ( .a ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_3645, MixColumnsIns_n26}), .c ({new_AGEMA_signal_3734, MixColumnsIns_n28}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U60 ( .a ({new_AGEMA_signal_3636, MixColumnsIns_n25}), .b ({new_AGEMA_signal_3566, MixColumnsIns_n24}), .c ({new_AGEMA_signal_3735, MixColumnsOutput[24]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U59 ( .a ({new_AGEMA_signal_3576, MixColumnsIns_n23}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3636, MixColumnsIns_n25}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U58 ( .a ({new_AGEMA_signal_3637, MixColumnsIns_n22}), .b ({new_AGEMA_signal_3562, MixColumnsIns_n42}), .c ({new_AGEMA_signal_3736, MixColumnsOutput[23]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U57 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3562, MixColumnsIns_n42}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U56 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3568, MixColumnsIns_n21}), .c ({new_AGEMA_signal_3637, MixColumnsIns_n22}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U55 ( .a ({new_AGEMA_signal_3638, MixColumnsIns_n20}), .b ({new_AGEMA_signal_3563, MixColumnsIns_n40}), .c ({new_AGEMA_signal_3737, MixColumnsOutput[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U54 ( .a ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .b ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3563, MixColumnsIns_n40}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U53 ( .a ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .b ({new_AGEMA_signal_3570, MixColumnsIns_n19}), .c ({new_AGEMA_signal_3638, MixColumnsIns_n20}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U52 ( .a ({new_AGEMA_signal_3639, MixColumnsIns_n18}), .b ({new_AGEMA_signal_3564, MixColumnsIns_n35}), .c ({new_AGEMA_signal_3738, MixColumnsOutput[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U51 ( .a ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .b ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_3564, MixColumnsIns_n35}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U50 ( .a ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .b ({new_AGEMA_signal_3572, MixColumnsIns_n17}), .c ({new_AGEMA_signal_3639, MixColumnsIns_n18}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U49 ( .a ({new_AGEMA_signal_3739, MixColumnsIns_n16}), .b ({new_AGEMA_signal_3640, MixColumnsIns_n33}), .c ({new_AGEMA_signal_3872, MixColumnsOutput[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U48 ( .a ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .b ({new_AGEMA_signal_3581, MixColumnsIns_DoubleBytes[20]}), .c ({new_AGEMA_signal_3640, MixColumnsIns_n33}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U47 ( .a ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .b ({new_AGEMA_signal_3651, MixColumnsIns_n15}), .c ({new_AGEMA_signal_3739, MixColumnsIns_n16}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U46 ( .a ({new_AGEMA_signal_3740, MixColumnsIns_n14}), .b ({new_AGEMA_signal_3641, MixColumnsIns_n27}), .c ({new_AGEMA_signal_3873, MixColumnsOutput[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U45 ( .a ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .b ({new_AGEMA_signal_3580, MixColumnsIns_DoubleBytes[25]}), .c ({new_AGEMA_signal_3641, MixColumnsIns_n27}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U44 ( .a ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .b ({new_AGEMA_signal_3642, MixColumnsIns_n62}), .c ({new_AGEMA_signal_3740, MixColumnsIns_n14}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U43 ( .a ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .b ({new_AGEMA_signal_3589, MixColumnsIns_DoubleBytes[1]}), .c ({new_AGEMA_signal_3642, MixColumnsIns_n62}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U42 ( .a ({new_AGEMA_signal_3741, MixColumnsIns_n13}), .b ({new_AGEMA_signal_3643, MixColumnsIns_n31}), .c ({new_AGEMA_signal_3874, MixColumnsOutput[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U41 ( .a ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .b ({new_AGEMA_signal_3582, MixColumnsIns_DoubleBytes[19]}), .c ({new_AGEMA_signal_3643, MixColumnsIns_n31}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U40 ( .a ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .b ({new_AGEMA_signal_3653, MixColumnsIns_n12}), .c ({new_AGEMA_signal_3741, MixColumnsIns_n13}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U39 ( .a ({new_AGEMA_signal_3644, MixColumnsIns_n11}), .b ({new_AGEMA_signal_3565, MixColumnsIns_n29}), .c ({new_AGEMA_signal_3742, MixColumnsOutput[18]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U38 ( .a ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .b ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_3565, MixColumnsIns_n29}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U37 ( .a ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .b ({new_AGEMA_signal_3574, MixColumnsIns_n10}), .c ({new_AGEMA_signal_3644, MixColumnsIns_n11}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U36 ( .a ({new_AGEMA_signal_3743, MixColumnsIns_n9}), .b ({new_AGEMA_signal_3645, MixColumnsIns_n26}), .c ({new_AGEMA_signal_3875, MixColumnsOutput[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U35 ( .a ({new_AGEMA_signal_3583, MixColumnsIns_DoubleBytes[17]}), .b ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_3645, MixColumnsIns_n26}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U34 ( .a ({new_AGEMA_signal_3646, MixColumnsIns_n63}), .b ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_3743, MixColumnsIns_n9}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U33 ( .a ({new_AGEMA_signal_3586, MixColumnsIns_DoubleBytes[9]}), .b ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_3646, MixColumnsIns_n63}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U32 ( .a ({new_AGEMA_signal_3647, MixColumnsIns_n8}), .b ({new_AGEMA_signal_3566, MixColumnsIns_n24}), .c ({new_AGEMA_signal_3744, MixColumnsOutput[16]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U31 ( .a ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .b ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3566, MixColumnsIns_n24}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U30 ( .a ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .b ({new_AGEMA_signal_3567, MixColumnsIns_n60}), .c ({new_AGEMA_signal_3647, MixColumnsIns_n8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U29 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3567, MixColumnsIns_n60}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U28 ( .a ({new_AGEMA_signal_3648, MixColumnsIns_n7}), .b ({new_AGEMA_signal_3568, MixColumnsIns_n21}), .c ({new_AGEMA_signal_3745, MixColumnsOutput[15]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U27 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3568, MixColumnsIns_n21}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U26 ( .a ({new_AGEMA_signal_3569, MixColumnsIns_n56}), .b ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3648, MixColumnsIns_n7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U25 ( .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3569, MixColumnsIns_n56}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U24 ( .a ({new_AGEMA_signal_3649, MixColumnsIns_n6}), .b ({new_AGEMA_signal_3570, MixColumnsIns_n19}), .c ({new_AGEMA_signal_3746, MixColumnsOutput[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U23 ( .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .b ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3570, MixColumnsIns_n19}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U22 ( .a ({new_AGEMA_signal_3571, MixColumnsIns_n53}), .b ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3649, MixColumnsIns_n6}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U21 ( .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3571, MixColumnsIns_n53}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U20 ( .a ({new_AGEMA_signal_3650, MixColumnsIns_n5}), .b ({new_AGEMA_signal_3572, MixColumnsIns_n17}), .c ({new_AGEMA_signal_3747, MixColumnsOutput[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U19 ( .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .b ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_3572, MixColumnsIns_n17}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U18 ( .a ({new_AGEMA_signal_3573, MixColumnsIns_n50}), .b ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3650, MixColumnsIns_n5}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U17 ( .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3573, MixColumnsIns_n50}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U16 ( .a ({new_AGEMA_signal_3748, MixColumnsIns_n4}), .b ({new_AGEMA_signal_3651, MixColumnsIns_n15}), .c ({new_AGEMA_signal_3876, MixColumnsOutput[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U15 ( .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .b ({new_AGEMA_signal_3584, MixColumnsIns_DoubleBytes[12]}), .c ({new_AGEMA_signal_3651, MixColumnsIns_n15}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U14 ( .a ({new_AGEMA_signal_3652, MixColumnsIns_n47}), .b ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_3748, MixColumnsIns_n4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U13 ( .a ({new_AGEMA_signal_3587, MixColumnsIns_DoubleBytes[4]}), .b ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_3652, MixColumnsIns_n47}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U12 ( .a ({new_AGEMA_signal_3749, MixColumnsIns_n3}), .b ({new_AGEMA_signal_3653, MixColumnsIns_n12}), .c ({new_AGEMA_signal_3877, MixColumnsOutput[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U11 ( .a ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .b ({new_AGEMA_signal_3585, MixColumnsIns_DoubleBytes[11]}), .c ({new_AGEMA_signal_3653, MixColumnsIns_n12}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U10 ( .a ({new_AGEMA_signal_3654, MixColumnsIns_n44}), .b ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_3749, MixColumnsIns_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U9 ( .a ({new_AGEMA_signal_3588, MixColumnsIns_DoubleBytes[3]}), .b ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_3654, MixColumnsIns_n44}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U8 ( .a ({new_AGEMA_signal_3655, MixColumnsIns_n2}), .b ({new_AGEMA_signal_3574, MixColumnsIns_n10}), .c ({new_AGEMA_signal_3750, MixColumnsOutput[10]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U7 ( .a ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .b ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_3574, MixColumnsIns_n10}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U6 ( .a ({new_AGEMA_signal_3575, MixColumnsIns_n37}), .b ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3655, MixColumnsIns_n2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U5 ( .a ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .b ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3575, MixColumnsIns_n37}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U4 ( .a ({new_AGEMA_signal_3656, MixColumnsIns_n1}), .b ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3751, MixColumnsOutput[0]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U3 ( .a ({new_AGEMA_signal_3577, MixColumnsIns_n59}), .b ({new_AGEMA_signal_3576, MixColumnsIns_n23}), .c ({new_AGEMA_signal_3656, MixColumnsIns_n1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U2 ( .a ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .b ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3576, MixColumnsIns_n23}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_U1 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3577, MixColumnsIns_n59}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_3578, MixColumnsIns_DoubleBytes[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3579, MixColumnsIns_DoubleBytes[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .b ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3580, MixColumnsIns_DoubleBytes[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_3581, MixColumnsIns_DoubleBytes[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3582, MixColumnsIns_DoubleBytes[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .b ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3583, MixColumnsIns_DoubleBytes[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_3584, MixColumnsIns_DoubleBytes[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3585, MixColumnsIns_DoubleBytes[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .b ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3586, MixColumnsIns_DoubleBytes[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .c ({new_AGEMA_signal_3587, MixColumnsIns_DoubleBytes[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .c ({new_AGEMA_signal_3588, MixColumnsIns_DoubleBytes[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) MixColumnsIns_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3589, MixColumnsIns_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_0_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3751, MixColumnsOutput[0]}), .a ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3878, ColumnOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_1_U1 ( .s (new_AGEMA_signal_5377), .b ({new_AGEMA_signal_3873, MixColumnsOutput[1]}), .a ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_4023, ColumnOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_2_U1 ( .s (new_AGEMA_signal_5377), .b ({new_AGEMA_signal_3729, MixColumnsOutput[2]}), .a ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .c ({new_AGEMA_signal_3879, ColumnOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_3_U1 ( .s (new_AGEMA_signal_5377), .b ({new_AGEMA_signal_3868, MixColumnsOutput[3]}), .a ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .c ({new_AGEMA_signal_4024, ColumnOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_4_U1 ( .s (new_AGEMA_signal_5377), .b ({new_AGEMA_signal_3867, MixColumnsOutput[4]}), .a ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_4025, ColumnOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_5_U1 ( .s (new_AGEMA_signal_5377), .b ({new_AGEMA_signal_3724, MixColumnsOutput[5]}), .a ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_3880, ColumnOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_6_U1 ( .s (new_AGEMA_signal_5377), .b ({new_AGEMA_signal_3723, MixColumnsOutput[6]}), .a ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_3881, ColumnOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_7_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3722, MixColumnsOutput[7]}), .a ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_3882, ColumnOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_8_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3721, MixColumnsOutput[8]}), .a ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3883, ColumnOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_9_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3866, MixColumnsOutput[9]}), .a ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_4026, ColumnOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_10_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3750, MixColumnsOutput[10]}), .a ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3884, ColumnOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_11_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3877, MixColumnsOutput[11]}), .a ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_4027, ColumnOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_12_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3876, MixColumnsOutput[12]}), .a ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_4028, ColumnOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_13_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3747, MixColumnsOutput[13]}), .a ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3885, ColumnOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_14_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3746, MixColumnsOutput[14]}), .a ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3886, ColumnOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_15_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3745, MixColumnsOutput[15]}), .a ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_3887, ColumnOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_16_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3744, MixColumnsOutput[16]}), .a ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3888, ColumnOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_17_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3875, MixColumnsOutput[17]}), .a ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_4029, ColumnOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_18_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3742, MixColumnsOutput[18]}), .a ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3889, ColumnOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_19_U1 ( .s (new_AGEMA_signal_5373), .b ({new_AGEMA_signal_3874, MixColumnsOutput[19]}), .a ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_4030, ColumnOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_20_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3872, MixColumnsOutput[20]}), .a ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_4031, ColumnOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_21_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3738, MixColumnsOutput[21]}), .a ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3890, ColumnOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_22_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3737, MixColumnsOutput[22]}), .a ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3891, ColumnOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_23_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3736, MixColumnsOutput[23]}), .a ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3892, ColumnOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_24_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3735, MixColumnsOutput[24]}), .a ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3893, ColumnOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_25_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3871, MixColumnsOutput[25]}), .a ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_4032, ColumnOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_26_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3733, MixColumnsOutput[26]}), .a ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3894, ColumnOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_27_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3870, MixColumnsOutput[27]}), .a ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_4033, ColumnOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_28_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3869, MixColumnsOutput[28]}), .a ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_4034, ColumnOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_29_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3730, MixColumnsOutput[29]}), .a ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3895, ColumnOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_30_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3728, MixColumnsOutput[30]}), .a ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3896, ColumnOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxMCOut_mux_inst_31_U1 ( .s (new_AGEMA_signal_5381), .b ({new_AGEMA_signal_3727, MixColumnsOutput[31]}), .a ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3897, ColumnOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_0_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3878, ColumnOutput[0]}), .a ({new_AGEMA_signal_5393, new_AGEMA_signal_5389}), .c ({new_AGEMA_signal_4035, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_1_U1 ( .s (new_AGEMA_signal_5397), .b ({new_AGEMA_signal_4023, ColumnOutput[1]}), .a ({new_AGEMA_signal_5405, new_AGEMA_signal_5401}), .c ({new_AGEMA_signal_4195, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_2_U1 ( .s (new_AGEMA_signal_5409), .b ({new_AGEMA_signal_3879, ColumnOutput[2]}), .a ({new_AGEMA_signal_5417, new_AGEMA_signal_5413}), .c ({new_AGEMA_signal_4036, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_3_U1 ( .s (new_AGEMA_signal_5421), .b ({new_AGEMA_signal_4024, ColumnOutput[3]}), .a ({new_AGEMA_signal_5429, new_AGEMA_signal_5425}), .c ({new_AGEMA_signal_4196, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_4_U1 ( .s (new_AGEMA_signal_5433), .b ({new_AGEMA_signal_4025, ColumnOutput[4]}), .a ({new_AGEMA_signal_5441, new_AGEMA_signal_5437}), .c ({new_AGEMA_signal_4197, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_5_U1 ( .s (new_AGEMA_signal_5445), .b ({new_AGEMA_signal_3880, ColumnOutput[5]}), .a ({new_AGEMA_signal_5453, new_AGEMA_signal_5449}), .c ({new_AGEMA_signal_4037, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_6_U1 ( .s (new_AGEMA_signal_5457), .b ({new_AGEMA_signal_3881, ColumnOutput[6]}), .a ({new_AGEMA_signal_5465, new_AGEMA_signal_5461}), .c ({new_AGEMA_signal_4038, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_7_U1 ( .s (new_AGEMA_signal_5397), .b ({new_AGEMA_signal_3882, ColumnOutput[7]}), .a ({new_AGEMA_signal_5473, new_AGEMA_signal_5469}), .c ({new_AGEMA_signal_4039, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_8_U1 ( .s (new_AGEMA_signal_5433), .b ({new_AGEMA_signal_3883, ColumnOutput[8]}), .a ({new_AGEMA_signal_5481, new_AGEMA_signal_5477}), .c ({new_AGEMA_signal_4040, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_9_U1 ( .s (new_AGEMA_signal_5397), .b ({new_AGEMA_signal_4026, ColumnOutput[9]}), .a ({new_AGEMA_signal_5489, new_AGEMA_signal_5485}), .c ({new_AGEMA_signal_4198, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_10_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3884, ColumnOutput[10]}), .a ({new_AGEMA_signal_5497, new_AGEMA_signal_5493}), .c ({new_AGEMA_signal_4041, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_11_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_4027, ColumnOutput[11]}), .a ({new_AGEMA_signal_5505, new_AGEMA_signal_5501}), .c ({new_AGEMA_signal_4199, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_12_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_4028, ColumnOutput[12]}), .a ({new_AGEMA_signal_5513, new_AGEMA_signal_5509}), .c ({new_AGEMA_signal_4200, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_13_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3885, ColumnOutput[13]}), .a ({new_AGEMA_signal_5521, new_AGEMA_signal_5517}), .c ({new_AGEMA_signal_4042, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_14_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3886, ColumnOutput[14]}), .a ({new_AGEMA_signal_5529, new_AGEMA_signal_5525}), .c ({new_AGEMA_signal_4043, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_15_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3887, ColumnOutput[15]}), .a ({new_AGEMA_signal_5537, new_AGEMA_signal_5533}), .c ({new_AGEMA_signal_4044, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_16_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3888, ColumnOutput[16]}), .a ({new_AGEMA_signal_5545, new_AGEMA_signal_5541}), .c ({new_AGEMA_signal_4045, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_17_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_4029, ColumnOutput[17]}), .a ({new_AGEMA_signal_5553, new_AGEMA_signal_5549}), .c ({new_AGEMA_signal_4201, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_18_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_3889, ColumnOutput[18]}), .a ({new_AGEMA_signal_5561, new_AGEMA_signal_5557}), .c ({new_AGEMA_signal_4046, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_19_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_4030, ColumnOutput[19]}), .a ({new_AGEMA_signal_5569, new_AGEMA_signal_5565}), .c ({new_AGEMA_signal_4202, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_20_U1 ( .s (new_AGEMA_signal_5409), .b ({new_AGEMA_signal_4031, ColumnOutput[20]}), .a ({new_AGEMA_signal_5577, new_AGEMA_signal_5573}), .c ({new_AGEMA_signal_4203, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_21_U1 ( .s (new_AGEMA_signal_5421), .b ({new_AGEMA_signal_3890, ColumnOutput[21]}), .a ({new_AGEMA_signal_5585, new_AGEMA_signal_5581}), .c ({new_AGEMA_signal_4047, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_22_U1 ( .s (new_AGEMA_signal_5433), .b ({new_AGEMA_signal_3891, ColumnOutput[22]}), .a ({new_AGEMA_signal_5593, new_AGEMA_signal_5589}), .c ({new_AGEMA_signal_4048, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_23_U1 ( .s (new_AGEMA_signal_5445), .b ({new_AGEMA_signal_3892, ColumnOutput[23]}), .a ({new_AGEMA_signal_5601, new_AGEMA_signal_5597}), .c ({new_AGEMA_signal_4049, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_24_U1 ( .s (new_AGEMA_signal_5457), .b ({new_AGEMA_signal_3893, ColumnOutput[24]}), .a ({new_AGEMA_signal_5609, new_AGEMA_signal_5605}), .c ({new_AGEMA_signal_4050, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_25_U1 ( .s (new_AGEMA_signal_5433), .b ({new_AGEMA_signal_4032, ColumnOutput[25]}), .a ({new_AGEMA_signal_5617, new_AGEMA_signal_5613}), .c ({new_AGEMA_signal_4204, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_26_U1 ( .s (new_AGEMA_signal_5445), .b ({new_AGEMA_signal_3894, ColumnOutput[26]}), .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5621}), .c ({new_AGEMA_signal_4051, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_27_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_4033, ColumnOutput[27]}), .a ({new_AGEMA_signal_5633, new_AGEMA_signal_5629}), .c ({new_AGEMA_signal_4205, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_28_U1 ( .s (new_AGEMA_signal_5385), .b ({new_AGEMA_signal_4034, ColumnOutput[28]}), .a ({new_AGEMA_signal_5641, new_AGEMA_signal_5637}), .c ({new_AGEMA_signal_4206, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_29_U1 ( .s (new_AGEMA_signal_5397), .b ({new_AGEMA_signal_3895, ColumnOutput[29]}), .a ({new_AGEMA_signal_5649, new_AGEMA_signal_5645}), .c ({new_AGEMA_signal_4052, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_30_U1 ( .s (new_AGEMA_signal_5409), .b ({new_AGEMA_signal_3896, ColumnOutput[30]}), .a ({new_AGEMA_signal_5657, new_AGEMA_signal_5653}), .c ({new_AGEMA_signal_4053, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxRound_mux_inst_31_U1 ( .s (new_AGEMA_signal_5421), .b ({new_AGEMA_signal_3897, ColumnOutput[31]}), .a ({new_AGEMA_signal_5665, new_AGEMA_signal_5661}), .c ({new_AGEMA_signal_4054, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3991, RoundKeyOutput[0]}), .a ({new_AGEMA_signal_5673, new_AGEMA_signal_5669}), .c ({new_AGEMA_signal_4056, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4126, RoundKeyOutput[1]}), .a ({new_AGEMA_signal_5681, new_AGEMA_signal_5677}), .c ({new_AGEMA_signal_4208, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4127, RoundKeyOutput[2]}), .a ({new_AGEMA_signal_5689, new_AGEMA_signal_5685}), .c ({new_AGEMA_signal_4210, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4128, RoundKeyOutput[3]}), .a ({new_AGEMA_signal_5697, new_AGEMA_signal_5693}), .c ({new_AGEMA_signal_4212, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4129, RoundKeyOutput[4]}), .a ({new_AGEMA_signal_5705, new_AGEMA_signal_5701}), .c ({new_AGEMA_signal_4214, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4130, RoundKeyOutput[5]}), .a ({new_AGEMA_signal_5713, new_AGEMA_signal_5709}), .c ({new_AGEMA_signal_4216, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4131, RoundKeyOutput[6]}), .a ({new_AGEMA_signal_5721, new_AGEMA_signal_5717}), .c ({new_AGEMA_signal_4218, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4132, RoundKeyOutput[7]}), .a ({new_AGEMA_signal_5729, new_AGEMA_signal_5725}), .c ({new_AGEMA_signal_4220, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3992, RoundKeyOutput[8]}), .a ({new_AGEMA_signal_5737, new_AGEMA_signal_5733}), .c ({new_AGEMA_signal_4058, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4133, RoundKeyOutput[9]}), .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5741}), .c ({new_AGEMA_signal_4222, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4134, RoundKeyOutput[10]}), .a ({new_AGEMA_signal_5753, new_AGEMA_signal_5749}), .c ({new_AGEMA_signal_4224, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4135, RoundKeyOutput[11]}), .a ({new_AGEMA_signal_5761, new_AGEMA_signal_5757}), .c ({new_AGEMA_signal_4226, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4136, RoundKeyOutput[12]}), .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5765}), .c ({new_AGEMA_signal_4228, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4137, RoundKeyOutput[13]}), .a ({new_AGEMA_signal_5777, new_AGEMA_signal_5773}), .c ({new_AGEMA_signal_4230, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4138, RoundKeyOutput[14]}), .a ({new_AGEMA_signal_5785, new_AGEMA_signal_5781}), .c ({new_AGEMA_signal_4232, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4139, RoundKeyOutput[15]}), .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5789}), .c ({new_AGEMA_signal_4234, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3993, RoundKeyOutput[16]}), .a ({new_AGEMA_signal_5801, new_AGEMA_signal_5797}), .c ({new_AGEMA_signal_4060, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4140, RoundKeyOutput[17]}), .a ({new_AGEMA_signal_5809, new_AGEMA_signal_5805}), .c ({new_AGEMA_signal_4236, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4141, RoundKeyOutput[18]}), .a ({new_AGEMA_signal_5817, new_AGEMA_signal_5813}), .c ({new_AGEMA_signal_4238, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4142, RoundKeyOutput[19]}), .a ({new_AGEMA_signal_5825, new_AGEMA_signal_5821}), .c ({new_AGEMA_signal_4240, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4143, RoundKeyOutput[20]}), .a ({new_AGEMA_signal_5833, new_AGEMA_signal_5829}), .c ({new_AGEMA_signal_4242, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4144, RoundKeyOutput[21]}), .a ({new_AGEMA_signal_5841, new_AGEMA_signal_5837}), .c ({new_AGEMA_signal_4244, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4145, RoundKeyOutput[22]}), .a ({new_AGEMA_signal_5849, new_AGEMA_signal_5845}), .c ({new_AGEMA_signal_4246, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4146, RoundKeyOutput[23]}), .a ({new_AGEMA_signal_5857, new_AGEMA_signal_5853}), .c ({new_AGEMA_signal_4248, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4147, RoundKeyOutput[24]}), .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5861}), .c ({new_AGEMA_signal_4250, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4265, RoundKeyOutput[25]}), .a ({new_AGEMA_signal_5873, new_AGEMA_signal_5869}), .c ({new_AGEMA_signal_4297, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4266, RoundKeyOutput[26]}), .a ({new_AGEMA_signal_5881, new_AGEMA_signal_5877}), .c ({new_AGEMA_signal_4299, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4267, RoundKeyOutput[27]}), .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5885}), .c ({new_AGEMA_signal_4301, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4268, RoundKeyOutput[28]}), .a ({new_AGEMA_signal_5897, new_AGEMA_signal_5893}), .c ({new_AGEMA_signal_4303, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4269, RoundKeyOutput[29]}), .a ({new_AGEMA_signal_5905, new_AGEMA_signal_5901}), .c ({new_AGEMA_signal_4305, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4270, RoundKeyOutput[30]}), .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5909}), .c ({new_AGEMA_signal_4307, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4271, RoundKeyOutput[31]}), .a ({new_AGEMA_signal_5921, new_AGEMA_signal_5917}), .c ({new_AGEMA_signal_4309, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3834, RoundKeyOutput[32]}), .a ({new_AGEMA_signal_5929, new_AGEMA_signal_5925}), .c ({new_AGEMA_signal_3899, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3994, RoundKeyOutput[33]}), .a ({new_AGEMA_signal_5937, new_AGEMA_signal_5933}), .c ({new_AGEMA_signal_4062, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3995, RoundKeyOutput[34]}), .a ({new_AGEMA_signal_5945, new_AGEMA_signal_5941}), .c ({new_AGEMA_signal_4064, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3996, RoundKeyOutput[35]}), .a ({new_AGEMA_signal_5953, new_AGEMA_signal_5949}), .c ({new_AGEMA_signal_4066, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3997, RoundKeyOutput[36]}), .a ({new_AGEMA_signal_5961, new_AGEMA_signal_5957}), .c ({new_AGEMA_signal_4068, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3998, RoundKeyOutput[37]}), .a ({new_AGEMA_signal_5969, new_AGEMA_signal_5965}), .c ({new_AGEMA_signal_4070, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3999, RoundKeyOutput[38]}), .a ({new_AGEMA_signal_5977, new_AGEMA_signal_5973}), .c ({new_AGEMA_signal_4072, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4000, RoundKeyOutput[39]}), .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5981}), .c ({new_AGEMA_signal_4074, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3835, RoundKeyOutput[40]}), .a ({new_AGEMA_signal_5993, new_AGEMA_signal_5989}), .c ({new_AGEMA_signal_3901, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4001, RoundKeyOutput[41]}), .a ({new_AGEMA_signal_6001, new_AGEMA_signal_5997}), .c ({new_AGEMA_signal_4076, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4002, RoundKeyOutput[42]}), .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6005}), .c ({new_AGEMA_signal_4078, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4003, RoundKeyOutput[43]}), .a ({new_AGEMA_signal_6017, new_AGEMA_signal_6013}), .c ({new_AGEMA_signal_4080, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4004, RoundKeyOutput[44]}), .a ({new_AGEMA_signal_6025, new_AGEMA_signal_6021}), .c ({new_AGEMA_signal_4082, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4005, RoundKeyOutput[45]}), .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6029}), .c ({new_AGEMA_signal_4084, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4006, RoundKeyOutput[46]}), .a ({new_AGEMA_signal_6041, new_AGEMA_signal_6037}), .c ({new_AGEMA_signal_4086, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4007, RoundKeyOutput[47]}), .a ({new_AGEMA_signal_6049, new_AGEMA_signal_6045}), .c ({new_AGEMA_signal_4088, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3836, RoundKeyOutput[48]}), .a ({new_AGEMA_signal_6057, new_AGEMA_signal_6053}), .c ({new_AGEMA_signal_3903, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4008, RoundKeyOutput[49]}), .a ({new_AGEMA_signal_6065, new_AGEMA_signal_6061}), .c ({new_AGEMA_signal_4090, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4009, RoundKeyOutput[50]}), .a ({new_AGEMA_signal_6073, new_AGEMA_signal_6069}), .c ({new_AGEMA_signal_4092, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4010, RoundKeyOutput[51]}), .a ({new_AGEMA_signal_6081, new_AGEMA_signal_6077}), .c ({new_AGEMA_signal_4094, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4011, RoundKeyOutput[52]}), .a ({new_AGEMA_signal_6089, new_AGEMA_signal_6085}), .c ({new_AGEMA_signal_4096, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4012, RoundKeyOutput[53]}), .a ({new_AGEMA_signal_6097, new_AGEMA_signal_6093}), .c ({new_AGEMA_signal_4098, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4013, RoundKeyOutput[54]}), .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6101}), .c ({new_AGEMA_signal_4100, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4014, RoundKeyOutput[55]}), .a ({new_AGEMA_signal_6113, new_AGEMA_signal_6109}), .c ({new_AGEMA_signal_4102, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4015, RoundKeyOutput[56]}), .a ({new_AGEMA_signal_6121, new_AGEMA_signal_6117}), .c ({new_AGEMA_signal_4104, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4148, RoundKeyOutput[57]}), .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6125}), .c ({new_AGEMA_signal_4252, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4149, RoundKeyOutput[58]}), .a ({new_AGEMA_signal_6137, new_AGEMA_signal_6133}), .c ({new_AGEMA_signal_4254, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4150, RoundKeyOutput[59]}), .a ({new_AGEMA_signal_6145, new_AGEMA_signal_6141}), .c ({new_AGEMA_signal_4256, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4151, RoundKeyOutput[60]}), .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6149}), .c ({new_AGEMA_signal_4258, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4152, RoundKeyOutput[61]}), .a ({new_AGEMA_signal_6161, new_AGEMA_signal_6157}), .c ({new_AGEMA_signal_4260, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4153, RoundKeyOutput[62]}), .a ({new_AGEMA_signal_6169, new_AGEMA_signal_6165}), .c ({new_AGEMA_signal_4262, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4154, RoundKeyOutput[63]}), .a ({new_AGEMA_signal_6177, new_AGEMA_signal_6173}), .c ({new_AGEMA_signal_4264, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3695, RoundKeyOutput[64]}), .a ({new_AGEMA_signal_6185, new_AGEMA_signal_6181}), .c ({new_AGEMA_signal_3753, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3837, RoundKeyOutput[65]}), .a ({new_AGEMA_signal_6193, new_AGEMA_signal_6189}), .c ({new_AGEMA_signal_3905, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3838, RoundKeyOutput[66]}), .a ({new_AGEMA_signal_6201, new_AGEMA_signal_6197}), .c ({new_AGEMA_signal_3907, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3839, RoundKeyOutput[67]}), .a ({new_AGEMA_signal_6209, new_AGEMA_signal_6205}), .c ({new_AGEMA_signal_3909, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3840, RoundKeyOutput[68]}), .a ({new_AGEMA_signal_6217, new_AGEMA_signal_6213}), .c ({new_AGEMA_signal_3911, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3841, RoundKeyOutput[69]}), .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6221}), .c ({new_AGEMA_signal_3913, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3842, RoundKeyOutput[70]}), .a ({new_AGEMA_signal_6233, new_AGEMA_signal_6229}), .c ({new_AGEMA_signal_3915, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3843, RoundKeyOutput[71]}), .a ({new_AGEMA_signal_6241, new_AGEMA_signal_6237}), .c ({new_AGEMA_signal_3917, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3696, RoundKeyOutput[72]}), .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6245}), .c ({new_AGEMA_signal_3755, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3844, RoundKeyOutput[73]}), .a ({new_AGEMA_signal_6257, new_AGEMA_signal_6253}), .c ({new_AGEMA_signal_3919, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3845, RoundKeyOutput[74]}), .a ({new_AGEMA_signal_6265, new_AGEMA_signal_6261}), .c ({new_AGEMA_signal_3921, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3846, RoundKeyOutput[75]}), .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6269}), .c ({new_AGEMA_signal_3923, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3847, RoundKeyOutput[76]}), .a ({new_AGEMA_signal_6281, new_AGEMA_signal_6277}), .c ({new_AGEMA_signal_3925, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3848, RoundKeyOutput[77]}), .a ({new_AGEMA_signal_6289, new_AGEMA_signal_6285}), .c ({new_AGEMA_signal_3927, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3849, RoundKeyOutput[78]}), .a ({new_AGEMA_signal_6297, new_AGEMA_signal_6293}), .c ({new_AGEMA_signal_3929, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3850, RoundKeyOutput[79]}), .a ({new_AGEMA_signal_6305, new_AGEMA_signal_6301}), .c ({new_AGEMA_signal_3931, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3697, RoundKeyOutput[80]}), .a ({new_AGEMA_signal_6313, new_AGEMA_signal_6309}), .c ({new_AGEMA_signal_3757, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3851, RoundKeyOutput[81]}), .a ({new_AGEMA_signal_6321, new_AGEMA_signal_6317}), .c ({new_AGEMA_signal_3933, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3852, RoundKeyOutput[82]}), .a ({new_AGEMA_signal_6329, new_AGEMA_signal_6325}), .c ({new_AGEMA_signal_3935, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3853, RoundKeyOutput[83]}), .a ({new_AGEMA_signal_6337, new_AGEMA_signal_6333}), .c ({new_AGEMA_signal_3937, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3854, RoundKeyOutput[84]}), .a ({new_AGEMA_signal_6345, new_AGEMA_signal_6341}), .c ({new_AGEMA_signal_3939, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3855, RoundKeyOutput[85]}), .a ({new_AGEMA_signal_6353, new_AGEMA_signal_6349}), .c ({new_AGEMA_signal_3941, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3856, RoundKeyOutput[86]}), .a ({new_AGEMA_signal_6361, new_AGEMA_signal_6357}), .c ({new_AGEMA_signal_3943, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3857, RoundKeyOutput[87]}), .a ({new_AGEMA_signal_6369, new_AGEMA_signal_6365}), .c ({new_AGEMA_signal_3945, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3858, RoundKeyOutput[88]}), .a ({new_AGEMA_signal_6377, new_AGEMA_signal_6373}), .c ({new_AGEMA_signal_3947, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4016, RoundKeyOutput[89]}), .a ({new_AGEMA_signal_6385, new_AGEMA_signal_6381}), .c ({new_AGEMA_signal_4106, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4017, RoundKeyOutput[90]}), .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6389}), .c ({new_AGEMA_signal_4108, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4018, RoundKeyOutput[91]}), .a ({new_AGEMA_signal_6401, new_AGEMA_signal_6397}), .c ({new_AGEMA_signal_4110, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4019, RoundKeyOutput[92]}), .a ({new_AGEMA_signal_6409, new_AGEMA_signal_6405}), .c ({new_AGEMA_signal_4112, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4020, RoundKeyOutput[93]}), .a ({new_AGEMA_signal_6417, new_AGEMA_signal_6413}), .c ({new_AGEMA_signal_4114, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4021, RoundKeyOutput[94]}), .a ({new_AGEMA_signal_6425, new_AGEMA_signal_6421}), .c ({new_AGEMA_signal_4116, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_4022, RoundKeyOutput[95]}), .a ({new_AGEMA_signal_6433, new_AGEMA_signal_6429}), .c ({new_AGEMA_signal_4118, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3622, RoundKeyOutput[96]}), .a ({new_AGEMA_signal_6441, new_AGEMA_signal_6437}), .c ({new_AGEMA_signal_3658, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3698, RoundKeyOutput[97]}), .a ({new_AGEMA_signal_6449, new_AGEMA_signal_6445}), .c ({new_AGEMA_signal_3759, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3699, RoundKeyOutput[98]}), .a ({new_AGEMA_signal_6457, new_AGEMA_signal_6453}), .c ({new_AGEMA_signal_3761, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3700, RoundKeyOutput[99]}), .a ({new_AGEMA_signal_6465, new_AGEMA_signal_6461}), .c ({new_AGEMA_signal_3763, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3701, RoundKeyOutput[100]}), .a ({new_AGEMA_signal_6473, new_AGEMA_signal_6469}), .c ({new_AGEMA_signal_3765, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3702, RoundKeyOutput[101]}), .a ({new_AGEMA_signal_6481, new_AGEMA_signal_6477}), .c ({new_AGEMA_signal_3767, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3703, RoundKeyOutput[102]}), .a ({new_AGEMA_signal_6489, new_AGEMA_signal_6485}), .c ({new_AGEMA_signal_3769, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3704, RoundKeyOutput[103]}), .a ({new_AGEMA_signal_6497, new_AGEMA_signal_6493}), .c ({new_AGEMA_signal_3771, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3623, RoundKeyOutput[104]}), .a ({new_AGEMA_signal_6505, new_AGEMA_signal_6501}), .c ({new_AGEMA_signal_3660, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3705, RoundKeyOutput[105]}), .a ({new_AGEMA_signal_6513, new_AGEMA_signal_6509}), .c ({new_AGEMA_signal_3773, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3706, RoundKeyOutput[106]}), .a ({new_AGEMA_signal_6521, new_AGEMA_signal_6517}), .c ({new_AGEMA_signal_3775, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3707, RoundKeyOutput[107]}), .a ({new_AGEMA_signal_6529, new_AGEMA_signal_6525}), .c ({new_AGEMA_signal_3777, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3708, RoundKeyOutput[108]}), .a ({new_AGEMA_signal_6537, new_AGEMA_signal_6533}), .c ({new_AGEMA_signal_3779, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3709, RoundKeyOutput[109]}), .a ({new_AGEMA_signal_6545, new_AGEMA_signal_6541}), .c ({new_AGEMA_signal_3781, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3710, RoundKeyOutput[110]}), .a ({new_AGEMA_signal_6553, new_AGEMA_signal_6549}), .c ({new_AGEMA_signal_3783, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3711, RoundKeyOutput[111]}), .a ({new_AGEMA_signal_6561, new_AGEMA_signal_6557}), .c ({new_AGEMA_signal_3785, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3624, RoundKeyOutput[112]}), .a ({new_AGEMA_signal_6569, new_AGEMA_signal_6565}), .c ({new_AGEMA_signal_3662, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3712, RoundKeyOutput[113]}), .a ({new_AGEMA_signal_6577, new_AGEMA_signal_6573}), .c ({new_AGEMA_signal_3787, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3713, RoundKeyOutput[114]}), .a ({new_AGEMA_signal_6585, new_AGEMA_signal_6581}), .c ({new_AGEMA_signal_3789, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3714, RoundKeyOutput[115]}), .a ({new_AGEMA_signal_6593, new_AGEMA_signal_6589}), .c ({new_AGEMA_signal_3791, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3715, RoundKeyOutput[116]}), .a ({new_AGEMA_signal_6601, new_AGEMA_signal_6597}), .c ({new_AGEMA_signal_3793, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3716, RoundKeyOutput[117]}), .a ({new_AGEMA_signal_6609, new_AGEMA_signal_6605}), .c ({new_AGEMA_signal_3795, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3717, RoundKeyOutput[118]}), .a ({new_AGEMA_signal_6617, new_AGEMA_signal_6613}), .c ({new_AGEMA_signal_3797, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3718, RoundKeyOutput[119]}), .a ({new_AGEMA_signal_6625, new_AGEMA_signal_6621}), .c ({new_AGEMA_signal_3799, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3719, RoundKeyOutput[120]}), .a ({new_AGEMA_signal_6633, new_AGEMA_signal_6629}), .c ({new_AGEMA_signal_3801, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3859, RoundKeyOutput[121]}), .a ({new_AGEMA_signal_6641, new_AGEMA_signal_6637}), .c ({new_AGEMA_signal_3949, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3860, RoundKeyOutput[122]}), .a ({new_AGEMA_signal_6649, new_AGEMA_signal_6645}), .c ({new_AGEMA_signal_3951, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3861, RoundKeyOutput[123]}), .a ({new_AGEMA_signal_6657, new_AGEMA_signal_6653}), .c ({new_AGEMA_signal_3953, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3862, RoundKeyOutput[124]}), .a ({new_AGEMA_signal_6665, new_AGEMA_signal_6661}), .c ({new_AGEMA_signal_3955, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3863, RoundKeyOutput[125]}), .a ({new_AGEMA_signal_6673, new_AGEMA_signal_6669}), .c ({new_AGEMA_signal_3957, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3864, RoundKeyOutput[126]}), .a ({new_AGEMA_signal_6681, new_AGEMA_signal_6677}), .c ({new_AGEMA_signal_3959, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (new_AGEMA_signal_4681), .b ({new_AGEMA_signal_3865, RoundKeyOutput[127]}), .a ({new_AGEMA_signal_6689, new_AGEMA_signal_6685}), .c ({new_AGEMA_signal_3961, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_6697, new_AGEMA_signal_6693}), .b ({new_AGEMA_signal_3803, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_3962, KeyExpansionOutput[9]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_6705, new_AGEMA_signal_6701}), .b ({new_AGEMA_signal_3664, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_3802, KeyExpansionOutput[8]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_6713, new_AGEMA_signal_6709}), .b ({new_AGEMA_signal_3804, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_3963, KeyExpansionOutput[7]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_6721, new_AGEMA_signal_6717}), .b ({new_AGEMA_signal_3805, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_3964, KeyExpansionOutput[6]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_6729, new_AGEMA_signal_6725}), .b ({new_AGEMA_signal_3806, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_3965, KeyExpansionOutput[5]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_6737, new_AGEMA_signal_6733}), .b ({new_AGEMA_signal_3807, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_3966, KeyExpansionOutput[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_6745, new_AGEMA_signal_6741}), .b ({new_AGEMA_signal_3663, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_3803, KeyExpansionOutput[41]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6749}), .b ({new_AGEMA_signal_3609, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_3663, KeyExpansionOutput[73]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_6761, new_AGEMA_signal_6757}), .b ({new_AGEMA_signal_3590, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_3664, KeyExpansionOutput[40]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_6769, new_AGEMA_signal_6765}), .b ({new_AGEMA_signal_3555, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_3590, KeyExpansionOutput[72]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_6777, new_AGEMA_signal_6773}), .b ({new_AGEMA_signal_3808, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_3967, KeyExpansionOutput[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_6785, new_AGEMA_signal_6781}), .b ({new_AGEMA_signal_3665, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_3804, KeyExpansionOutput[39]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_6793, new_AGEMA_signal_6789}), .b ({new_AGEMA_signal_3610, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_3665, KeyExpansionOutput[71]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_6801, new_AGEMA_signal_6797}), .b ({new_AGEMA_signal_3666, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_3805, KeyExpansionOutput[38]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_6809, new_AGEMA_signal_6805}), .b ({new_AGEMA_signal_3611, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_3666, KeyExpansionOutput[70]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_6817, new_AGEMA_signal_6813}), .b ({new_AGEMA_signal_3667, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_3806, KeyExpansionOutput[37]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_6825, new_AGEMA_signal_6821}), .b ({new_AGEMA_signal_3612, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_3667, KeyExpansionOutput[69]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_6833, new_AGEMA_signal_6829}), .b ({new_AGEMA_signal_3668, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_3807, KeyExpansionOutput[36]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_6841, new_AGEMA_signal_6837}), .b ({new_AGEMA_signal_3613, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_3668, KeyExpansionOutput[68]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_6849, new_AGEMA_signal_6845}), .b ({new_AGEMA_signal_3669, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_3808, KeyExpansionOutput[35]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_6857, new_AGEMA_signal_6853}), .b ({new_AGEMA_signal_3591, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_3669, KeyExpansionOutput[67]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_6865, new_AGEMA_signal_6861}), .b ({new_AGEMA_signal_3551, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_3591, KeyExpansionOutput[99]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6869}), .b ({new_AGEMA_signal_3968, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_4119, KeyExpansionOutput[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_6881, new_AGEMA_signal_6877}), .b ({new_AGEMA_signal_3809, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_3968, KeyExpansionOutput[63]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_6889, new_AGEMA_signal_6885}), .b ({new_AGEMA_signal_3685, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_3809, KeyExpansionOutput[95]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_6897, new_AGEMA_signal_6893}), .b ({new_AGEMA_signal_3969, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_4120, KeyExpansionOutput[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_6905, new_AGEMA_signal_6901}), .b ({new_AGEMA_signal_3810, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_3969, KeyExpansionOutput[62]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_6913, new_AGEMA_signal_6909}), .b ({new_AGEMA_signal_3686, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_3810, KeyExpansionOutput[94]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_6921, new_AGEMA_signal_6917}), .b ({new_AGEMA_signal_3811, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_3970, KeyExpansionOutput[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_6929, new_AGEMA_signal_6925}), .b ({new_AGEMA_signal_3670, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_3811, KeyExpansionOutput[34]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_6937, new_AGEMA_signal_6933}), .b ({new_AGEMA_signal_3592, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_3670, KeyExpansionOutput[66]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_6945, new_AGEMA_signal_6941}), .b ({new_AGEMA_signal_3552, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_3592, KeyExpansionOutput[98]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_6953, new_AGEMA_signal_6949}), .b ({new_AGEMA_signal_3971, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_4121, KeyExpansionOutput[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_6961, new_AGEMA_signal_6957}), .b ({new_AGEMA_signal_3812, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_3971, KeyExpansionOutput[61]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_6969, new_AGEMA_signal_6965}), .b ({new_AGEMA_signal_3687, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_3812, KeyExpansionOutput[93]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_6977, new_AGEMA_signal_6973}), .b ({new_AGEMA_signal_3972, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_4122, KeyExpansionOutput[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_6985, new_AGEMA_signal_6981}), .b ({new_AGEMA_signal_3813, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_3972, KeyExpansionOutput[60]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_6993, new_AGEMA_signal_6989}), .b ({new_AGEMA_signal_3688, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_3813, KeyExpansionOutput[92]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_7001, new_AGEMA_signal_6997}), .b ({new_AGEMA_signal_3973, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_4123, KeyExpansionOutput[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_7009, new_AGEMA_signal_7005}), .b ({new_AGEMA_signal_3814, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_3973, KeyExpansionOutput[59]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_7017, new_AGEMA_signal_7013}), .b ({new_AGEMA_signal_3689, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_3814, KeyExpansionOutput[91]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_7025, new_AGEMA_signal_7021}), .b ({new_AGEMA_signal_3974, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_4124, KeyExpansionOutput[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_7033, new_AGEMA_signal_7029}), .b ({new_AGEMA_signal_3815, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_3974, KeyExpansionOutput[58]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_7041, new_AGEMA_signal_7037}), .b ({new_AGEMA_signal_3690, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_3815, KeyExpansionOutput[90]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_7049, new_AGEMA_signal_7045}), .b ({new_AGEMA_signal_3975, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_4125, KeyExpansionOutput[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_7057, new_AGEMA_signal_7053}), .b ({new_AGEMA_signal_3816, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_3975, KeyExpansionOutput[57]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_7065, new_AGEMA_signal_7061}), .b ({new_AGEMA_signal_3691, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_3816, KeyExpansionOutput[89]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_7073, new_AGEMA_signal_7069}), .b ({new_AGEMA_signal_3817, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_3976, KeyExpansionOutput[24]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_7081, new_AGEMA_signal_7077}), .b ({new_AGEMA_signal_3671, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_3817, KeyExpansionOutput[56]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_7089, new_AGEMA_signal_7085}), .b ({new_AGEMA_signal_3595, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_3671, KeyExpansionOutput[88]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_7097, new_AGEMA_signal_7093}), .b ({new_AGEMA_signal_3818, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_3977, KeyExpansionOutput[23]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_7105, new_AGEMA_signal_7101}), .b ({new_AGEMA_signal_3672, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_3818, KeyExpansionOutput[55]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_7113, new_AGEMA_signal_7109}), .b ({new_AGEMA_signal_3596, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_3672, KeyExpansionOutput[87]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_7121, new_AGEMA_signal_7117}), .b ({new_AGEMA_signal_3819, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_3978, KeyExpansionOutput[22]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_7129, new_AGEMA_signal_7125}), .b ({new_AGEMA_signal_3673, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_3819, KeyExpansionOutput[54]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_7137, new_AGEMA_signal_7133}), .b ({new_AGEMA_signal_3597, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_3673, KeyExpansionOutput[86]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_7145, new_AGEMA_signal_7141}), .b ({new_AGEMA_signal_3820, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_3979, KeyExpansionOutput[21]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_7153, new_AGEMA_signal_7149}), .b ({new_AGEMA_signal_3674, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_3820, KeyExpansionOutput[53]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_7161, new_AGEMA_signal_7157}), .b ({new_AGEMA_signal_3598, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_3674, KeyExpansionOutput[85]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_7169, new_AGEMA_signal_7165}), .b ({new_AGEMA_signal_3821, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_3980, KeyExpansionOutput[20]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_7177, new_AGEMA_signal_7173}), .b ({new_AGEMA_signal_3675, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_3821, KeyExpansionOutput[52]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_7185, new_AGEMA_signal_7181}), .b ({new_AGEMA_signal_3599, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_3675, KeyExpansionOutput[84]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_7193, new_AGEMA_signal_7189}), .b ({new_AGEMA_signal_3822, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_3981, KeyExpansionOutput[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_7201, new_AGEMA_signal_7197}), .b ({new_AGEMA_signal_3676, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_3822, KeyExpansionOutput[33]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_7209, new_AGEMA_signal_7205}), .b ({new_AGEMA_signal_3593, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_3676, KeyExpansionOutput[65]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_7217, new_AGEMA_signal_7213}), .b ({new_AGEMA_signal_3553, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_3593, KeyExpansionOutput[97]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_7225, new_AGEMA_signal_7221}), .b ({new_AGEMA_signal_3823, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_3982, KeyExpansionOutput[19]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_7233, new_AGEMA_signal_7229}), .b ({new_AGEMA_signal_3677, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_3823, KeyExpansionOutput[51]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_7241, new_AGEMA_signal_7237}), .b ({new_AGEMA_signal_3600, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_3677, KeyExpansionOutput[83]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_7249, new_AGEMA_signal_7245}), .b ({new_AGEMA_signal_3824, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_3983, KeyExpansionOutput[18]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_7257, new_AGEMA_signal_7253}), .b ({new_AGEMA_signal_3678, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_3824, KeyExpansionOutput[50]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_7265, new_AGEMA_signal_7261}), .b ({new_AGEMA_signal_3601, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_3678, KeyExpansionOutput[82]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_7273, new_AGEMA_signal_7269}), .b ({new_AGEMA_signal_3825, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_3984, KeyExpansionOutput[17]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_7281, new_AGEMA_signal_7277}), .b ({new_AGEMA_signal_3679, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_3825, KeyExpansionOutput[49]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_7289, new_AGEMA_signal_7285}), .b ({new_AGEMA_signal_3602, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_3679, KeyExpansionOutput[81]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_7297, new_AGEMA_signal_7293}), .b ({new_AGEMA_signal_3680, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_3826, KeyExpansionOutput[16]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_7305, new_AGEMA_signal_7301}), .b ({new_AGEMA_signal_3594, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_3680, KeyExpansionOutput[48]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_7313, new_AGEMA_signal_7309}), .b ({new_AGEMA_signal_3554, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_3594, KeyExpansionOutput[80]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_7321, new_AGEMA_signal_7317}), .b ({new_AGEMA_signal_3827, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_3985, KeyExpansionOutput[15]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_7329, new_AGEMA_signal_7325}), .b ({new_AGEMA_signal_3681, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_3827, KeyExpansionOutput[47]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_7337, new_AGEMA_signal_7333}), .b ({new_AGEMA_signal_3603, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_3681, KeyExpansionOutput[79]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_7345, new_AGEMA_signal_7341}), .b ({new_AGEMA_signal_3828, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_3986, KeyExpansionOutput[14]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_7353, new_AGEMA_signal_7349}), .b ({new_AGEMA_signal_3682, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_3828, KeyExpansionOutput[46]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_7361, new_AGEMA_signal_7357}), .b ({new_AGEMA_signal_3604, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_3682, KeyExpansionOutput[78]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_7369, new_AGEMA_signal_7365}), .b ({new_AGEMA_signal_3829, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_3987, KeyExpansionOutput[13]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_7377, new_AGEMA_signal_7373}), .b ({new_AGEMA_signal_3683, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_3829, KeyExpansionOutput[45]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_7385, new_AGEMA_signal_7381}), .b ({new_AGEMA_signal_3605, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_3683, KeyExpansionOutput[77]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_7393, new_AGEMA_signal_7389}), .b ({new_AGEMA_signal_3830, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_3988, KeyExpansionOutput[12]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_7401, new_AGEMA_signal_7397}), .b ({new_AGEMA_signal_3684, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_3830, KeyExpansionOutput[44]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_7409, new_AGEMA_signal_7405}), .b ({new_AGEMA_signal_3606, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_3684, KeyExpansionOutput[76]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_7417, new_AGEMA_signal_7413}), .b ({new_AGEMA_signal_3615, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_3685, KeyExpansionOutput[127]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_7425, new_AGEMA_signal_7421}), .b ({new_AGEMA_signal_3616, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_3686, KeyExpansionOutput[126]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_7433, new_AGEMA_signal_7429}), .b ({new_AGEMA_signal_3617, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_3687, KeyExpansionOutput[125]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_7441, new_AGEMA_signal_7437}), .b ({new_AGEMA_signal_3618, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_3688, KeyExpansionOutput[124]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_7449, new_AGEMA_signal_7445}), .b ({new_AGEMA_signal_3619, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_3689, KeyExpansionOutput[123]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_7457, new_AGEMA_signal_7453}), .b ({new_AGEMA_signal_3620, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_3690, KeyExpansionOutput[122]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_7465, new_AGEMA_signal_7461}), .b ({new_AGEMA_signal_3621, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_3691, KeyExpansionOutput[121]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_7473, new_AGEMA_signal_7469}), .b ({new_AGEMA_signal_3557, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_3595, KeyExpansionOutput[120]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_7481, new_AGEMA_signal_7477}), .b ({new_AGEMA_signal_3831, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_3989, KeyExpansionOutput[11]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_7489, new_AGEMA_signal_7485}), .b ({new_AGEMA_signal_3692, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_3831, KeyExpansionOutput[43]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7493}), .b ({new_AGEMA_signal_3607, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_3692, KeyExpansionOutput[75]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_7505, new_AGEMA_signal_7501}), .b ({new_AGEMA_signal_3533, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_3596, KeyExpansionOutput[119]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_7513, new_AGEMA_signal_7509}), .b ({new_AGEMA_signal_3534, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_3597, KeyExpansionOutput[118]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7517}), .b ({new_AGEMA_signal_3535, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_3598, KeyExpansionOutput[117]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_7529, new_AGEMA_signal_7525}), .b ({new_AGEMA_signal_3536, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_3599, KeyExpansionOutput[116]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_7537, new_AGEMA_signal_7533}), .b ({new_AGEMA_signal_3537, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_3600, KeyExpansionOutput[115]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_7545, new_AGEMA_signal_7541}), .b ({new_AGEMA_signal_3538, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_3601, KeyExpansionOutput[114]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_7553, new_AGEMA_signal_7549}), .b ({new_AGEMA_signal_3539, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_3602, KeyExpansionOutput[113]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_7561, new_AGEMA_signal_7557}), .b ({new_AGEMA_signal_3503, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_3554, KeyExpansionOutput[112]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_7569, new_AGEMA_signal_7565}), .b ({new_AGEMA_signal_3540, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_3603, KeyExpansionOutput[111]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_7577, new_AGEMA_signal_7573}), .b ({new_AGEMA_signal_3541, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_3604, KeyExpansionOutput[110]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_7585, new_AGEMA_signal_7581}), .b ({new_AGEMA_signal_3832, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_3990, KeyExpansionOutput[10]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_7593, new_AGEMA_signal_7589}), .b ({new_AGEMA_signal_3693, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_3832, KeyExpansionOutput[42]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_7601, new_AGEMA_signal_7597}), .b ({new_AGEMA_signal_3608, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_3693, KeyExpansionOutput[74]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_7609, new_AGEMA_signal_7605}), .b ({new_AGEMA_signal_3542, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_3605, KeyExpansionOutput[109]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_7617, new_AGEMA_signal_7613}), .b ({new_AGEMA_signal_3543, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_3606, KeyExpansionOutput[108]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_7625, new_AGEMA_signal_7621}), .b ({new_AGEMA_signal_3544, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_3607, KeyExpansionOutput[107]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_7633, new_AGEMA_signal_7629}), .b ({new_AGEMA_signal_3545, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_3608, KeyExpansionOutput[106]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7637}), .b ({new_AGEMA_signal_3546, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_3609, KeyExpansionOutput[105]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_7649, new_AGEMA_signal_7645}), .b ({new_AGEMA_signal_3514, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_3555, KeyExpansionOutput[104]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_7657, new_AGEMA_signal_7653}), .b ({new_AGEMA_signal_3547, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_3610, KeyExpansionOutput[103]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_7665, new_AGEMA_signal_7661}), .b ({new_AGEMA_signal_3548, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_3611, KeyExpansionOutput[102]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_7673, new_AGEMA_signal_7669}), .b ({new_AGEMA_signal_3549, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_3612, KeyExpansionOutput[101]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_7681, new_AGEMA_signal_7677}), .b ({new_AGEMA_signal_3550, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_3613, KeyExpansionOutput[100]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_7689, new_AGEMA_signal_7685}), .b ({new_AGEMA_signal_3694, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_3833, KeyExpansionOutput[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_7697, new_AGEMA_signal_7693}), .b ({new_AGEMA_signal_3614, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_3694, KeyExpansionOutput[32]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_7705, new_AGEMA_signal_7701}), .b ({new_AGEMA_signal_3556, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_3614, KeyExpansionOutput[64]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_7713, new_AGEMA_signal_7709}), .b ({new_AGEMA_signal_3525, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_3556, KeyExpansionOutput[96]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({1'b0, new_AGEMA_signal_7717}), .b ({new_AGEMA_signal_3526, MixColumnsIns_DoubleBytes[0]}), .c ({new_AGEMA_signal_3615, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({1'b0, new_AGEMA_signal_7721}), .b ({new_AGEMA_signal_3527, MixColumnsIns_DoubleBytes[7]}), .c ({new_AGEMA_signal_3616, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({1'b0, new_AGEMA_signal_7725}), .b ({new_AGEMA_signal_3528, MixColumnsIns_DoubleBytes[6]}), .c ({new_AGEMA_signal_3617, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({1'b0, new_AGEMA_signal_7729}), .b ({new_AGEMA_signal_3529, MixColumnsIns_DoubleBytes[5]}), .c ({new_AGEMA_signal_3618, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({1'b0, new_AGEMA_signal_7733}), .b ({new_AGEMA_signal_3530, SubBytesOutput[3]}), .c ({new_AGEMA_signal_3619, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({1'b0, new_AGEMA_signal_7737}), .b ({new_AGEMA_signal_3531, SubBytesOutput[2]}), .c ({new_AGEMA_signal_3620, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({1'b0, new_AGEMA_signal_7741}), .b ({new_AGEMA_signal_3532, MixColumnsIns_DoubleBytes[2]}), .c ({new_AGEMA_signal_3621, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({1'b0, new_AGEMA_signal_7745}), .b ({new_AGEMA_signal_3492, SubBytesOutput[0]}), .c ({new_AGEMA_signal_3557, KeyExpansionIns_tmp[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_0_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7689, new_AGEMA_signal_7685}), .a ({new_AGEMA_signal_3833, KeyExpansionOutput[0]}), .c ({new_AGEMA_signal_3991, RoundKeyOutput[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_1_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7193, new_AGEMA_signal_7189}), .a ({new_AGEMA_signal_3981, KeyExpansionOutput[1]}), .c ({new_AGEMA_signal_4126, RoundKeyOutput[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_2_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6917}), .a ({new_AGEMA_signal_3970, KeyExpansionOutput[2]}), .c ({new_AGEMA_signal_4127, RoundKeyOutput[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_3_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6777, new_AGEMA_signal_6773}), .a ({new_AGEMA_signal_3967, KeyExpansionOutput[3]}), .c ({new_AGEMA_signal_4128, RoundKeyOutput[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_4_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6737, new_AGEMA_signal_6733}), .a ({new_AGEMA_signal_3966, KeyExpansionOutput[4]}), .c ({new_AGEMA_signal_4129, RoundKeyOutput[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_5_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_6729, new_AGEMA_signal_6725}), .a ({new_AGEMA_signal_3965, KeyExpansionOutput[5]}), .c ({new_AGEMA_signal_4130, RoundKeyOutput[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_6_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6721, new_AGEMA_signal_6717}), .a ({new_AGEMA_signal_3964, KeyExpansionOutput[6]}), .c ({new_AGEMA_signal_4131, RoundKeyOutput[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_7_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6713, new_AGEMA_signal_6709}), .a ({new_AGEMA_signal_3963, KeyExpansionOutput[7]}), .c ({new_AGEMA_signal_4132, RoundKeyOutput[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_8_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_6705, new_AGEMA_signal_6701}), .a ({new_AGEMA_signal_3802, KeyExpansionOutput[8]}), .c ({new_AGEMA_signal_3992, RoundKeyOutput[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_9_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6697, new_AGEMA_signal_6693}), .a ({new_AGEMA_signal_3962, KeyExpansionOutput[9]}), .c ({new_AGEMA_signal_4133, RoundKeyOutput[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_10_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7585, new_AGEMA_signal_7581}), .a ({new_AGEMA_signal_3990, KeyExpansionOutput[10]}), .c ({new_AGEMA_signal_4134, RoundKeyOutput[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_11_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7481, new_AGEMA_signal_7477}), .a ({new_AGEMA_signal_3989, KeyExpansionOutput[11]}), .c ({new_AGEMA_signal_4135, RoundKeyOutput[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_12_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7393, new_AGEMA_signal_7389}), .a ({new_AGEMA_signal_3988, KeyExpansionOutput[12]}), .c ({new_AGEMA_signal_4136, RoundKeyOutput[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_13_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7369, new_AGEMA_signal_7365}), .a ({new_AGEMA_signal_3987, KeyExpansionOutput[13]}), .c ({new_AGEMA_signal_4137, RoundKeyOutput[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_14_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7345, new_AGEMA_signal_7341}), .a ({new_AGEMA_signal_3986, KeyExpansionOutput[14]}), .c ({new_AGEMA_signal_4138, RoundKeyOutput[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_15_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7321, new_AGEMA_signal_7317}), .a ({new_AGEMA_signal_3985, KeyExpansionOutput[15]}), .c ({new_AGEMA_signal_4139, RoundKeyOutput[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_16_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7297, new_AGEMA_signal_7293}), .a ({new_AGEMA_signal_3826, KeyExpansionOutput[16]}), .c ({new_AGEMA_signal_3993, RoundKeyOutput[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_17_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7273, new_AGEMA_signal_7269}), .a ({new_AGEMA_signal_3984, KeyExpansionOutput[17]}), .c ({new_AGEMA_signal_4140, RoundKeyOutput[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_18_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7249, new_AGEMA_signal_7245}), .a ({new_AGEMA_signal_3983, KeyExpansionOutput[18]}), .c ({new_AGEMA_signal_4141, RoundKeyOutput[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_19_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7225, new_AGEMA_signal_7221}), .a ({new_AGEMA_signal_3982, KeyExpansionOutput[19]}), .c ({new_AGEMA_signal_4142, RoundKeyOutput[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_20_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7169, new_AGEMA_signal_7165}), .a ({new_AGEMA_signal_3980, KeyExpansionOutput[20]}), .c ({new_AGEMA_signal_4143, RoundKeyOutput[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_21_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7145, new_AGEMA_signal_7141}), .a ({new_AGEMA_signal_3979, KeyExpansionOutput[21]}), .c ({new_AGEMA_signal_4144, RoundKeyOutput[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_22_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7121, new_AGEMA_signal_7117}), .a ({new_AGEMA_signal_3978, KeyExpansionOutput[22]}), .c ({new_AGEMA_signal_4145, RoundKeyOutput[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_23_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7097, new_AGEMA_signal_7093}), .a ({new_AGEMA_signal_3977, KeyExpansionOutput[23]}), .c ({new_AGEMA_signal_4146, RoundKeyOutput[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_24_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7073, new_AGEMA_signal_7069}), .a ({new_AGEMA_signal_3976, KeyExpansionOutput[24]}), .c ({new_AGEMA_signal_4147, RoundKeyOutput[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_25_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7049, new_AGEMA_signal_7045}), .a ({new_AGEMA_signal_4125, KeyExpansionOutput[25]}), .c ({new_AGEMA_signal_4265, RoundKeyOutput[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_26_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7025, new_AGEMA_signal_7021}), .a ({new_AGEMA_signal_4124, KeyExpansionOutput[26]}), .c ({new_AGEMA_signal_4266, RoundKeyOutput[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_27_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7001, new_AGEMA_signal_6997}), .a ({new_AGEMA_signal_4123, KeyExpansionOutput[27]}), .c ({new_AGEMA_signal_4267, RoundKeyOutput[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_28_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_6977, new_AGEMA_signal_6973}), .a ({new_AGEMA_signal_4122, KeyExpansionOutput[28]}), .c ({new_AGEMA_signal_4268, RoundKeyOutput[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_29_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_6953, new_AGEMA_signal_6949}), .a ({new_AGEMA_signal_4121, KeyExpansionOutput[29]}), .c ({new_AGEMA_signal_4269, RoundKeyOutput[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_30_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6897, new_AGEMA_signal_6893}), .a ({new_AGEMA_signal_4120, KeyExpansionOutput[30]}), .c ({new_AGEMA_signal_4270, RoundKeyOutput[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_31_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_6873, new_AGEMA_signal_6869}), .a ({new_AGEMA_signal_4119, KeyExpansionOutput[31]}), .c ({new_AGEMA_signal_4271, RoundKeyOutput[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_32_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7697, new_AGEMA_signal_7693}), .a ({new_AGEMA_signal_3694, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_3834, RoundKeyOutput[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_33_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7201, new_AGEMA_signal_7197}), .a ({new_AGEMA_signal_3822, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_3994, RoundKeyOutput[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_34_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6929, new_AGEMA_signal_6925}), .a ({new_AGEMA_signal_3811, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_3995, RoundKeyOutput[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_35_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6845}), .a ({new_AGEMA_signal_3808, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_3996, RoundKeyOutput[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_36_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_6833, new_AGEMA_signal_6829}), .a ({new_AGEMA_signal_3807, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_3997, RoundKeyOutput[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_37_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_6817, new_AGEMA_signal_6813}), .a ({new_AGEMA_signal_3806, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_3998, RoundKeyOutput[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_38_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6801, new_AGEMA_signal_6797}), .a ({new_AGEMA_signal_3805, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_3999, RoundKeyOutput[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_39_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_6785, new_AGEMA_signal_6781}), .a ({new_AGEMA_signal_3804, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_4000, RoundKeyOutput[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_40_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6761, new_AGEMA_signal_6757}), .a ({new_AGEMA_signal_3664, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_3835, RoundKeyOutput[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_41_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6745, new_AGEMA_signal_6741}), .a ({new_AGEMA_signal_3803, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_4001, RoundKeyOutput[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_42_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7593, new_AGEMA_signal_7589}), .a ({new_AGEMA_signal_3832, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_4002, RoundKeyOutput[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_43_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7489, new_AGEMA_signal_7485}), .a ({new_AGEMA_signal_3831, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_4003, RoundKeyOutput[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_44_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7397}), .a ({new_AGEMA_signal_3830, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_4004, RoundKeyOutput[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_45_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7373}), .a ({new_AGEMA_signal_3829, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_4005, RoundKeyOutput[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_46_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7353, new_AGEMA_signal_7349}), .a ({new_AGEMA_signal_3828, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_4006, RoundKeyOutput[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_47_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7329, new_AGEMA_signal_7325}), .a ({new_AGEMA_signal_3827, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_4007, RoundKeyOutput[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_48_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7305, new_AGEMA_signal_7301}), .a ({new_AGEMA_signal_3680, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_3836, RoundKeyOutput[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_49_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7281, new_AGEMA_signal_7277}), .a ({new_AGEMA_signal_3825, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_4008, RoundKeyOutput[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_50_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7257, new_AGEMA_signal_7253}), .a ({new_AGEMA_signal_3824, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_4009, RoundKeyOutput[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_51_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7229}), .a ({new_AGEMA_signal_3823, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_4010, RoundKeyOutput[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_52_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7177, new_AGEMA_signal_7173}), .a ({new_AGEMA_signal_3821, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_4011, RoundKeyOutput[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_53_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7153, new_AGEMA_signal_7149}), .a ({new_AGEMA_signal_3820, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_4012, RoundKeyOutput[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_54_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7129, new_AGEMA_signal_7125}), .a ({new_AGEMA_signal_3819, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_4013, RoundKeyOutput[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_55_U1 ( .s (new_AGEMA_signal_7769), .b ({new_AGEMA_signal_7105, new_AGEMA_signal_7101}), .a ({new_AGEMA_signal_3818, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_4014, RoundKeyOutput[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_56_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7081, new_AGEMA_signal_7077}), .a ({new_AGEMA_signal_3817, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_4015, RoundKeyOutput[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_57_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7057, new_AGEMA_signal_7053}), .a ({new_AGEMA_signal_3975, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_4148, RoundKeyOutput[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_58_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7033, new_AGEMA_signal_7029}), .a ({new_AGEMA_signal_3974, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_4149, RoundKeyOutput[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_59_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7009, new_AGEMA_signal_7005}), .a ({new_AGEMA_signal_3973, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_4150, RoundKeyOutput[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_60_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6985, new_AGEMA_signal_6981}), .a ({new_AGEMA_signal_3972, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_4151, RoundKeyOutput[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_61_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6961, new_AGEMA_signal_6957}), .a ({new_AGEMA_signal_3971, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_4152, RoundKeyOutput[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_62_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6905, new_AGEMA_signal_6901}), .a ({new_AGEMA_signal_3969, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_4153, RoundKeyOutput[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_63_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6881, new_AGEMA_signal_6877}), .a ({new_AGEMA_signal_3968, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_4154, RoundKeyOutput[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_64_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7705, new_AGEMA_signal_7701}), .a ({new_AGEMA_signal_3614, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_3695, RoundKeyOutput[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_65_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_7209, new_AGEMA_signal_7205}), .a ({new_AGEMA_signal_3676, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_3837, RoundKeyOutput[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_66_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6937, new_AGEMA_signal_6933}), .a ({new_AGEMA_signal_3670, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_3838, RoundKeyOutput[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_67_U1 ( .s (new_AGEMA_signal_7765), .b ({new_AGEMA_signal_6857, new_AGEMA_signal_6853}), .a ({new_AGEMA_signal_3669, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_3839, RoundKeyOutput[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_68_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6841, new_AGEMA_signal_6837}), .a ({new_AGEMA_signal_3668, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_3840, RoundKeyOutput[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_69_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6821}), .a ({new_AGEMA_signal_3667, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_3841, RoundKeyOutput[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_70_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6809, new_AGEMA_signal_6805}), .a ({new_AGEMA_signal_3666, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_3842, RoundKeyOutput[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_71_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6793, new_AGEMA_signal_6789}), .a ({new_AGEMA_signal_3665, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_3843, RoundKeyOutput[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_72_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6769, new_AGEMA_signal_6765}), .a ({new_AGEMA_signal_3590, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_3696, RoundKeyOutput[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_73_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_6753, new_AGEMA_signal_6749}), .a ({new_AGEMA_signal_3663, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_3844, RoundKeyOutput[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_74_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7601, new_AGEMA_signal_7597}), .a ({new_AGEMA_signal_3693, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_3845, RoundKeyOutput[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_75_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7493}), .a ({new_AGEMA_signal_3692, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_3846, RoundKeyOutput[75]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_76_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7409, new_AGEMA_signal_7405}), .a ({new_AGEMA_signal_3684, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_3847, RoundKeyOutput[76]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_77_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7385, new_AGEMA_signal_7381}), .a ({new_AGEMA_signal_3683, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_3848, RoundKeyOutput[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_78_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7361, new_AGEMA_signal_7357}), .a ({new_AGEMA_signal_3682, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_3849, RoundKeyOutput[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_79_U1 ( .s (new_AGEMA_signal_7761), .b ({new_AGEMA_signal_7337, new_AGEMA_signal_7333}), .a ({new_AGEMA_signal_3681, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_3850, RoundKeyOutput[79]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_80_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7313, new_AGEMA_signal_7309}), .a ({new_AGEMA_signal_3594, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_3697, RoundKeyOutput[80]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_81_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7289, new_AGEMA_signal_7285}), .a ({new_AGEMA_signal_3679, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_3851, RoundKeyOutput[81]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_82_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7265, new_AGEMA_signal_7261}), .a ({new_AGEMA_signal_3678, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_3852, RoundKeyOutput[82]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_83_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7241, new_AGEMA_signal_7237}), .a ({new_AGEMA_signal_3677, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_3853, RoundKeyOutput[83]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_84_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7185, new_AGEMA_signal_7181}), .a ({new_AGEMA_signal_3675, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_3854, RoundKeyOutput[84]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_85_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7157}), .a ({new_AGEMA_signal_3674, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_3855, RoundKeyOutput[85]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_86_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7133}), .a ({new_AGEMA_signal_3673, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_3856, RoundKeyOutput[86]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_87_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7113, new_AGEMA_signal_7109}), .a ({new_AGEMA_signal_3672, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_3857, RoundKeyOutput[87]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_88_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7085}), .a ({new_AGEMA_signal_3671, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_3858, RoundKeyOutput[88]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_89_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7061}), .a ({new_AGEMA_signal_3816, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_4016, RoundKeyOutput[89]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_90_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7041, new_AGEMA_signal_7037}), .a ({new_AGEMA_signal_3815, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_4017, RoundKeyOutput[90]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_91_U1 ( .s (new_AGEMA_signal_7757), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7013}), .a ({new_AGEMA_signal_3814, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_4018, RoundKeyOutput[91]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_92_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6993, new_AGEMA_signal_6989}), .a ({new_AGEMA_signal_3813, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_4019, RoundKeyOutput[92]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_93_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6969, new_AGEMA_signal_6965}), .a ({new_AGEMA_signal_3812, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_4020, RoundKeyOutput[93]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_94_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6913, new_AGEMA_signal_6909}), .a ({new_AGEMA_signal_3810, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_4021, RoundKeyOutput[94]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_95_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6889, new_AGEMA_signal_6885}), .a ({new_AGEMA_signal_3809, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_4022, RoundKeyOutput[95]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_96_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7713, new_AGEMA_signal_7709}), .a ({new_AGEMA_signal_3556, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_3622, RoundKeyOutput[96]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_97_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7217, new_AGEMA_signal_7213}), .a ({new_AGEMA_signal_3593, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_3698, RoundKeyOutput[97]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_98_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6945, new_AGEMA_signal_6941}), .a ({new_AGEMA_signal_3592, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_3699, RoundKeyOutput[98]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_99_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_6865, new_AGEMA_signal_6861}), .a ({new_AGEMA_signal_3591, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_3700, RoundKeyOutput[99]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_100_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7681, new_AGEMA_signal_7677}), .a ({new_AGEMA_signal_3613, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_3701, RoundKeyOutput[100]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_101_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7673, new_AGEMA_signal_7669}), .a ({new_AGEMA_signal_3612, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_3702, RoundKeyOutput[101]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_102_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7661}), .a ({new_AGEMA_signal_3611, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_3703, RoundKeyOutput[102]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_103_U1 ( .s (new_AGEMA_signal_7753), .b ({new_AGEMA_signal_7657, new_AGEMA_signal_7653}), .a ({new_AGEMA_signal_3610, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_3704, RoundKeyOutput[103]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_104_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7649, new_AGEMA_signal_7645}), .a ({new_AGEMA_signal_3555, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_3623, RoundKeyOutput[104]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_105_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7641, new_AGEMA_signal_7637}), .a ({new_AGEMA_signal_3609, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_3705, RoundKeyOutput[105]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_106_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7633, new_AGEMA_signal_7629}), .a ({new_AGEMA_signal_3608, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_3706, RoundKeyOutput[106]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_107_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7625, new_AGEMA_signal_7621}), .a ({new_AGEMA_signal_3607, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_3707, RoundKeyOutput[107]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_108_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7617, new_AGEMA_signal_7613}), .a ({new_AGEMA_signal_3606, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_3708, RoundKeyOutput[108]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_109_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7609, new_AGEMA_signal_7605}), .a ({new_AGEMA_signal_3605, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_3709, RoundKeyOutput[109]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_110_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7577, new_AGEMA_signal_7573}), .a ({new_AGEMA_signal_3604, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_3710, RoundKeyOutput[110]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_111_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7569, new_AGEMA_signal_7565}), .a ({new_AGEMA_signal_3603, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_3711, RoundKeyOutput[111]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_112_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7561, new_AGEMA_signal_7557}), .a ({new_AGEMA_signal_3554, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_3624, RoundKeyOutput[112]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_113_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7553, new_AGEMA_signal_7549}), .a ({new_AGEMA_signal_3602, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_3712, RoundKeyOutput[113]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_114_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7545, new_AGEMA_signal_7541}), .a ({new_AGEMA_signal_3601, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_3713, RoundKeyOutput[114]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_115_U1 ( .s (new_AGEMA_signal_7749), .b ({new_AGEMA_signal_7537, new_AGEMA_signal_7533}), .a ({new_AGEMA_signal_3600, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_3714, RoundKeyOutput[115]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_116_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7529, new_AGEMA_signal_7525}), .a ({new_AGEMA_signal_3599, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_3715, RoundKeyOutput[116]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_117_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7521, new_AGEMA_signal_7517}), .a ({new_AGEMA_signal_3598, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_3716, RoundKeyOutput[117]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_118_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7513, new_AGEMA_signal_7509}), .a ({new_AGEMA_signal_3597, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_3717, RoundKeyOutput[118]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_119_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7505, new_AGEMA_signal_7501}), .a ({new_AGEMA_signal_3596, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_3718, RoundKeyOutput[119]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_120_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7469}), .a ({new_AGEMA_signal_3595, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_3719, RoundKeyOutput[120]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_121_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7465, new_AGEMA_signal_7461}), .a ({new_AGEMA_signal_3691, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_3859, RoundKeyOutput[121]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_122_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7457, new_AGEMA_signal_7453}), .a ({new_AGEMA_signal_3690, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_3860, RoundKeyOutput[122]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_123_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7445}), .a ({new_AGEMA_signal_3689, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_3861, RoundKeyOutput[123]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_124_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7441, new_AGEMA_signal_7437}), .a ({new_AGEMA_signal_3688, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_3862, RoundKeyOutput[124]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_125_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7433, new_AGEMA_signal_7429}), .a ({new_AGEMA_signal_3687, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_3863, RoundKeyOutput[125]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_126_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7425, new_AGEMA_signal_7421}), .a ({new_AGEMA_signal_3686, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_3864, RoundKeyOutput[126]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MuxKeyExpansion_mux_inst_127_U1 ( .s (new_AGEMA_signal_7773), .b ({new_AGEMA_signal_7417, new_AGEMA_signal_7413}), .a ({new_AGEMA_signal_3685, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_3865, RoundKeyOutput[127]}) ) ;
    buf_clk new_AGEMA_reg_buffer_2160 ( .C (clk), .D (new_AGEMA_signal_4680), .Q (new_AGEMA_signal_4681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2164 ( .C (clk), .D (new_AGEMA_signal_4684), .Q (new_AGEMA_signal_4685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2168 ( .C (clk), .D (new_AGEMA_signal_4688), .Q (new_AGEMA_signal_4689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2172 ( .C (clk), .D (new_AGEMA_signal_4692), .Q (new_AGEMA_signal_4693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2176 ( .C (clk), .D (new_AGEMA_signal_4696), .Q (new_AGEMA_signal_4697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2180 ( .C (clk), .D (new_AGEMA_signal_4700), .Q (new_AGEMA_signal_4701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2184 ( .C (clk), .D (new_AGEMA_signal_4704), .Q (new_AGEMA_signal_4705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2188 ( .C (clk), .D (new_AGEMA_signal_4708), .Q (new_AGEMA_signal_4709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2192 ( .C (clk), .D (new_AGEMA_signal_4712), .Q (new_AGEMA_signal_4713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2196 ( .C (clk), .D (new_AGEMA_signal_4716), .Q (new_AGEMA_signal_4717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2200 ( .C (clk), .D (new_AGEMA_signal_4720), .Q (new_AGEMA_signal_4721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2204 ( .C (clk), .D (new_AGEMA_signal_4724), .Q (new_AGEMA_signal_4725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2208 ( .C (clk), .D (new_AGEMA_signal_4728), .Q (new_AGEMA_signal_4729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2212 ( .C (clk), .D (new_AGEMA_signal_4732), .Q (new_AGEMA_signal_4733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2216 ( .C (clk), .D (new_AGEMA_signal_4736), .Q (new_AGEMA_signal_4737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2220 ( .C (clk), .D (new_AGEMA_signal_4740), .Q (new_AGEMA_signal_4741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2224 ( .C (clk), .D (new_AGEMA_signal_4744), .Q (new_AGEMA_signal_4745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2228 ( .C (clk), .D (new_AGEMA_signal_4748), .Q (new_AGEMA_signal_4749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2232 ( .C (clk), .D (new_AGEMA_signal_4752), .Q (new_AGEMA_signal_4753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2236 ( .C (clk), .D (new_AGEMA_signal_4756), .Q (new_AGEMA_signal_4757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2240 ( .C (clk), .D (new_AGEMA_signal_4760), .Q (new_AGEMA_signal_4761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2244 ( .C (clk), .D (new_AGEMA_signal_4764), .Q (new_AGEMA_signal_4765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2248 ( .C (clk), .D (new_AGEMA_signal_4768), .Q (new_AGEMA_signal_4769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2252 ( .C (clk), .D (new_AGEMA_signal_4772), .Q (new_AGEMA_signal_4773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2256 ( .C (clk), .D (new_AGEMA_signal_4776), .Q (new_AGEMA_signal_4777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2260 ( .C (clk), .D (new_AGEMA_signal_4780), .Q (new_AGEMA_signal_4781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2264 ( .C (clk), .D (new_AGEMA_signal_4784), .Q (new_AGEMA_signal_4785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2268 ( .C (clk), .D (new_AGEMA_signal_4788), .Q (new_AGEMA_signal_4789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2272 ( .C (clk), .D (new_AGEMA_signal_4792), .Q (new_AGEMA_signal_4793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2276 ( .C (clk), .D (new_AGEMA_signal_4796), .Q (new_AGEMA_signal_4797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2280 ( .C (clk), .D (new_AGEMA_signal_4800), .Q (new_AGEMA_signal_4801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2284 ( .C (clk), .D (new_AGEMA_signal_4804), .Q (new_AGEMA_signal_4805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2288 ( .C (clk), .D (new_AGEMA_signal_4808), .Q (new_AGEMA_signal_4809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2292 ( .C (clk), .D (new_AGEMA_signal_4812), .Q (new_AGEMA_signal_4813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2296 ( .C (clk), .D (new_AGEMA_signal_4816), .Q (new_AGEMA_signal_4817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2300 ( .C (clk), .D (new_AGEMA_signal_4820), .Q (new_AGEMA_signal_4821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2304 ( .C (clk), .D (new_AGEMA_signal_4824), .Q (new_AGEMA_signal_4825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2308 ( .C (clk), .D (new_AGEMA_signal_4828), .Q (new_AGEMA_signal_4829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2312 ( .C (clk), .D (new_AGEMA_signal_4832), .Q (new_AGEMA_signal_4833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2316 ( .C (clk), .D (new_AGEMA_signal_4836), .Q (new_AGEMA_signal_4837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2320 ( .C (clk), .D (new_AGEMA_signal_4840), .Q (new_AGEMA_signal_4841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2324 ( .C (clk), .D (new_AGEMA_signal_4844), .Q (new_AGEMA_signal_4845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2328 ( .C (clk), .D (new_AGEMA_signal_4848), .Q (new_AGEMA_signal_4849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2332 ( .C (clk), .D (new_AGEMA_signal_4852), .Q (new_AGEMA_signal_4853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2336 ( .C (clk), .D (new_AGEMA_signal_4856), .Q (new_AGEMA_signal_4857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2340 ( .C (clk), .D (new_AGEMA_signal_4860), .Q (new_AGEMA_signal_4861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2344 ( .C (clk), .D (new_AGEMA_signal_4864), .Q (new_AGEMA_signal_4865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2348 ( .C (clk), .D (new_AGEMA_signal_4868), .Q (new_AGEMA_signal_4869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2352 ( .C (clk), .D (new_AGEMA_signal_4872), .Q (new_AGEMA_signal_4873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2356 ( .C (clk), .D (new_AGEMA_signal_4876), .Q (new_AGEMA_signal_4877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2360 ( .C (clk), .D (new_AGEMA_signal_4880), .Q (new_AGEMA_signal_4881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2364 ( .C (clk), .D (new_AGEMA_signal_4884), .Q (new_AGEMA_signal_4885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2368 ( .C (clk), .D (new_AGEMA_signal_4888), .Q (new_AGEMA_signal_4889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2372 ( .C (clk), .D (new_AGEMA_signal_4892), .Q (new_AGEMA_signal_4893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2376 ( .C (clk), .D (new_AGEMA_signal_4896), .Q (new_AGEMA_signal_4897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2380 ( .C (clk), .D (new_AGEMA_signal_4900), .Q (new_AGEMA_signal_4901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2384 ( .C (clk), .D (new_AGEMA_signal_4904), .Q (new_AGEMA_signal_4905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2388 ( .C (clk), .D (new_AGEMA_signal_4908), .Q (new_AGEMA_signal_4909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2392 ( .C (clk), .D (new_AGEMA_signal_4912), .Q (new_AGEMA_signal_4913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2396 ( .C (clk), .D (new_AGEMA_signal_4916), .Q (new_AGEMA_signal_4917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2400 ( .C (clk), .D (new_AGEMA_signal_4920), .Q (new_AGEMA_signal_4921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2404 ( .C (clk), .D (new_AGEMA_signal_4924), .Q (new_AGEMA_signal_4925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2408 ( .C (clk), .D (new_AGEMA_signal_4928), .Q (new_AGEMA_signal_4929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2412 ( .C (clk), .D (new_AGEMA_signal_4932), .Q (new_AGEMA_signal_4933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2416 ( .C (clk), .D (new_AGEMA_signal_4936), .Q (new_AGEMA_signal_4937) ) ;
    buf_clk new_AGEMA_reg_buffer_2852 ( .C (clk), .D (new_AGEMA_signal_5372), .Q (new_AGEMA_signal_5373) ) ;
    buf_clk new_AGEMA_reg_buffer_2856 ( .C (clk), .D (new_AGEMA_signal_5376), .Q (new_AGEMA_signal_5377) ) ;
    buf_clk new_AGEMA_reg_buffer_2860 ( .C (clk), .D (new_AGEMA_signal_5380), .Q (new_AGEMA_signal_5381) ) ;
    buf_clk new_AGEMA_reg_buffer_2864 ( .C (clk), .D (new_AGEMA_signal_5384), .Q (new_AGEMA_signal_5385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2868 ( .C (clk), .D (new_AGEMA_signal_5388), .Q (new_AGEMA_signal_5389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2872 ( .C (clk), .D (new_AGEMA_signal_5392), .Q (new_AGEMA_signal_5393) ) ;
    buf_clk new_AGEMA_reg_buffer_2876 ( .C (clk), .D (new_AGEMA_signal_5396), .Q (new_AGEMA_signal_5397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2880 ( .C (clk), .D (new_AGEMA_signal_5400), .Q (new_AGEMA_signal_5401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2884 ( .C (clk), .D (new_AGEMA_signal_5404), .Q (new_AGEMA_signal_5405) ) ;
    buf_clk new_AGEMA_reg_buffer_2888 ( .C (clk), .D (new_AGEMA_signal_5408), .Q (new_AGEMA_signal_5409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2892 ( .C (clk), .D (new_AGEMA_signal_5412), .Q (new_AGEMA_signal_5413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2896 ( .C (clk), .D (new_AGEMA_signal_5416), .Q (new_AGEMA_signal_5417) ) ;
    buf_clk new_AGEMA_reg_buffer_2900 ( .C (clk), .D (new_AGEMA_signal_5420), .Q (new_AGEMA_signal_5421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2904 ( .C (clk), .D (new_AGEMA_signal_5424), .Q (new_AGEMA_signal_5425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2908 ( .C (clk), .D (new_AGEMA_signal_5428), .Q (new_AGEMA_signal_5429) ) ;
    buf_clk new_AGEMA_reg_buffer_2912 ( .C (clk), .D (new_AGEMA_signal_5432), .Q (new_AGEMA_signal_5433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2916 ( .C (clk), .D (new_AGEMA_signal_5436), .Q (new_AGEMA_signal_5437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2920 ( .C (clk), .D (new_AGEMA_signal_5440), .Q (new_AGEMA_signal_5441) ) ;
    buf_clk new_AGEMA_reg_buffer_2924 ( .C (clk), .D (new_AGEMA_signal_5444), .Q (new_AGEMA_signal_5445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2928 ( .C (clk), .D (new_AGEMA_signal_5448), .Q (new_AGEMA_signal_5449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2932 ( .C (clk), .D (new_AGEMA_signal_5452), .Q (new_AGEMA_signal_5453) ) ;
    buf_clk new_AGEMA_reg_buffer_2936 ( .C (clk), .D (new_AGEMA_signal_5456), .Q (new_AGEMA_signal_5457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2940 ( .C (clk), .D (new_AGEMA_signal_5460), .Q (new_AGEMA_signal_5461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2944 ( .C (clk), .D (new_AGEMA_signal_5464), .Q (new_AGEMA_signal_5465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2948 ( .C (clk), .D (new_AGEMA_signal_5468), .Q (new_AGEMA_signal_5469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2952 ( .C (clk), .D (new_AGEMA_signal_5472), .Q (new_AGEMA_signal_5473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2956 ( .C (clk), .D (new_AGEMA_signal_5476), .Q (new_AGEMA_signal_5477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2960 ( .C (clk), .D (new_AGEMA_signal_5480), .Q (new_AGEMA_signal_5481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2964 ( .C (clk), .D (new_AGEMA_signal_5484), .Q (new_AGEMA_signal_5485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2968 ( .C (clk), .D (new_AGEMA_signal_5488), .Q (new_AGEMA_signal_5489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2972 ( .C (clk), .D (new_AGEMA_signal_5492), .Q (new_AGEMA_signal_5493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2976 ( .C (clk), .D (new_AGEMA_signal_5496), .Q (new_AGEMA_signal_5497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2980 ( .C (clk), .D (new_AGEMA_signal_5500), .Q (new_AGEMA_signal_5501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2984 ( .C (clk), .D (new_AGEMA_signal_5504), .Q (new_AGEMA_signal_5505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2988 ( .C (clk), .D (new_AGEMA_signal_5508), .Q (new_AGEMA_signal_5509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2992 ( .C (clk), .D (new_AGEMA_signal_5512), .Q (new_AGEMA_signal_5513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_2996 ( .C (clk), .D (new_AGEMA_signal_5516), .Q (new_AGEMA_signal_5517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3000 ( .C (clk), .D (new_AGEMA_signal_5520), .Q (new_AGEMA_signal_5521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3004 ( .C (clk), .D (new_AGEMA_signal_5524), .Q (new_AGEMA_signal_5525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3008 ( .C (clk), .D (new_AGEMA_signal_5528), .Q (new_AGEMA_signal_5529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3012 ( .C (clk), .D (new_AGEMA_signal_5532), .Q (new_AGEMA_signal_5533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3016 ( .C (clk), .D (new_AGEMA_signal_5536), .Q (new_AGEMA_signal_5537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3020 ( .C (clk), .D (new_AGEMA_signal_5540), .Q (new_AGEMA_signal_5541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3024 ( .C (clk), .D (new_AGEMA_signal_5544), .Q (new_AGEMA_signal_5545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3028 ( .C (clk), .D (new_AGEMA_signal_5548), .Q (new_AGEMA_signal_5549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3032 ( .C (clk), .D (new_AGEMA_signal_5552), .Q (new_AGEMA_signal_5553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3036 ( .C (clk), .D (new_AGEMA_signal_5556), .Q (new_AGEMA_signal_5557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3040 ( .C (clk), .D (new_AGEMA_signal_5560), .Q (new_AGEMA_signal_5561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3044 ( .C (clk), .D (new_AGEMA_signal_5564), .Q (new_AGEMA_signal_5565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3048 ( .C (clk), .D (new_AGEMA_signal_5568), .Q (new_AGEMA_signal_5569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3052 ( .C (clk), .D (new_AGEMA_signal_5572), .Q (new_AGEMA_signal_5573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3056 ( .C (clk), .D (new_AGEMA_signal_5576), .Q (new_AGEMA_signal_5577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3060 ( .C (clk), .D (new_AGEMA_signal_5580), .Q (new_AGEMA_signal_5581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3064 ( .C (clk), .D (new_AGEMA_signal_5584), .Q (new_AGEMA_signal_5585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3068 ( .C (clk), .D (new_AGEMA_signal_5588), .Q (new_AGEMA_signal_5589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3072 ( .C (clk), .D (new_AGEMA_signal_5592), .Q (new_AGEMA_signal_5593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3076 ( .C (clk), .D (new_AGEMA_signal_5596), .Q (new_AGEMA_signal_5597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3080 ( .C (clk), .D (new_AGEMA_signal_5600), .Q (new_AGEMA_signal_5601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3084 ( .C (clk), .D (new_AGEMA_signal_5604), .Q (new_AGEMA_signal_5605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3088 ( .C (clk), .D (new_AGEMA_signal_5608), .Q (new_AGEMA_signal_5609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3092 ( .C (clk), .D (new_AGEMA_signal_5612), .Q (new_AGEMA_signal_5613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3096 ( .C (clk), .D (new_AGEMA_signal_5616), .Q (new_AGEMA_signal_5617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3100 ( .C (clk), .D (new_AGEMA_signal_5620), .Q (new_AGEMA_signal_5621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3104 ( .C (clk), .D (new_AGEMA_signal_5624), .Q (new_AGEMA_signal_5625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3108 ( .C (clk), .D (new_AGEMA_signal_5628), .Q (new_AGEMA_signal_5629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3112 ( .C (clk), .D (new_AGEMA_signal_5632), .Q (new_AGEMA_signal_5633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3116 ( .C (clk), .D (new_AGEMA_signal_5636), .Q (new_AGEMA_signal_5637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3120 ( .C (clk), .D (new_AGEMA_signal_5640), .Q (new_AGEMA_signal_5641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3124 ( .C (clk), .D (new_AGEMA_signal_5644), .Q (new_AGEMA_signal_5645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3128 ( .C (clk), .D (new_AGEMA_signal_5648), .Q (new_AGEMA_signal_5649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3132 ( .C (clk), .D (new_AGEMA_signal_5652), .Q (new_AGEMA_signal_5653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3136 ( .C (clk), .D (new_AGEMA_signal_5656), .Q (new_AGEMA_signal_5657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3140 ( .C (clk), .D (new_AGEMA_signal_5660), .Q (new_AGEMA_signal_5661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3144 ( .C (clk), .D (new_AGEMA_signal_5664), .Q (new_AGEMA_signal_5665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3148 ( .C (clk), .D (new_AGEMA_signal_5668), .Q (new_AGEMA_signal_5669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3152 ( .C (clk), .D (new_AGEMA_signal_5672), .Q (new_AGEMA_signal_5673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3156 ( .C (clk), .D (new_AGEMA_signal_5676), .Q (new_AGEMA_signal_5677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3160 ( .C (clk), .D (new_AGEMA_signal_5680), .Q (new_AGEMA_signal_5681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3164 ( .C (clk), .D (new_AGEMA_signal_5684), .Q (new_AGEMA_signal_5685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3168 ( .C (clk), .D (new_AGEMA_signal_5688), .Q (new_AGEMA_signal_5689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3172 ( .C (clk), .D (new_AGEMA_signal_5692), .Q (new_AGEMA_signal_5693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3176 ( .C (clk), .D (new_AGEMA_signal_5696), .Q (new_AGEMA_signal_5697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3180 ( .C (clk), .D (new_AGEMA_signal_5700), .Q (new_AGEMA_signal_5701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3184 ( .C (clk), .D (new_AGEMA_signal_5704), .Q (new_AGEMA_signal_5705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3188 ( .C (clk), .D (new_AGEMA_signal_5708), .Q (new_AGEMA_signal_5709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3192 ( .C (clk), .D (new_AGEMA_signal_5712), .Q (new_AGEMA_signal_5713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3196 ( .C (clk), .D (new_AGEMA_signal_5716), .Q (new_AGEMA_signal_5717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3200 ( .C (clk), .D (new_AGEMA_signal_5720), .Q (new_AGEMA_signal_5721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3204 ( .C (clk), .D (new_AGEMA_signal_5724), .Q (new_AGEMA_signal_5725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3208 ( .C (clk), .D (new_AGEMA_signal_5728), .Q (new_AGEMA_signal_5729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3212 ( .C (clk), .D (new_AGEMA_signal_5732), .Q (new_AGEMA_signal_5733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3216 ( .C (clk), .D (new_AGEMA_signal_5736), .Q (new_AGEMA_signal_5737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3220 ( .C (clk), .D (new_AGEMA_signal_5740), .Q (new_AGEMA_signal_5741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3224 ( .C (clk), .D (new_AGEMA_signal_5744), .Q (new_AGEMA_signal_5745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3228 ( .C (clk), .D (new_AGEMA_signal_5748), .Q (new_AGEMA_signal_5749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3232 ( .C (clk), .D (new_AGEMA_signal_5752), .Q (new_AGEMA_signal_5753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3236 ( .C (clk), .D (new_AGEMA_signal_5756), .Q (new_AGEMA_signal_5757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3240 ( .C (clk), .D (new_AGEMA_signal_5760), .Q (new_AGEMA_signal_5761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3244 ( .C (clk), .D (new_AGEMA_signal_5764), .Q (new_AGEMA_signal_5765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3248 ( .C (clk), .D (new_AGEMA_signal_5768), .Q (new_AGEMA_signal_5769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3252 ( .C (clk), .D (new_AGEMA_signal_5772), .Q (new_AGEMA_signal_5773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3256 ( .C (clk), .D (new_AGEMA_signal_5776), .Q (new_AGEMA_signal_5777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3260 ( .C (clk), .D (new_AGEMA_signal_5780), .Q (new_AGEMA_signal_5781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3264 ( .C (clk), .D (new_AGEMA_signal_5784), .Q (new_AGEMA_signal_5785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3268 ( .C (clk), .D (new_AGEMA_signal_5788), .Q (new_AGEMA_signal_5789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3272 ( .C (clk), .D (new_AGEMA_signal_5792), .Q (new_AGEMA_signal_5793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3276 ( .C (clk), .D (new_AGEMA_signal_5796), .Q (new_AGEMA_signal_5797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3280 ( .C (clk), .D (new_AGEMA_signal_5800), .Q (new_AGEMA_signal_5801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3284 ( .C (clk), .D (new_AGEMA_signal_5804), .Q (new_AGEMA_signal_5805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3288 ( .C (clk), .D (new_AGEMA_signal_5808), .Q (new_AGEMA_signal_5809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3292 ( .C (clk), .D (new_AGEMA_signal_5812), .Q (new_AGEMA_signal_5813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3296 ( .C (clk), .D (new_AGEMA_signal_5816), .Q (new_AGEMA_signal_5817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3300 ( .C (clk), .D (new_AGEMA_signal_5820), .Q (new_AGEMA_signal_5821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3304 ( .C (clk), .D (new_AGEMA_signal_5824), .Q (new_AGEMA_signal_5825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3308 ( .C (clk), .D (new_AGEMA_signal_5828), .Q (new_AGEMA_signal_5829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3312 ( .C (clk), .D (new_AGEMA_signal_5832), .Q (new_AGEMA_signal_5833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3316 ( .C (clk), .D (new_AGEMA_signal_5836), .Q (new_AGEMA_signal_5837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3320 ( .C (clk), .D (new_AGEMA_signal_5840), .Q (new_AGEMA_signal_5841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3324 ( .C (clk), .D (new_AGEMA_signal_5844), .Q (new_AGEMA_signal_5845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3328 ( .C (clk), .D (new_AGEMA_signal_5848), .Q (new_AGEMA_signal_5849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3332 ( .C (clk), .D (new_AGEMA_signal_5852), .Q (new_AGEMA_signal_5853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3336 ( .C (clk), .D (new_AGEMA_signal_5856), .Q (new_AGEMA_signal_5857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3340 ( .C (clk), .D (new_AGEMA_signal_5860), .Q (new_AGEMA_signal_5861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3344 ( .C (clk), .D (new_AGEMA_signal_5864), .Q (new_AGEMA_signal_5865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3348 ( .C (clk), .D (new_AGEMA_signal_5868), .Q (new_AGEMA_signal_5869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3352 ( .C (clk), .D (new_AGEMA_signal_5872), .Q (new_AGEMA_signal_5873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3356 ( .C (clk), .D (new_AGEMA_signal_5876), .Q (new_AGEMA_signal_5877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3360 ( .C (clk), .D (new_AGEMA_signal_5880), .Q (new_AGEMA_signal_5881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3364 ( .C (clk), .D (new_AGEMA_signal_5884), .Q (new_AGEMA_signal_5885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3368 ( .C (clk), .D (new_AGEMA_signal_5888), .Q (new_AGEMA_signal_5889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3372 ( .C (clk), .D (new_AGEMA_signal_5892), .Q (new_AGEMA_signal_5893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3376 ( .C (clk), .D (new_AGEMA_signal_5896), .Q (new_AGEMA_signal_5897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3380 ( .C (clk), .D (new_AGEMA_signal_5900), .Q (new_AGEMA_signal_5901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3384 ( .C (clk), .D (new_AGEMA_signal_5904), .Q (new_AGEMA_signal_5905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3388 ( .C (clk), .D (new_AGEMA_signal_5908), .Q (new_AGEMA_signal_5909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3392 ( .C (clk), .D (new_AGEMA_signal_5912), .Q (new_AGEMA_signal_5913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3396 ( .C (clk), .D (new_AGEMA_signal_5916), .Q (new_AGEMA_signal_5917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3400 ( .C (clk), .D (new_AGEMA_signal_5920), .Q (new_AGEMA_signal_5921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3404 ( .C (clk), .D (new_AGEMA_signal_5924), .Q (new_AGEMA_signal_5925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3408 ( .C (clk), .D (new_AGEMA_signal_5928), .Q (new_AGEMA_signal_5929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3412 ( .C (clk), .D (new_AGEMA_signal_5932), .Q (new_AGEMA_signal_5933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3416 ( .C (clk), .D (new_AGEMA_signal_5936), .Q (new_AGEMA_signal_5937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3420 ( .C (clk), .D (new_AGEMA_signal_5940), .Q (new_AGEMA_signal_5941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3424 ( .C (clk), .D (new_AGEMA_signal_5944), .Q (new_AGEMA_signal_5945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3428 ( .C (clk), .D (new_AGEMA_signal_5948), .Q (new_AGEMA_signal_5949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3432 ( .C (clk), .D (new_AGEMA_signal_5952), .Q (new_AGEMA_signal_5953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3436 ( .C (clk), .D (new_AGEMA_signal_5956), .Q (new_AGEMA_signal_5957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3440 ( .C (clk), .D (new_AGEMA_signal_5960), .Q (new_AGEMA_signal_5961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3444 ( .C (clk), .D (new_AGEMA_signal_5964), .Q (new_AGEMA_signal_5965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3448 ( .C (clk), .D (new_AGEMA_signal_5968), .Q (new_AGEMA_signal_5969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3452 ( .C (clk), .D (new_AGEMA_signal_5972), .Q (new_AGEMA_signal_5973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3456 ( .C (clk), .D (new_AGEMA_signal_5976), .Q (new_AGEMA_signal_5977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3460 ( .C (clk), .D (new_AGEMA_signal_5980), .Q (new_AGEMA_signal_5981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3464 ( .C (clk), .D (new_AGEMA_signal_5984), .Q (new_AGEMA_signal_5985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3468 ( .C (clk), .D (new_AGEMA_signal_5988), .Q (new_AGEMA_signal_5989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3472 ( .C (clk), .D (new_AGEMA_signal_5992), .Q (new_AGEMA_signal_5993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3476 ( .C (clk), .D (new_AGEMA_signal_5996), .Q (new_AGEMA_signal_5997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3480 ( .C (clk), .D (new_AGEMA_signal_6000), .Q (new_AGEMA_signal_6001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3484 ( .C (clk), .D (new_AGEMA_signal_6004), .Q (new_AGEMA_signal_6005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3488 ( .C (clk), .D (new_AGEMA_signal_6008), .Q (new_AGEMA_signal_6009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3492 ( .C (clk), .D (new_AGEMA_signal_6012), .Q (new_AGEMA_signal_6013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3496 ( .C (clk), .D (new_AGEMA_signal_6016), .Q (new_AGEMA_signal_6017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3500 ( .C (clk), .D (new_AGEMA_signal_6020), .Q (new_AGEMA_signal_6021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3504 ( .C (clk), .D (new_AGEMA_signal_6024), .Q (new_AGEMA_signal_6025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3508 ( .C (clk), .D (new_AGEMA_signal_6028), .Q (new_AGEMA_signal_6029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3512 ( .C (clk), .D (new_AGEMA_signal_6032), .Q (new_AGEMA_signal_6033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3516 ( .C (clk), .D (new_AGEMA_signal_6036), .Q (new_AGEMA_signal_6037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3520 ( .C (clk), .D (new_AGEMA_signal_6040), .Q (new_AGEMA_signal_6041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3524 ( .C (clk), .D (new_AGEMA_signal_6044), .Q (new_AGEMA_signal_6045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3528 ( .C (clk), .D (new_AGEMA_signal_6048), .Q (new_AGEMA_signal_6049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3532 ( .C (clk), .D (new_AGEMA_signal_6052), .Q (new_AGEMA_signal_6053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3536 ( .C (clk), .D (new_AGEMA_signal_6056), .Q (new_AGEMA_signal_6057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3540 ( .C (clk), .D (new_AGEMA_signal_6060), .Q (new_AGEMA_signal_6061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3544 ( .C (clk), .D (new_AGEMA_signal_6064), .Q (new_AGEMA_signal_6065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3548 ( .C (clk), .D (new_AGEMA_signal_6068), .Q (new_AGEMA_signal_6069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3552 ( .C (clk), .D (new_AGEMA_signal_6072), .Q (new_AGEMA_signal_6073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3556 ( .C (clk), .D (new_AGEMA_signal_6076), .Q (new_AGEMA_signal_6077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3560 ( .C (clk), .D (new_AGEMA_signal_6080), .Q (new_AGEMA_signal_6081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3564 ( .C (clk), .D (new_AGEMA_signal_6084), .Q (new_AGEMA_signal_6085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3568 ( .C (clk), .D (new_AGEMA_signal_6088), .Q (new_AGEMA_signal_6089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3572 ( .C (clk), .D (new_AGEMA_signal_6092), .Q (new_AGEMA_signal_6093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3576 ( .C (clk), .D (new_AGEMA_signal_6096), .Q (new_AGEMA_signal_6097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3580 ( .C (clk), .D (new_AGEMA_signal_6100), .Q (new_AGEMA_signal_6101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3584 ( .C (clk), .D (new_AGEMA_signal_6104), .Q (new_AGEMA_signal_6105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3588 ( .C (clk), .D (new_AGEMA_signal_6108), .Q (new_AGEMA_signal_6109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3592 ( .C (clk), .D (new_AGEMA_signal_6112), .Q (new_AGEMA_signal_6113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3596 ( .C (clk), .D (new_AGEMA_signal_6116), .Q (new_AGEMA_signal_6117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3600 ( .C (clk), .D (new_AGEMA_signal_6120), .Q (new_AGEMA_signal_6121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3604 ( .C (clk), .D (new_AGEMA_signal_6124), .Q (new_AGEMA_signal_6125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3608 ( .C (clk), .D (new_AGEMA_signal_6128), .Q (new_AGEMA_signal_6129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3612 ( .C (clk), .D (new_AGEMA_signal_6132), .Q (new_AGEMA_signal_6133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3616 ( .C (clk), .D (new_AGEMA_signal_6136), .Q (new_AGEMA_signal_6137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3620 ( .C (clk), .D (new_AGEMA_signal_6140), .Q (new_AGEMA_signal_6141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3624 ( .C (clk), .D (new_AGEMA_signal_6144), .Q (new_AGEMA_signal_6145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3628 ( .C (clk), .D (new_AGEMA_signal_6148), .Q (new_AGEMA_signal_6149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3632 ( .C (clk), .D (new_AGEMA_signal_6152), .Q (new_AGEMA_signal_6153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3636 ( .C (clk), .D (new_AGEMA_signal_6156), .Q (new_AGEMA_signal_6157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3640 ( .C (clk), .D (new_AGEMA_signal_6160), .Q (new_AGEMA_signal_6161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3644 ( .C (clk), .D (new_AGEMA_signal_6164), .Q (new_AGEMA_signal_6165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3648 ( .C (clk), .D (new_AGEMA_signal_6168), .Q (new_AGEMA_signal_6169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3652 ( .C (clk), .D (new_AGEMA_signal_6172), .Q (new_AGEMA_signal_6173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3656 ( .C (clk), .D (new_AGEMA_signal_6176), .Q (new_AGEMA_signal_6177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3660 ( .C (clk), .D (new_AGEMA_signal_6180), .Q (new_AGEMA_signal_6181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3664 ( .C (clk), .D (new_AGEMA_signal_6184), .Q (new_AGEMA_signal_6185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3668 ( .C (clk), .D (new_AGEMA_signal_6188), .Q (new_AGEMA_signal_6189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3672 ( .C (clk), .D (new_AGEMA_signal_6192), .Q (new_AGEMA_signal_6193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3676 ( .C (clk), .D (new_AGEMA_signal_6196), .Q (new_AGEMA_signal_6197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3680 ( .C (clk), .D (new_AGEMA_signal_6200), .Q (new_AGEMA_signal_6201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3684 ( .C (clk), .D (new_AGEMA_signal_6204), .Q (new_AGEMA_signal_6205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3688 ( .C (clk), .D (new_AGEMA_signal_6208), .Q (new_AGEMA_signal_6209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3692 ( .C (clk), .D (new_AGEMA_signal_6212), .Q (new_AGEMA_signal_6213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3696 ( .C (clk), .D (new_AGEMA_signal_6216), .Q (new_AGEMA_signal_6217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3700 ( .C (clk), .D (new_AGEMA_signal_6220), .Q (new_AGEMA_signal_6221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3704 ( .C (clk), .D (new_AGEMA_signal_6224), .Q (new_AGEMA_signal_6225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3708 ( .C (clk), .D (new_AGEMA_signal_6228), .Q (new_AGEMA_signal_6229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3712 ( .C (clk), .D (new_AGEMA_signal_6232), .Q (new_AGEMA_signal_6233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3716 ( .C (clk), .D (new_AGEMA_signal_6236), .Q (new_AGEMA_signal_6237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3720 ( .C (clk), .D (new_AGEMA_signal_6240), .Q (new_AGEMA_signal_6241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3724 ( .C (clk), .D (new_AGEMA_signal_6244), .Q (new_AGEMA_signal_6245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3728 ( .C (clk), .D (new_AGEMA_signal_6248), .Q (new_AGEMA_signal_6249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3732 ( .C (clk), .D (new_AGEMA_signal_6252), .Q (new_AGEMA_signal_6253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3736 ( .C (clk), .D (new_AGEMA_signal_6256), .Q (new_AGEMA_signal_6257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3740 ( .C (clk), .D (new_AGEMA_signal_6260), .Q (new_AGEMA_signal_6261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3744 ( .C (clk), .D (new_AGEMA_signal_6264), .Q (new_AGEMA_signal_6265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3748 ( .C (clk), .D (new_AGEMA_signal_6268), .Q (new_AGEMA_signal_6269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3752 ( .C (clk), .D (new_AGEMA_signal_6272), .Q (new_AGEMA_signal_6273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3756 ( .C (clk), .D (new_AGEMA_signal_6276), .Q (new_AGEMA_signal_6277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3760 ( .C (clk), .D (new_AGEMA_signal_6280), .Q (new_AGEMA_signal_6281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3764 ( .C (clk), .D (new_AGEMA_signal_6284), .Q (new_AGEMA_signal_6285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3768 ( .C (clk), .D (new_AGEMA_signal_6288), .Q (new_AGEMA_signal_6289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3772 ( .C (clk), .D (new_AGEMA_signal_6292), .Q (new_AGEMA_signal_6293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3776 ( .C (clk), .D (new_AGEMA_signal_6296), .Q (new_AGEMA_signal_6297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3780 ( .C (clk), .D (new_AGEMA_signal_6300), .Q (new_AGEMA_signal_6301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3784 ( .C (clk), .D (new_AGEMA_signal_6304), .Q (new_AGEMA_signal_6305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3788 ( .C (clk), .D (new_AGEMA_signal_6308), .Q (new_AGEMA_signal_6309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3792 ( .C (clk), .D (new_AGEMA_signal_6312), .Q (new_AGEMA_signal_6313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3796 ( .C (clk), .D (new_AGEMA_signal_6316), .Q (new_AGEMA_signal_6317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3800 ( .C (clk), .D (new_AGEMA_signal_6320), .Q (new_AGEMA_signal_6321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3804 ( .C (clk), .D (new_AGEMA_signal_6324), .Q (new_AGEMA_signal_6325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3808 ( .C (clk), .D (new_AGEMA_signal_6328), .Q (new_AGEMA_signal_6329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3812 ( .C (clk), .D (new_AGEMA_signal_6332), .Q (new_AGEMA_signal_6333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3816 ( .C (clk), .D (new_AGEMA_signal_6336), .Q (new_AGEMA_signal_6337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3820 ( .C (clk), .D (new_AGEMA_signal_6340), .Q (new_AGEMA_signal_6341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3824 ( .C (clk), .D (new_AGEMA_signal_6344), .Q (new_AGEMA_signal_6345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3828 ( .C (clk), .D (new_AGEMA_signal_6348), .Q (new_AGEMA_signal_6349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3832 ( .C (clk), .D (new_AGEMA_signal_6352), .Q (new_AGEMA_signal_6353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3836 ( .C (clk), .D (new_AGEMA_signal_6356), .Q (new_AGEMA_signal_6357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3840 ( .C (clk), .D (new_AGEMA_signal_6360), .Q (new_AGEMA_signal_6361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3844 ( .C (clk), .D (new_AGEMA_signal_6364), .Q (new_AGEMA_signal_6365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3848 ( .C (clk), .D (new_AGEMA_signal_6368), .Q (new_AGEMA_signal_6369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3852 ( .C (clk), .D (new_AGEMA_signal_6372), .Q (new_AGEMA_signal_6373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3856 ( .C (clk), .D (new_AGEMA_signal_6376), .Q (new_AGEMA_signal_6377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3860 ( .C (clk), .D (new_AGEMA_signal_6380), .Q (new_AGEMA_signal_6381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3864 ( .C (clk), .D (new_AGEMA_signal_6384), .Q (new_AGEMA_signal_6385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3868 ( .C (clk), .D (new_AGEMA_signal_6388), .Q (new_AGEMA_signal_6389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3872 ( .C (clk), .D (new_AGEMA_signal_6392), .Q (new_AGEMA_signal_6393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3876 ( .C (clk), .D (new_AGEMA_signal_6396), .Q (new_AGEMA_signal_6397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3880 ( .C (clk), .D (new_AGEMA_signal_6400), .Q (new_AGEMA_signal_6401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3884 ( .C (clk), .D (new_AGEMA_signal_6404), .Q (new_AGEMA_signal_6405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3888 ( .C (clk), .D (new_AGEMA_signal_6408), .Q (new_AGEMA_signal_6409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3892 ( .C (clk), .D (new_AGEMA_signal_6412), .Q (new_AGEMA_signal_6413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3896 ( .C (clk), .D (new_AGEMA_signal_6416), .Q (new_AGEMA_signal_6417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3900 ( .C (clk), .D (new_AGEMA_signal_6420), .Q (new_AGEMA_signal_6421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3904 ( .C (clk), .D (new_AGEMA_signal_6424), .Q (new_AGEMA_signal_6425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3908 ( .C (clk), .D (new_AGEMA_signal_6428), .Q (new_AGEMA_signal_6429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3912 ( .C (clk), .D (new_AGEMA_signal_6432), .Q (new_AGEMA_signal_6433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3916 ( .C (clk), .D (new_AGEMA_signal_6436), .Q (new_AGEMA_signal_6437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3920 ( .C (clk), .D (new_AGEMA_signal_6440), .Q (new_AGEMA_signal_6441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3924 ( .C (clk), .D (new_AGEMA_signal_6444), .Q (new_AGEMA_signal_6445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3928 ( .C (clk), .D (new_AGEMA_signal_6448), .Q (new_AGEMA_signal_6449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3932 ( .C (clk), .D (new_AGEMA_signal_6452), .Q (new_AGEMA_signal_6453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3936 ( .C (clk), .D (new_AGEMA_signal_6456), .Q (new_AGEMA_signal_6457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3940 ( .C (clk), .D (new_AGEMA_signal_6460), .Q (new_AGEMA_signal_6461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3944 ( .C (clk), .D (new_AGEMA_signal_6464), .Q (new_AGEMA_signal_6465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3948 ( .C (clk), .D (new_AGEMA_signal_6468), .Q (new_AGEMA_signal_6469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3952 ( .C (clk), .D (new_AGEMA_signal_6472), .Q (new_AGEMA_signal_6473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3956 ( .C (clk), .D (new_AGEMA_signal_6476), .Q (new_AGEMA_signal_6477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3960 ( .C (clk), .D (new_AGEMA_signal_6480), .Q (new_AGEMA_signal_6481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3964 ( .C (clk), .D (new_AGEMA_signal_6484), .Q (new_AGEMA_signal_6485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3968 ( .C (clk), .D (new_AGEMA_signal_6488), .Q (new_AGEMA_signal_6489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3972 ( .C (clk), .D (new_AGEMA_signal_6492), .Q (new_AGEMA_signal_6493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3976 ( .C (clk), .D (new_AGEMA_signal_6496), .Q (new_AGEMA_signal_6497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3980 ( .C (clk), .D (new_AGEMA_signal_6500), .Q (new_AGEMA_signal_6501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3984 ( .C (clk), .D (new_AGEMA_signal_6504), .Q (new_AGEMA_signal_6505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3988 ( .C (clk), .D (new_AGEMA_signal_6508), .Q (new_AGEMA_signal_6509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3992 ( .C (clk), .D (new_AGEMA_signal_6512), .Q (new_AGEMA_signal_6513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_3996 ( .C (clk), .D (new_AGEMA_signal_6516), .Q (new_AGEMA_signal_6517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4000 ( .C (clk), .D (new_AGEMA_signal_6520), .Q (new_AGEMA_signal_6521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4004 ( .C (clk), .D (new_AGEMA_signal_6524), .Q (new_AGEMA_signal_6525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4008 ( .C (clk), .D (new_AGEMA_signal_6528), .Q (new_AGEMA_signal_6529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4012 ( .C (clk), .D (new_AGEMA_signal_6532), .Q (new_AGEMA_signal_6533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4016 ( .C (clk), .D (new_AGEMA_signal_6536), .Q (new_AGEMA_signal_6537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4020 ( .C (clk), .D (new_AGEMA_signal_6540), .Q (new_AGEMA_signal_6541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4024 ( .C (clk), .D (new_AGEMA_signal_6544), .Q (new_AGEMA_signal_6545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4028 ( .C (clk), .D (new_AGEMA_signal_6548), .Q (new_AGEMA_signal_6549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4032 ( .C (clk), .D (new_AGEMA_signal_6552), .Q (new_AGEMA_signal_6553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4036 ( .C (clk), .D (new_AGEMA_signal_6556), .Q (new_AGEMA_signal_6557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4040 ( .C (clk), .D (new_AGEMA_signal_6560), .Q (new_AGEMA_signal_6561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4044 ( .C (clk), .D (new_AGEMA_signal_6564), .Q (new_AGEMA_signal_6565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4048 ( .C (clk), .D (new_AGEMA_signal_6568), .Q (new_AGEMA_signal_6569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4052 ( .C (clk), .D (new_AGEMA_signal_6572), .Q (new_AGEMA_signal_6573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4056 ( .C (clk), .D (new_AGEMA_signal_6576), .Q (new_AGEMA_signal_6577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4060 ( .C (clk), .D (new_AGEMA_signal_6580), .Q (new_AGEMA_signal_6581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4064 ( .C (clk), .D (new_AGEMA_signal_6584), .Q (new_AGEMA_signal_6585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4068 ( .C (clk), .D (new_AGEMA_signal_6588), .Q (new_AGEMA_signal_6589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4072 ( .C (clk), .D (new_AGEMA_signal_6592), .Q (new_AGEMA_signal_6593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4076 ( .C (clk), .D (new_AGEMA_signal_6596), .Q (new_AGEMA_signal_6597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4080 ( .C (clk), .D (new_AGEMA_signal_6600), .Q (new_AGEMA_signal_6601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4084 ( .C (clk), .D (new_AGEMA_signal_6604), .Q (new_AGEMA_signal_6605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4088 ( .C (clk), .D (new_AGEMA_signal_6608), .Q (new_AGEMA_signal_6609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4092 ( .C (clk), .D (new_AGEMA_signal_6612), .Q (new_AGEMA_signal_6613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4096 ( .C (clk), .D (new_AGEMA_signal_6616), .Q (new_AGEMA_signal_6617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4100 ( .C (clk), .D (new_AGEMA_signal_6620), .Q (new_AGEMA_signal_6621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4104 ( .C (clk), .D (new_AGEMA_signal_6624), .Q (new_AGEMA_signal_6625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4108 ( .C (clk), .D (new_AGEMA_signal_6628), .Q (new_AGEMA_signal_6629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4112 ( .C (clk), .D (new_AGEMA_signal_6632), .Q (new_AGEMA_signal_6633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4116 ( .C (clk), .D (new_AGEMA_signal_6636), .Q (new_AGEMA_signal_6637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4120 ( .C (clk), .D (new_AGEMA_signal_6640), .Q (new_AGEMA_signal_6641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4124 ( .C (clk), .D (new_AGEMA_signal_6644), .Q (new_AGEMA_signal_6645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4128 ( .C (clk), .D (new_AGEMA_signal_6648), .Q (new_AGEMA_signal_6649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4132 ( .C (clk), .D (new_AGEMA_signal_6652), .Q (new_AGEMA_signal_6653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4136 ( .C (clk), .D (new_AGEMA_signal_6656), .Q (new_AGEMA_signal_6657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4140 ( .C (clk), .D (new_AGEMA_signal_6660), .Q (new_AGEMA_signal_6661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4144 ( .C (clk), .D (new_AGEMA_signal_6664), .Q (new_AGEMA_signal_6665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4148 ( .C (clk), .D (new_AGEMA_signal_6668), .Q (new_AGEMA_signal_6669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4152 ( .C (clk), .D (new_AGEMA_signal_6672), .Q (new_AGEMA_signal_6673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4156 ( .C (clk), .D (new_AGEMA_signal_6676), .Q (new_AGEMA_signal_6677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4160 ( .C (clk), .D (new_AGEMA_signal_6680), .Q (new_AGEMA_signal_6681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4164 ( .C (clk), .D (new_AGEMA_signal_6684), .Q (new_AGEMA_signal_6685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4168 ( .C (clk), .D (new_AGEMA_signal_6688), .Q (new_AGEMA_signal_6689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4172 ( .C (clk), .D (new_AGEMA_signal_6692), .Q (new_AGEMA_signal_6693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4176 ( .C (clk), .D (new_AGEMA_signal_6696), .Q (new_AGEMA_signal_6697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4180 ( .C (clk), .D (new_AGEMA_signal_6700), .Q (new_AGEMA_signal_6701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4184 ( .C (clk), .D (new_AGEMA_signal_6704), .Q (new_AGEMA_signal_6705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4188 ( .C (clk), .D (new_AGEMA_signal_6708), .Q (new_AGEMA_signal_6709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4192 ( .C (clk), .D (new_AGEMA_signal_6712), .Q (new_AGEMA_signal_6713) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4196 ( .C (clk), .D (new_AGEMA_signal_6716), .Q (new_AGEMA_signal_6717) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4200 ( .C (clk), .D (new_AGEMA_signal_6720), .Q (new_AGEMA_signal_6721) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4204 ( .C (clk), .D (new_AGEMA_signal_6724), .Q (new_AGEMA_signal_6725) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4208 ( .C (clk), .D (new_AGEMA_signal_6728), .Q (new_AGEMA_signal_6729) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4212 ( .C (clk), .D (new_AGEMA_signal_6732), .Q (new_AGEMA_signal_6733) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4216 ( .C (clk), .D (new_AGEMA_signal_6736), .Q (new_AGEMA_signal_6737) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4220 ( .C (clk), .D (new_AGEMA_signal_6740), .Q (new_AGEMA_signal_6741) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4224 ( .C (clk), .D (new_AGEMA_signal_6744), .Q (new_AGEMA_signal_6745) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4228 ( .C (clk), .D (new_AGEMA_signal_6748), .Q (new_AGEMA_signal_6749) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4232 ( .C (clk), .D (new_AGEMA_signal_6752), .Q (new_AGEMA_signal_6753) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4236 ( .C (clk), .D (new_AGEMA_signal_6756), .Q (new_AGEMA_signal_6757) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4240 ( .C (clk), .D (new_AGEMA_signal_6760), .Q (new_AGEMA_signal_6761) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4244 ( .C (clk), .D (new_AGEMA_signal_6764), .Q (new_AGEMA_signal_6765) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4248 ( .C (clk), .D (new_AGEMA_signal_6768), .Q (new_AGEMA_signal_6769) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4252 ( .C (clk), .D (new_AGEMA_signal_6772), .Q (new_AGEMA_signal_6773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4256 ( .C (clk), .D (new_AGEMA_signal_6776), .Q (new_AGEMA_signal_6777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4260 ( .C (clk), .D (new_AGEMA_signal_6780), .Q (new_AGEMA_signal_6781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4264 ( .C (clk), .D (new_AGEMA_signal_6784), .Q (new_AGEMA_signal_6785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4268 ( .C (clk), .D (new_AGEMA_signal_6788), .Q (new_AGEMA_signal_6789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4272 ( .C (clk), .D (new_AGEMA_signal_6792), .Q (new_AGEMA_signal_6793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4276 ( .C (clk), .D (new_AGEMA_signal_6796), .Q (new_AGEMA_signal_6797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4280 ( .C (clk), .D (new_AGEMA_signal_6800), .Q (new_AGEMA_signal_6801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4284 ( .C (clk), .D (new_AGEMA_signal_6804), .Q (new_AGEMA_signal_6805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4288 ( .C (clk), .D (new_AGEMA_signal_6808), .Q (new_AGEMA_signal_6809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4292 ( .C (clk), .D (new_AGEMA_signal_6812), .Q (new_AGEMA_signal_6813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4296 ( .C (clk), .D (new_AGEMA_signal_6816), .Q (new_AGEMA_signal_6817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4300 ( .C (clk), .D (new_AGEMA_signal_6820), .Q (new_AGEMA_signal_6821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4304 ( .C (clk), .D (new_AGEMA_signal_6824), .Q (new_AGEMA_signal_6825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4308 ( .C (clk), .D (new_AGEMA_signal_6828), .Q (new_AGEMA_signal_6829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4312 ( .C (clk), .D (new_AGEMA_signal_6832), .Q (new_AGEMA_signal_6833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4316 ( .C (clk), .D (new_AGEMA_signal_6836), .Q (new_AGEMA_signal_6837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4320 ( .C (clk), .D (new_AGEMA_signal_6840), .Q (new_AGEMA_signal_6841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4324 ( .C (clk), .D (new_AGEMA_signal_6844), .Q (new_AGEMA_signal_6845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4328 ( .C (clk), .D (new_AGEMA_signal_6848), .Q (new_AGEMA_signal_6849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4332 ( .C (clk), .D (new_AGEMA_signal_6852), .Q (new_AGEMA_signal_6853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4336 ( .C (clk), .D (new_AGEMA_signal_6856), .Q (new_AGEMA_signal_6857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4340 ( .C (clk), .D (new_AGEMA_signal_6860), .Q (new_AGEMA_signal_6861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4344 ( .C (clk), .D (new_AGEMA_signal_6864), .Q (new_AGEMA_signal_6865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4348 ( .C (clk), .D (new_AGEMA_signal_6868), .Q (new_AGEMA_signal_6869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4352 ( .C (clk), .D (new_AGEMA_signal_6872), .Q (new_AGEMA_signal_6873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4356 ( .C (clk), .D (new_AGEMA_signal_6876), .Q (new_AGEMA_signal_6877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4360 ( .C (clk), .D (new_AGEMA_signal_6880), .Q (new_AGEMA_signal_6881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4364 ( .C (clk), .D (new_AGEMA_signal_6884), .Q (new_AGEMA_signal_6885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4368 ( .C (clk), .D (new_AGEMA_signal_6888), .Q (new_AGEMA_signal_6889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4372 ( .C (clk), .D (new_AGEMA_signal_6892), .Q (new_AGEMA_signal_6893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4376 ( .C (clk), .D (new_AGEMA_signal_6896), .Q (new_AGEMA_signal_6897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4380 ( .C (clk), .D (new_AGEMA_signal_6900), .Q (new_AGEMA_signal_6901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4384 ( .C (clk), .D (new_AGEMA_signal_6904), .Q (new_AGEMA_signal_6905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4388 ( .C (clk), .D (new_AGEMA_signal_6908), .Q (new_AGEMA_signal_6909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4392 ( .C (clk), .D (new_AGEMA_signal_6912), .Q (new_AGEMA_signal_6913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4396 ( .C (clk), .D (new_AGEMA_signal_6916), .Q (new_AGEMA_signal_6917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4400 ( .C (clk), .D (new_AGEMA_signal_6920), .Q (new_AGEMA_signal_6921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4404 ( .C (clk), .D (new_AGEMA_signal_6924), .Q (new_AGEMA_signal_6925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4408 ( .C (clk), .D (new_AGEMA_signal_6928), .Q (new_AGEMA_signal_6929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4412 ( .C (clk), .D (new_AGEMA_signal_6932), .Q (new_AGEMA_signal_6933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4416 ( .C (clk), .D (new_AGEMA_signal_6936), .Q (new_AGEMA_signal_6937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4420 ( .C (clk), .D (new_AGEMA_signal_6940), .Q (new_AGEMA_signal_6941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4424 ( .C (clk), .D (new_AGEMA_signal_6944), .Q (new_AGEMA_signal_6945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4428 ( .C (clk), .D (new_AGEMA_signal_6948), .Q (new_AGEMA_signal_6949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4432 ( .C (clk), .D (new_AGEMA_signal_6952), .Q (new_AGEMA_signal_6953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4436 ( .C (clk), .D (new_AGEMA_signal_6956), .Q (new_AGEMA_signal_6957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4440 ( .C (clk), .D (new_AGEMA_signal_6960), .Q (new_AGEMA_signal_6961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4444 ( .C (clk), .D (new_AGEMA_signal_6964), .Q (new_AGEMA_signal_6965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4448 ( .C (clk), .D (new_AGEMA_signal_6968), .Q (new_AGEMA_signal_6969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4452 ( .C (clk), .D (new_AGEMA_signal_6972), .Q (new_AGEMA_signal_6973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4456 ( .C (clk), .D (new_AGEMA_signal_6976), .Q (new_AGEMA_signal_6977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4460 ( .C (clk), .D (new_AGEMA_signal_6980), .Q (new_AGEMA_signal_6981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4464 ( .C (clk), .D (new_AGEMA_signal_6984), .Q (new_AGEMA_signal_6985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4468 ( .C (clk), .D (new_AGEMA_signal_6988), .Q (new_AGEMA_signal_6989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4472 ( .C (clk), .D (new_AGEMA_signal_6992), .Q (new_AGEMA_signal_6993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4476 ( .C (clk), .D (new_AGEMA_signal_6996), .Q (new_AGEMA_signal_6997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4480 ( .C (clk), .D (new_AGEMA_signal_7000), .Q (new_AGEMA_signal_7001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4484 ( .C (clk), .D (new_AGEMA_signal_7004), .Q (new_AGEMA_signal_7005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4488 ( .C (clk), .D (new_AGEMA_signal_7008), .Q (new_AGEMA_signal_7009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4492 ( .C (clk), .D (new_AGEMA_signal_7012), .Q (new_AGEMA_signal_7013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4496 ( .C (clk), .D (new_AGEMA_signal_7016), .Q (new_AGEMA_signal_7017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4500 ( .C (clk), .D (new_AGEMA_signal_7020), .Q (new_AGEMA_signal_7021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4504 ( .C (clk), .D (new_AGEMA_signal_7024), .Q (new_AGEMA_signal_7025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4508 ( .C (clk), .D (new_AGEMA_signal_7028), .Q (new_AGEMA_signal_7029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4512 ( .C (clk), .D (new_AGEMA_signal_7032), .Q (new_AGEMA_signal_7033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4516 ( .C (clk), .D (new_AGEMA_signal_7036), .Q (new_AGEMA_signal_7037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4520 ( .C (clk), .D (new_AGEMA_signal_7040), .Q (new_AGEMA_signal_7041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4524 ( .C (clk), .D (new_AGEMA_signal_7044), .Q (new_AGEMA_signal_7045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4528 ( .C (clk), .D (new_AGEMA_signal_7048), .Q (new_AGEMA_signal_7049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4532 ( .C (clk), .D (new_AGEMA_signal_7052), .Q (new_AGEMA_signal_7053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4536 ( .C (clk), .D (new_AGEMA_signal_7056), .Q (new_AGEMA_signal_7057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4540 ( .C (clk), .D (new_AGEMA_signal_7060), .Q (new_AGEMA_signal_7061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4544 ( .C (clk), .D (new_AGEMA_signal_7064), .Q (new_AGEMA_signal_7065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4548 ( .C (clk), .D (new_AGEMA_signal_7068), .Q (new_AGEMA_signal_7069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4552 ( .C (clk), .D (new_AGEMA_signal_7072), .Q (new_AGEMA_signal_7073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4556 ( .C (clk), .D (new_AGEMA_signal_7076), .Q (new_AGEMA_signal_7077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4560 ( .C (clk), .D (new_AGEMA_signal_7080), .Q (new_AGEMA_signal_7081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4564 ( .C (clk), .D (new_AGEMA_signal_7084), .Q (new_AGEMA_signal_7085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4568 ( .C (clk), .D (new_AGEMA_signal_7088), .Q (new_AGEMA_signal_7089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4572 ( .C (clk), .D (new_AGEMA_signal_7092), .Q (new_AGEMA_signal_7093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4576 ( .C (clk), .D (new_AGEMA_signal_7096), .Q (new_AGEMA_signal_7097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4580 ( .C (clk), .D (new_AGEMA_signal_7100), .Q (new_AGEMA_signal_7101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4584 ( .C (clk), .D (new_AGEMA_signal_7104), .Q (new_AGEMA_signal_7105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4588 ( .C (clk), .D (new_AGEMA_signal_7108), .Q (new_AGEMA_signal_7109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4592 ( .C (clk), .D (new_AGEMA_signal_7112), .Q (new_AGEMA_signal_7113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4596 ( .C (clk), .D (new_AGEMA_signal_7116), .Q (new_AGEMA_signal_7117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4600 ( .C (clk), .D (new_AGEMA_signal_7120), .Q (new_AGEMA_signal_7121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4604 ( .C (clk), .D (new_AGEMA_signal_7124), .Q (new_AGEMA_signal_7125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4608 ( .C (clk), .D (new_AGEMA_signal_7128), .Q (new_AGEMA_signal_7129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4612 ( .C (clk), .D (new_AGEMA_signal_7132), .Q (new_AGEMA_signal_7133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4616 ( .C (clk), .D (new_AGEMA_signal_7136), .Q (new_AGEMA_signal_7137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4620 ( .C (clk), .D (new_AGEMA_signal_7140), .Q (new_AGEMA_signal_7141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4624 ( .C (clk), .D (new_AGEMA_signal_7144), .Q (new_AGEMA_signal_7145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4628 ( .C (clk), .D (new_AGEMA_signal_7148), .Q (new_AGEMA_signal_7149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4632 ( .C (clk), .D (new_AGEMA_signal_7152), .Q (new_AGEMA_signal_7153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4636 ( .C (clk), .D (new_AGEMA_signal_7156), .Q (new_AGEMA_signal_7157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4640 ( .C (clk), .D (new_AGEMA_signal_7160), .Q (new_AGEMA_signal_7161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4644 ( .C (clk), .D (new_AGEMA_signal_7164), .Q (new_AGEMA_signal_7165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4648 ( .C (clk), .D (new_AGEMA_signal_7168), .Q (new_AGEMA_signal_7169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4652 ( .C (clk), .D (new_AGEMA_signal_7172), .Q (new_AGEMA_signal_7173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4656 ( .C (clk), .D (new_AGEMA_signal_7176), .Q (new_AGEMA_signal_7177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4660 ( .C (clk), .D (new_AGEMA_signal_7180), .Q (new_AGEMA_signal_7181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4664 ( .C (clk), .D (new_AGEMA_signal_7184), .Q (new_AGEMA_signal_7185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4668 ( .C (clk), .D (new_AGEMA_signal_7188), .Q (new_AGEMA_signal_7189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4672 ( .C (clk), .D (new_AGEMA_signal_7192), .Q (new_AGEMA_signal_7193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4676 ( .C (clk), .D (new_AGEMA_signal_7196), .Q (new_AGEMA_signal_7197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4680 ( .C (clk), .D (new_AGEMA_signal_7200), .Q (new_AGEMA_signal_7201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4684 ( .C (clk), .D (new_AGEMA_signal_7204), .Q (new_AGEMA_signal_7205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4688 ( .C (clk), .D (new_AGEMA_signal_7208), .Q (new_AGEMA_signal_7209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4692 ( .C (clk), .D (new_AGEMA_signal_7212), .Q (new_AGEMA_signal_7213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4696 ( .C (clk), .D (new_AGEMA_signal_7216), .Q (new_AGEMA_signal_7217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4700 ( .C (clk), .D (new_AGEMA_signal_7220), .Q (new_AGEMA_signal_7221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4704 ( .C (clk), .D (new_AGEMA_signal_7224), .Q (new_AGEMA_signal_7225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4708 ( .C (clk), .D (new_AGEMA_signal_7228), .Q (new_AGEMA_signal_7229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4712 ( .C (clk), .D (new_AGEMA_signal_7232), .Q (new_AGEMA_signal_7233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4716 ( .C (clk), .D (new_AGEMA_signal_7236), .Q (new_AGEMA_signal_7237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4720 ( .C (clk), .D (new_AGEMA_signal_7240), .Q (new_AGEMA_signal_7241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4724 ( .C (clk), .D (new_AGEMA_signal_7244), .Q (new_AGEMA_signal_7245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4728 ( .C (clk), .D (new_AGEMA_signal_7248), .Q (new_AGEMA_signal_7249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4732 ( .C (clk), .D (new_AGEMA_signal_7252), .Q (new_AGEMA_signal_7253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4736 ( .C (clk), .D (new_AGEMA_signal_7256), .Q (new_AGEMA_signal_7257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4740 ( .C (clk), .D (new_AGEMA_signal_7260), .Q (new_AGEMA_signal_7261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4744 ( .C (clk), .D (new_AGEMA_signal_7264), .Q (new_AGEMA_signal_7265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4748 ( .C (clk), .D (new_AGEMA_signal_7268), .Q (new_AGEMA_signal_7269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4752 ( .C (clk), .D (new_AGEMA_signal_7272), .Q (new_AGEMA_signal_7273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4756 ( .C (clk), .D (new_AGEMA_signal_7276), .Q (new_AGEMA_signal_7277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4760 ( .C (clk), .D (new_AGEMA_signal_7280), .Q (new_AGEMA_signal_7281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4764 ( .C (clk), .D (new_AGEMA_signal_7284), .Q (new_AGEMA_signal_7285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4768 ( .C (clk), .D (new_AGEMA_signal_7288), .Q (new_AGEMA_signal_7289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4772 ( .C (clk), .D (new_AGEMA_signal_7292), .Q (new_AGEMA_signal_7293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4776 ( .C (clk), .D (new_AGEMA_signal_7296), .Q (new_AGEMA_signal_7297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4780 ( .C (clk), .D (new_AGEMA_signal_7300), .Q (new_AGEMA_signal_7301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4784 ( .C (clk), .D (new_AGEMA_signal_7304), .Q (new_AGEMA_signal_7305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4788 ( .C (clk), .D (new_AGEMA_signal_7308), .Q (new_AGEMA_signal_7309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4792 ( .C (clk), .D (new_AGEMA_signal_7312), .Q (new_AGEMA_signal_7313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4796 ( .C (clk), .D (new_AGEMA_signal_7316), .Q (new_AGEMA_signal_7317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4800 ( .C (clk), .D (new_AGEMA_signal_7320), .Q (new_AGEMA_signal_7321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4804 ( .C (clk), .D (new_AGEMA_signal_7324), .Q (new_AGEMA_signal_7325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4808 ( .C (clk), .D (new_AGEMA_signal_7328), .Q (new_AGEMA_signal_7329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4812 ( .C (clk), .D (new_AGEMA_signal_7332), .Q (new_AGEMA_signal_7333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4816 ( .C (clk), .D (new_AGEMA_signal_7336), .Q (new_AGEMA_signal_7337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4820 ( .C (clk), .D (new_AGEMA_signal_7340), .Q (new_AGEMA_signal_7341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4824 ( .C (clk), .D (new_AGEMA_signal_7344), .Q (new_AGEMA_signal_7345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4828 ( .C (clk), .D (new_AGEMA_signal_7348), .Q (new_AGEMA_signal_7349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4832 ( .C (clk), .D (new_AGEMA_signal_7352), .Q (new_AGEMA_signal_7353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4836 ( .C (clk), .D (new_AGEMA_signal_7356), .Q (new_AGEMA_signal_7357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4840 ( .C (clk), .D (new_AGEMA_signal_7360), .Q (new_AGEMA_signal_7361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4844 ( .C (clk), .D (new_AGEMA_signal_7364), .Q (new_AGEMA_signal_7365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4848 ( .C (clk), .D (new_AGEMA_signal_7368), .Q (new_AGEMA_signal_7369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4852 ( .C (clk), .D (new_AGEMA_signal_7372), .Q (new_AGEMA_signal_7373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4856 ( .C (clk), .D (new_AGEMA_signal_7376), .Q (new_AGEMA_signal_7377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4860 ( .C (clk), .D (new_AGEMA_signal_7380), .Q (new_AGEMA_signal_7381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4864 ( .C (clk), .D (new_AGEMA_signal_7384), .Q (new_AGEMA_signal_7385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4868 ( .C (clk), .D (new_AGEMA_signal_7388), .Q (new_AGEMA_signal_7389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4872 ( .C (clk), .D (new_AGEMA_signal_7392), .Q (new_AGEMA_signal_7393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4876 ( .C (clk), .D (new_AGEMA_signal_7396), .Q (new_AGEMA_signal_7397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4880 ( .C (clk), .D (new_AGEMA_signal_7400), .Q (new_AGEMA_signal_7401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4884 ( .C (clk), .D (new_AGEMA_signal_7404), .Q (new_AGEMA_signal_7405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4888 ( .C (clk), .D (new_AGEMA_signal_7408), .Q (new_AGEMA_signal_7409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4892 ( .C (clk), .D (new_AGEMA_signal_7412), .Q (new_AGEMA_signal_7413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4896 ( .C (clk), .D (new_AGEMA_signal_7416), .Q (new_AGEMA_signal_7417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4900 ( .C (clk), .D (new_AGEMA_signal_7420), .Q (new_AGEMA_signal_7421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4904 ( .C (clk), .D (new_AGEMA_signal_7424), .Q (new_AGEMA_signal_7425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4908 ( .C (clk), .D (new_AGEMA_signal_7428), .Q (new_AGEMA_signal_7429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4912 ( .C (clk), .D (new_AGEMA_signal_7432), .Q (new_AGEMA_signal_7433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4916 ( .C (clk), .D (new_AGEMA_signal_7436), .Q (new_AGEMA_signal_7437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4920 ( .C (clk), .D (new_AGEMA_signal_7440), .Q (new_AGEMA_signal_7441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4924 ( .C (clk), .D (new_AGEMA_signal_7444), .Q (new_AGEMA_signal_7445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4928 ( .C (clk), .D (new_AGEMA_signal_7448), .Q (new_AGEMA_signal_7449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4932 ( .C (clk), .D (new_AGEMA_signal_7452), .Q (new_AGEMA_signal_7453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4936 ( .C (clk), .D (new_AGEMA_signal_7456), .Q (new_AGEMA_signal_7457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4940 ( .C (clk), .D (new_AGEMA_signal_7460), .Q (new_AGEMA_signal_7461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4944 ( .C (clk), .D (new_AGEMA_signal_7464), .Q (new_AGEMA_signal_7465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4948 ( .C (clk), .D (new_AGEMA_signal_7468), .Q (new_AGEMA_signal_7469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4952 ( .C (clk), .D (new_AGEMA_signal_7472), .Q (new_AGEMA_signal_7473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4956 ( .C (clk), .D (new_AGEMA_signal_7476), .Q (new_AGEMA_signal_7477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4960 ( .C (clk), .D (new_AGEMA_signal_7480), .Q (new_AGEMA_signal_7481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4964 ( .C (clk), .D (new_AGEMA_signal_7484), .Q (new_AGEMA_signal_7485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4968 ( .C (clk), .D (new_AGEMA_signal_7488), .Q (new_AGEMA_signal_7489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4972 ( .C (clk), .D (new_AGEMA_signal_7492), .Q (new_AGEMA_signal_7493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4976 ( .C (clk), .D (new_AGEMA_signal_7496), .Q (new_AGEMA_signal_7497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4980 ( .C (clk), .D (new_AGEMA_signal_7500), .Q (new_AGEMA_signal_7501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4984 ( .C (clk), .D (new_AGEMA_signal_7504), .Q (new_AGEMA_signal_7505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4988 ( .C (clk), .D (new_AGEMA_signal_7508), .Q (new_AGEMA_signal_7509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4992 ( .C (clk), .D (new_AGEMA_signal_7512), .Q (new_AGEMA_signal_7513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_4996 ( .C (clk), .D (new_AGEMA_signal_7516), .Q (new_AGEMA_signal_7517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5000 ( .C (clk), .D (new_AGEMA_signal_7520), .Q (new_AGEMA_signal_7521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5004 ( .C (clk), .D (new_AGEMA_signal_7524), .Q (new_AGEMA_signal_7525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5008 ( .C (clk), .D (new_AGEMA_signal_7528), .Q (new_AGEMA_signal_7529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5012 ( .C (clk), .D (new_AGEMA_signal_7532), .Q (new_AGEMA_signal_7533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5016 ( .C (clk), .D (new_AGEMA_signal_7536), .Q (new_AGEMA_signal_7537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5020 ( .C (clk), .D (new_AGEMA_signal_7540), .Q (new_AGEMA_signal_7541) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5024 ( .C (clk), .D (new_AGEMA_signal_7544), .Q (new_AGEMA_signal_7545) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5028 ( .C (clk), .D (new_AGEMA_signal_7548), .Q (new_AGEMA_signal_7549) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5032 ( .C (clk), .D (new_AGEMA_signal_7552), .Q (new_AGEMA_signal_7553) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5036 ( .C (clk), .D (new_AGEMA_signal_7556), .Q (new_AGEMA_signal_7557) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5040 ( .C (clk), .D (new_AGEMA_signal_7560), .Q (new_AGEMA_signal_7561) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5044 ( .C (clk), .D (new_AGEMA_signal_7564), .Q (new_AGEMA_signal_7565) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5048 ( .C (clk), .D (new_AGEMA_signal_7568), .Q (new_AGEMA_signal_7569) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5052 ( .C (clk), .D (new_AGEMA_signal_7572), .Q (new_AGEMA_signal_7573) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5056 ( .C (clk), .D (new_AGEMA_signal_7576), .Q (new_AGEMA_signal_7577) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5060 ( .C (clk), .D (new_AGEMA_signal_7580), .Q (new_AGEMA_signal_7581) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5064 ( .C (clk), .D (new_AGEMA_signal_7584), .Q (new_AGEMA_signal_7585) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5068 ( .C (clk), .D (new_AGEMA_signal_7588), .Q (new_AGEMA_signal_7589) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5072 ( .C (clk), .D (new_AGEMA_signal_7592), .Q (new_AGEMA_signal_7593) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5076 ( .C (clk), .D (new_AGEMA_signal_7596), .Q (new_AGEMA_signal_7597) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5080 ( .C (clk), .D (new_AGEMA_signal_7600), .Q (new_AGEMA_signal_7601) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5084 ( .C (clk), .D (new_AGEMA_signal_7604), .Q (new_AGEMA_signal_7605) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5088 ( .C (clk), .D (new_AGEMA_signal_7608), .Q (new_AGEMA_signal_7609) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5092 ( .C (clk), .D (new_AGEMA_signal_7612), .Q (new_AGEMA_signal_7613) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5096 ( .C (clk), .D (new_AGEMA_signal_7616), .Q (new_AGEMA_signal_7617) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5100 ( .C (clk), .D (new_AGEMA_signal_7620), .Q (new_AGEMA_signal_7621) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5104 ( .C (clk), .D (new_AGEMA_signal_7624), .Q (new_AGEMA_signal_7625) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5108 ( .C (clk), .D (new_AGEMA_signal_7628), .Q (new_AGEMA_signal_7629) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5112 ( .C (clk), .D (new_AGEMA_signal_7632), .Q (new_AGEMA_signal_7633) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5116 ( .C (clk), .D (new_AGEMA_signal_7636), .Q (new_AGEMA_signal_7637) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5120 ( .C (clk), .D (new_AGEMA_signal_7640), .Q (new_AGEMA_signal_7641) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5124 ( .C (clk), .D (new_AGEMA_signal_7644), .Q (new_AGEMA_signal_7645) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5128 ( .C (clk), .D (new_AGEMA_signal_7648), .Q (new_AGEMA_signal_7649) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5132 ( .C (clk), .D (new_AGEMA_signal_7652), .Q (new_AGEMA_signal_7653) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5136 ( .C (clk), .D (new_AGEMA_signal_7656), .Q (new_AGEMA_signal_7657) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5140 ( .C (clk), .D (new_AGEMA_signal_7660), .Q (new_AGEMA_signal_7661) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5144 ( .C (clk), .D (new_AGEMA_signal_7664), .Q (new_AGEMA_signal_7665) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5148 ( .C (clk), .D (new_AGEMA_signal_7668), .Q (new_AGEMA_signal_7669) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5152 ( .C (clk), .D (new_AGEMA_signal_7672), .Q (new_AGEMA_signal_7673) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5156 ( .C (clk), .D (new_AGEMA_signal_7676), .Q (new_AGEMA_signal_7677) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5160 ( .C (clk), .D (new_AGEMA_signal_7680), .Q (new_AGEMA_signal_7681) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5164 ( .C (clk), .D (new_AGEMA_signal_7684), .Q (new_AGEMA_signal_7685) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5168 ( .C (clk), .D (new_AGEMA_signal_7688), .Q (new_AGEMA_signal_7689) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5172 ( .C (clk), .D (new_AGEMA_signal_7692), .Q (new_AGEMA_signal_7693) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5176 ( .C (clk), .D (new_AGEMA_signal_7696), .Q (new_AGEMA_signal_7697) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5180 ( .C (clk), .D (new_AGEMA_signal_7700), .Q (new_AGEMA_signal_7701) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5184 ( .C (clk), .D (new_AGEMA_signal_7704), .Q (new_AGEMA_signal_7705) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5188 ( .C (clk), .D (new_AGEMA_signal_7708), .Q (new_AGEMA_signal_7709) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5192 ( .C (clk), .D (new_AGEMA_signal_7712), .Q (new_AGEMA_signal_7713) ) ;
    buf_clk new_AGEMA_reg_buffer_5196 ( .C (clk), .D (new_AGEMA_signal_7716), .Q (new_AGEMA_signal_7717) ) ;
    buf_clk new_AGEMA_reg_buffer_5200 ( .C (clk), .D (new_AGEMA_signal_7720), .Q (new_AGEMA_signal_7721) ) ;
    buf_clk new_AGEMA_reg_buffer_5204 ( .C (clk), .D (new_AGEMA_signal_7724), .Q (new_AGEMA_signal_7725) ) ;
    buf_clk new_AGEMA_reg_buffer_5208 ( .C (clk), .D (new_AGEMA_signal_7728), .Q (new_AGEMA_signal_7729) ) ;
    buf_clk new_AGEMA_reg_buffer_5212 ( .C (clk), .D (new_AGEMA_signal_7732), .Q (new_AGEMA_signal_7733) ) ;
    buf_clk new_AGEMA_reg_buffer_5216 ( .C (clk), .D (new_AGEMA_signal_7736), .Q (new_AGEMA_signal_7737) ) ;
    buf_clk new_AGEMA_reg_buffer_5220 ( .C (clk), .D (new_AGEMA_signal_7740), .Q (new_AGEMA_signal_7741) ) ;
    buf_clk new_AGEMA_reg_buffer_5224 ( .C (clk), .D (new_AGEMA_signal_7744), .Q (new_AGEMA_signal_7745) ) ;
    buf_clk new_AGEMA_reg_buffer_5228 ( .C (clk), .D (new_AGEMA_signal_7748), .Q (new_AGEMA_signal_7749) ) ;
    buf_clk new_AGEMA_reg_buffer_5232 ( .C (clk), .D (new_AGEMA_signal_7752), .Q (new_AGEMA_signal_7753) ) ;
    buf_clk new_AGEMA_reg_buffer_5236 ( .C (clk), .D (new_AGEMA_signal_7756), .Q (new_AGEMA_signal_7757) ) ;
    buf_clk new_AGEMA_reg_buffer_5240 ( .C (clk), .D (new_AGEMA_signal_7760), .Q (new_AGEMA_signal_7761) ) ;
    buf_clk new_AGEMA_reg_buffer_5244 ( .C (clk), .D (new_AGEMA_signal_7764), .Q (new_AGEMA_signal_7765) ) ;
    buf_clk new_AGEMA_reg_buffer_5248 ( .C (clk), .D (new_AGEMA_signal_7768), .Q (new_AGEMA_signal_7769) ) ;
    buf_clk new_AGEMA_reg_buffer_5252 ( .C (clk), .D (new_AGEMA_signal_7772), .Q (new_AGEMA_signal_7773) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5256 ( .C (clk), .D (new_AGEMA_signal_7776), .Q (new_AGEMA_signal_7777) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5260 ( .C (clk), .D (new_AGEMA_signal_7780), .Q (new_AGEMA_signal_7781) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5264 ( .C (clk), .D (new_AGEMA_signal_7784), .Q (new_AGEMA_signal_7785) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5268 ( .C (clk), .D (new_AGEMA_signal_7788), .Q (new_AGEMA_signal_7789) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5272 ( .C (clk), .D (new_AGEMA_signal_7792), .Q (new_AGEMA_signal_7793) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5276 ( .C (clk), .D (new_AGEMA_signal_7796), .Q (new_AGEMA_signal_7797) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5280 ( .C (clk), .D (new_AGEMA_signal_7800), .Q (new_AGEMA_signal_7801) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5284 ( .C (clk), .D (new_AGEMA_signal_7804), .Q (new_AGEMA_signal_7805) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5288 ( .C (clk), .D (new_AGEMA_signal_7808), .Q (new_AGEMA_signal_7809) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5292 ( .C (clk), .D (new_AGEMA_signal_7812), .Q (new_AGEMA_signal_7813) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5296 ( .C (clk), .D (new_AGEMA_signal_7816), .Q (new_AGEMA_signal_7817) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5300 ( .C (clk), .D (new_AGEMA_signal_7820), .Q (new_AGEMA_signal_7821) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5304 ( .C (clk), .D (new_AGEMA_signal_7824), .Q (new_AGEMA_signal_7825) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5308 ( .C (clk), .D (new_AGEMA_signal_7828), .Q (new_AGEMA_signal_7829) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5312 ( .C (clk), .D (new_AGEMA_signal_7832), .Q (new_AGEMA_signal_7833) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5316 ( .C (clk), .D (new_AGEMA_signal_7836), .Q (new_AGEMA_signal_7837) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5320 ( .C (clk), .D (new_AGEMA_signal_7840), .Q (new_AGEMA_signal_7841) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5324 ( .C (clk), .D (new_AGEMA_signal_7844), .Q (new_AGEMA_signal_7845) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5328 ( .C (clk), .D (new_AGEMA_signal_7848), .Q (new_AGEMA_signal_7849) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5332 ( .C (clk), .D (new_AGEMA_signal_7852), .Q (new_AGEMA_signal_7853) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5336 ( .C (clk), .D (new_AGEMA_signal_7856), .Q (new_AGEMA_signal_7857) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5340 ( .C (clk), .D (new_AGEMA_signal_7860), .Q (new_AGEMA_signal_7861) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5344 ( .C (clk), .D (new_AGEMA_signal_7864), .Q (new_AGEMA_signal_7865) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5348 ( .C (clk), .D (new_AGEMA_signal_7868), .Q (new_AGEMA_signal_7869) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5352 ( .C (clk), .D (new_AGEMA_signal_7872), .Q (new_AGEMA_signal_7873) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5356 ( .C (clk), .D (new_AGEMA_signal_7876), .Q (new_AGEMA_signal_7877) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5360 ( .C (clk), .D (new_AGEMA_signal_7880), .Q (new_AGEMA_signal_7881) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5364 ( .C (clk), .D (new_AGEMA_signal_7884), .Q (new_AGEMA_signal_7885) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5368 ( .C (clk), .D (new_AGEMA_signal_7888), .Q (new_AGEMA_signal_7889) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5372 ( .C (clk), .D (new_AGEMA_signal_7892), .Q (new_AGEMA_signal_7893) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5376 ( .C (clk), .D (new_AGEMA_signal_7896), .Q (new_AGEMA_signal_7897) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5380 ( .C (clk), .D (new_AGEMA_signal_7900), .Q (new_AGEMA_signal_7901) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5384 ( .C (clk), .D (new_AGEMA_signal_7904), .Q (new_AGEMA_signal_7905) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5388 ( .C (clk), .D (new_AGEMA_signal_7908), .Q (new_AGEMA_signal_7909) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5392 ( .C (clk), .D (new_AGEMA_signal_7912), .Q (new_AGEMA_signal_7913) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5396 ( .C (clk), .D (new_AGEMA_signal_7916), .Q (new_AGEMA_signal_7917) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5400 ( .C (clk), .D (new_AGEMA_signal_7920), .Q (new_AGEMA_signal_7921) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5404 ( .C (clk), .D (new_AGEMA_signal_7924), .Q (new_AGEMA_signal_7925) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5408 ( .C (clk), .D (new_AGEMA_signal_7928), .Q (new_AGEMA_signal_7929) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5412 ( .C (clk), .D (new_AGEMA_signal_7932), .Q (new_AGEMA_signal_7933) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5416 ( .C (clk), .D (new_AGEMA_signal_7936), .Q (new_AGEMA_signal_7937) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5420 ( .C (clk), .D (new_AGEMA_signal_7940), .Q (new_AGEMA_signal_7941) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5424 ( .C (clk), .D (new_AGEMA_signal_7944), .Q (new_AGEMA_signal_7945) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5428 ( .C (clk), .D (new_AGEMA_signal_7948), .Q (new_AGEMA_signal_7949) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5432 ( .C (clk), .D (new_AGEMA_signal_7952), .Q (new_AGEMA_signal_7953) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5436 ( .C (clk), .D (new_AGEMA_signal_7956), .Q (new_AGEMA_signal_7957) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5440 ( .C (clk), .D (new_AGEMA_signal_7960), .Q (new_AGEMA_signal_7961) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5444 ( .C (clk), .D (new_AGEMA_signal_7964), .Q (new_AGEMA_signal_7965) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5448 ( .C (clk), .D (new_AGEMA_signal_7968), .Q (new_AGEMA_signal_7969) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5452 ( .C (clk), .D (new_AGEMA_signal_7972), .Q (new_AGEMA_signal_7973) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5456 ( .C (clk), .D (new_AGEMA_signal_7976), .Q (new_AGEMA_signal_7977) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5460 ( .C (clk), .D (new_AGEMA_signal_7980), .Q (new_AGEMA_signal_7981) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5464 ( .C (clk), .D (new_AGEMA_signal_7984), .Q (new_AGEMA_signal_7985) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5468 ( .C (clk), .D (new_AGEMA_signal_7988), .Q (new_AGEMA_signal_7989) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5472 ( .C (clk), .D (new_AGEMA_signal_7992), .Q (new_AGEMA_signal_7993) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5476 ( .C (clk), .D (new_AGEMA_signal_7996), .Q (new_AGEMA_signal_7997) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5480 ( .C (clk), .D (new_AGEMA_signal_8000), .Q (new_AGEMA_signal_8001) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5484 ( .C (clk), .D (new_AGEMA_signal_8004), .Q (new_AGEMA_signal_8005) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5488 ( .C (clk), .D (new_AGEMA_signal_8008), .Q (new_AGEMA_signal_8009) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5492 ( .C (clk), .D (new_AGEMA_signal_8012), .Q (new_AGEMA_signal_8013) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5496 ( .C (clk), .D (new_AGEMA_signal_8016), .Q (new_AGEMA_signal_8017) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5500 ( .C (clk), .D (new_AGEMA_signal_8020), .Q (new_AGEMA_signal_8021) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5504 ( .C (clk), .D (new_AGEMA_signal_8024), .Q (new_AGEMA_signal_8025) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5508 ( .C (clk), .D (new_AGEMA_signal_8028), .Q (new_AGEMA_signal_8029) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5512 ( .C (clk), .D (new_AGEMA_signal_8032), .Q (new_AGEMA_signal_8033) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5516 ( .C (clk), .D (new_AGEMA_signal_8036), .Q (new_AGEMA_signal_8037) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5520 ( .C (clk), .D (new_AGEMA_signal_8040), .Q (new_AGEMA_signal_8041) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5524 ( .C (clk), .D (new_AGEMA_signal_8044), .Q (new_AGEMA_signal_8045) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5528 ( .C (clk), .D (new_AGEMA_signal_8048), .Q (new_AGEMA_signal_8049) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5532 ( .C (clk), .D (new_AGEMA_signal_8052), .Q (new_AGEMA_signal_8053) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5536 ( .C (clk), .D (new_AGEMA_signal_8056), .Q (new_AGEMA_signal_8057) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5540 ( .C (clk), .D (new_AGEMA_signal_8060), .Q (new_AGEMA_signal_8061) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5544 ( .C (clk), .D (new_AGEMA_signal_8064), .Q (new_AGEMA_signal_8065) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5548 ( .C (clk), .D (new_AGEMA_signal_8068), .Q (new_AGEMA_signal_8069) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5552 ( .C (clk), .D (new_AGEMA_signal_8072), .Q (new_AGEMA_signal_8073) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5556 ( .C (clk), .D (new_AGEMA_signal_8076), .Q (new_AGEMA_signal_8077) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5560 ( .C (clk), .D (new_AGEMA_signal_8080), .Q (new_AGEMA_signal_8081) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5564 ( .C (clk), .D (new_AGEMA_signal_8084), .Q (new_AGEMA_signal_8085) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5568 ( .C (clk), .D (new_AGEMA_signal_8088), .Q (new_AGEMA_signal_8089) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5572 ( .C (clk), .D (new_AGEMA_signal_8092), .Q (new_AGEMA_signal_8093) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5576 ( .C (clk), .D (new_AGEMA_signal_8096), .Q (new_AGEMA_signal_8097) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5580 ( .C (clk), .D (new_AGEMA_signal_8100), .Q (new_AGEMA_signal_8101) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5584 ( .C (clk), .D (new_AGEMA_signal_8104), .Q (new_AGEMA_signal_8105) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5588 ( .C (clk), .D (new_AGEMA_signal_8108), .Q (new_AGEMA_signal_8109) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5592 ( .C (clk), .D (new_AGEMA_signal_8112), .Q (new_AGEMA_signal_8113) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5596 ( .C (clk), .D (new_AGEMA_signal_8116), .Q (new_AGEMA_signal_8117) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5600 ( .C (clk), .D (new_AGEMA_signal_8120), .Q (new_AGEMA_signal_8121) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5604 ( .C (clk), .D (new_AGEMA_signal_8124), .Q (new_AGEMA_signal_8125) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5608 ( .C (clk), .D (new_AGEMA_signal_8128), .Q (new_AGEMA_signal_8129) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5612 ( .C (clk), .D (new_AGEMA_signal_8132), .Q (new_AGEMA_signal_8133) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5616 ( .C (clk), .D (new_AGEMA_signal_8136), .Q (new_AGEMA_signal_8137) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5620 ( .C (clk), .D (new_AGEMA_signal_8140), .Q (new_AGEMA_signal_8141) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5624 ( .C (clk), .D (new_AGEMA_signal_8144), .Q (new_AGEMA_signal_8145) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5628 ( .C (clk), .D (new_AGEMA_signal_8148), .Q (new_AGEMA_signal_8149) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5632 ( .C (clk), .D (new_AGEMA_signal_8152), .Q (new_AGEMA_signal_8153) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5636 ( .C (clk), .D (new_AGEMA_signal_8156), .Q (new_AGEMA_signal_8157) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5640 ( .C (clk), .D (new_AGEMA_signal_8160), .Q (new_AGEMA_signal_8161) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5644 ( .C (clk), .D (new_AGEMA_signal_8164), .Q (new_AGEMA_signal_8165) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5648 ( .C (clk), .D (new_AGEMA_signal_8168), .Q (new_AGEMA_signal_8169) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5652 ( .C (clk), .D (new_AGEMA_signal_8172), .Q (new_AGEMA_signal_8173) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5656 ( .C (clk), .D (new_AGEMA_signal_8176), .Q (new_AGEMA_signal_8177) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5660 ( .C (clk), .D (new_AGEMA_signal_8180), .Q (new_AGEMA_signal_8181) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5664 ( .C (clk), .D (new_AGEMA_signal_8184), .Q (new_AGEMA_signal_8185) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5668 ( .C (clk), .D (new_AGEMA_signal_8188), .Q (new_AGEMA_signal_8189) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5672 ( .C (clk), .D (new_AGEMA_signal_8192), .Q (new_AGEMA_signal_8193) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5676 ( .C (clk), .D (new_AGEMA_signal_8196), .Q (new_AGEMA_signal_8197) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5680 ( .C (clk), .D (new_AGEMA_signal_8200), .Q (new_AGEMA_signal_8201) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5684 ( .C (clk), .D (new_AGEMA_signal_8204), .Q (new_AGEMA_signal_8205) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5688 ( .C (clk), .D (new_AGEMA_signal_8208), .Q (new_AGEMA_signal_8209) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5692 ( .C (clk), .D (new_AGEMA_signal_8212), .Q (new_AGEMA_signal_8213) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5696 ( .C (clk), .D (new_AGEMA_signal_8216), .Q (new_AGEMA_signal_8217) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5700 ( .C (clk), .D (new_AGEMA_signal_8220), .Q (new_AGEMA_signal_8221) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5704 ( .C (clk), .D (new_AGEMA_signal_8224), .Q (new_AGEMA_signal_8225) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5708 ( .C (clk), .D (new_AGEMA_signal_8228), .Q (new_AGEMA_signal_8229) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5712 ( .C (clk), .D (new_AGEMA_signal_8232), .Q (new_AGEMA_signal_8233) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5716 ( .C (clk), .D (new_AGEMA_signal_8236), .Q (new_AGEMA_signal_8237) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5720 ( .C (clk), .D (new_AGEMA_signal_8240), .Q (new_AGEMA_signal_8241) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5724 ( .C (clk), .D (new_AGEMA_signal_8244), .Q (new_AGEMA_signal_8245) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5728 ( .C (clk), .D (new_AGEMA_signal_8248), .Q (new_AGEMA_signal_8249) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5732 ( .C (clk), .D (new_AGEMA_signal_8252), .Q (new_AGEMA_signal_8253) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5736 ( .C (clk), .D (new_AGEMA_signal_8256), .Q (new_AGEMA_signal_8257) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5740 ( .C (clk), .D (new_AGEMA_signal_8260), .Q (new_AGEMA_signal_8261) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5744 ( .C (clk), .D (new_AGEMA_signal_8264), .Q (new_AGEMA_signal_8265) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5748 ( .C (clk), .D (new_AGEMA_signal_8268), .Q (new_AGEMA_signal_8269) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5752 ( .C (clk), .D (new_AGEMA_signal_8272), .Q (new_AGEMA_signal_8273) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5756 ( .C (clk), .D (new_AGEMA_signal_8276), .Q (new_AGEMA_signal_8277) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5760 ( .C (clk), .D (new_AGEMA_signal_8280), .Q (new_AGEMA_signal_8281) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5764 ( .C (clk), .D (new_AGEMA_signal_8284), .Q (new_AGEMA_signal_8285) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5768 ( .C (clk), .D (new_AGEMA_signal_8288), .Q (new_AGEMA_signal_8289) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5772 ( .C (clk), .D (new_AGEMA_signal_8292), .Q (new_AGEMA_signal_8293) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5776 ( .C (clk), .D (new_AGEMA_signal_8296), .Q (new_AGEMA_signal_8297) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5780 ( .C (clk), .D (new_AGEMA_signal_8300), .Q (new_AGEMA_signal_8301) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5784 ( .C (clk), .D (new_AGEMA_signal_8304), .Q (new_AGEMA_signal_8305) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5788 ( .C (clk), .D (new_AGEMA_signal_8308), .Q (new_AGEMA_signal_8309) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5792 ( .C (clk), .D (new_AGEMA_signal_8312), .Q (new_AGEMA_signal_8313) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5796 ( .C (clk), .D (new_AGEMA_signal_8316), .Q (new_AGEMA_signal_8317) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5800 ( .C (clk), .D (new_AGEMA_signal_8320), .Q (new_AGEMA_signal_8321) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5804 ( .C (clk), .D (new_AGEMA_signal_8324), .Q (new_AGEMA_signal_8325) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5808 ( .C (clk), .D (new_AGEMA_signal_8328), .Q (new_AGEMA_signal_8329) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5812 ( .C (clk), .D (new_AGEMA_signal_8332), .Q (new_AGEMA_signal_8333) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5816 ( .C (clk), .D (new_AGEMA_signal_8336), .Q (new_AGEMA_signal_8337) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5820 ( .C (clk), .D (new_AGEMA_signal_8340), .Q (new_AGEMA_signal_8341) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5824 ( .C (clk), .D (new_AGEMA_signal_8344), .Q (new_AGEMA_signal_8345) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5828 ( .C (clk), .D (new_AGEMA_signal_8348), .Q (new_AGEMA_signal_8349) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5832 ( .C (clk), .D (new_AGEMA_signal_8352), .Q (new_AGEMA_signal_8353) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5836 ( .C (clk), .D (new_AGEMA_signal_8356), .Q (new_AGEMA_signal_8357) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5840 ( .C (clk), .D (new_AGEMA_signal_8360), .Q (new_AGEMA_signal_8361) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5844 ( .C (clk), .D (new_AGEMA_signal_8364), .Q (new_AGEMA_signal_8365) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5848 ( .C (clk), .D (new_AGEMA_signal_8368), .Q (new_AGEMA_signal_8369) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5852 ( .C (clk), .D (new_AGEMA_signal_8372), .Q (new_AGEMA_signal_8373) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5856 ( .C (clk), .D (new_AGEMA_signal_8376), .Q (new_AGEMA_signal_8377) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5860 ( .C (clk), .D (new_AGEMA_signal_8380), .Q (new_AGEMA_signal_8381) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5864 ( .C (clk), .D (new_AGEMA_signal_8384), .Q (new_AGEMA_signal_8385) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5868 ( .C (clk), .D (new_AGEMA_signal_8388), .Q (new_AGEMA_signal_8389) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5872 ( .C (clk), .D (new_AGEMA_signal_8392), .Q (new_AGEMA_signal_8393) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5876 ( .C (clk), .D (new_AGEMA_signal_8396), .Q (new_AGEMA_signal_8397) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5880 ( .C (clk), .D (new_AGEMA_signal_8400), .Q (new_AGEMA_signal_8401) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5884 ( .C (clk), .D (new_AGEMA_signal_8404), .Q (new_AGEMA_signal_8405) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5888 ( .C (clk), .D (new_AGEMA_signal_8408), .Q (new_AGEMA_signal_8409) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5892 ( .C (clk), .D (new_AGEMA_signal_8412), .Q (new_AGEMA_signal_8413) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5896 ( .C (clk), .D (new_AGEMA_signal_8416), .Q (new_AGEMA_signal_8417) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5900 ( .C (clk), .D (new_AGEMA_signal_8420), .Q (new_AGEMA_signal_8421) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5904 ( .C (clk), .D (new_AGEMA_signal_8424), .Q (new_AGEMA_signal_8425) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5908 ( .C (clk), .D (new_AGEMA_signal_8428), .Q (new_AGEMA_signal_8429) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5912 ( .C (clk), .D (new_AGEMA_signal_8432), .Q (new_AGEMA_signal_8433) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5916 ( .C (clk), .D (new_AGEMA_signal_8436), .Q (new_AGEMA_signal_8437) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5920 ( .C (clk), .D (new_AGEMA_signal_8440), .Q (new_AGEMA_signal_8441) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5924 ( .C (clk), .D (new_AGEMA_signal_8444), .Q (new_AGEMA_signal_8445) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5928 ( .C (clk), .D (new_AGEMA_signal_8448), .Q (new_AGEMA_signal_8449) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5932 ( .C (clk), .D (new_AGEMA_signal_8452), .Q (new_AGEMA_signal_8453) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5936 ( .C (clk), .D (new_AGEMA_signal_8456), .Q (new_AGEMA_signal_8457) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5940 ( .C (clk), .D (new_AGEMA_signal_8460), .Q (new_AGEMA_signal_8461) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5944 ( .C (clk), .D (new_AGEMA_signal_8464), .Q (new_AGEMA_signal_8465) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5948 ( .C (clk), .D (new_AGEMA_signal_8468), .Q (new_AGEMA_signal_8469) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5952 ( .C (clk), .D (new_AGEMA_signal_8472), .Q (new_AGEMA_signal_8473) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5956 ( .C (clk), .D (new_AGEMA_signal_8476), .Q (new_AGEMA_signal_8477) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5960 ( .C (clk), .D (new_AGEMA_signal_8480), .Q (new_AGEMA_signal_8481) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5964 ( .C (clk), .D (new_AGEMA_signal_8484), .Q (new_AGEMA_signal_8485) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5968 ( .C (clk), .D (new_AGEMA_signal_8488), .Q (new_AGEMA_signal_8489) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5972 ( .C (clk), .D (new_AGEMA_signal_8492), .Q (new_AGEMA_signal_8493) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5976 ( .C (clk), .D (new_AGEMA_signal_8496), .Q (new_AGEMA_signal_8497) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5980 ( .C (clk), .D (new_AGEMA_signal_8500), .Q (new_AGEMA_signal_8501) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5984 ( .C (clk), .D (new_AGEMA_signal_8504), .Q (new_AGEMA_signal_8505) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5988 ( .C (clk), .D (new_AGEMA_signal_8508), .Q (new_AGEMA_signal_8509) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5992 ( .C (clk), .D (new_AGEMA_signal_8512), .Q (new_AGEMA_signal_8513) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_5996 ( .C (clk), .D (new_AGEMA_signal_8516), .Q (new_AGEMA_signal_8517) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6000 ( .C (clk), .D (new_AGEMA_signal_8520), .Q (new_AGEMA_signal_8521) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6004 ( .C (clk), .D (new_AGEMA_signal_8524), .Q (new_AGEMA_signal_8525) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6008 ( .C (clk), .D (new_AGEMA_signal_8528), .Q (new_AGEMA_signal_8529) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6012 ( .C (clk), .D (new_AGEMA_signal_8532), .Q (new_AGEMA_signal_8533) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6016 ( .C (clk), .D (new_AGEMA_signal_8536), .Q (new_AGEMA_signal_8537) ) ;
    buf_sca_clk new_AGEMA_reg_sca_buffer_6020 ( .C (clk), .D (new_AGEMA_signal_8540), .Q (new_AGEMA_signal_8541) ) ;
    buf_clk new_AGEMA_reg_buffer_6024 ( .C (clk), .D (new_AGEMA_signal_8544), .Q (new_AGEMA_signal_8545) ) ;
    buf_clk new_AGEMA_reg_buffer_6028 ( .C (clk), .D (new_AGEMA_signal_8548), .Q (new_AGEMA_signal_8549) ) ;
    buf_clk new_AGEMA_reg_buffer_6032 ( .C (clk), .D (new_AGEMA_signal_8552), .Q (new_AGEMA_signal_8553) ) ;
    buf_clk new_AGEMA_reg_buffer_6036 ( .C (clk), .D (new_AGEMA_signal_8556), .Q (new_AGEMA_signal_8557) ) ;
    buf_clk new_AGEMA_reg_buffer_6040 ( .C (clk), .D (new_AGEMA_signal_8560), .Q (new_AGEMA_signal_8561) ) ;
    buf_clk new_AGEMA_reg_buffer_6044 ( .C (clk), .D (new_AGEMA_signal_8564), .Q (new_AGEMA_signal_8565) ) ;
    buf_clk new_AGEMA_reg_buffer_6048 ( .C (clk), .D (new_AGEMA_signal_8568), .Q (new_AGEMA_signal_8569) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4156, RoundReg_Inst_ff_SDE_0_next_state}), .clk (clk), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4273, RoundReg_Inst_ff_SDE_1_next_state}), .clk (clk), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4158, RoundReg_Inst_ff_SDE_2_next_state}), .clk (clk), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4275, RoundReg_Inst_ff_SDE_3_next_state}), .clk (clk), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4277, RoundReg_Inst_ff_SDE_4_next_state}), .clk (clk), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4160, RoundReg_Inst_ff_SDE_5_next_state}), .clk (clk), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4162, RoundReg_Inst_ff_SDE_6_next_state}), .clk (clk), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4164, RoundReg_Inst_ff_SDE_7_next_state}), .clk (clk), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4166, RoundReg_Inst_ff_SDE_8_next_state}), .clk (clk), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4279, RoundReg_Inst_ff_SDE_9_next_state}), .clk (clk), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4168, RoundReg_Inst_ff_SDE_10_next_state}), .clk (clk), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4281, RoundReg_Inst_ff_SDE_11_next_state}), .clk (clk), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4283, RoundReg_Inst_ff_SDE_12_next_state}), .clk (clk), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4170, RoundReg_Inst_ff_SDE_13_next_state}), .clk (clk), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4172, RoundReg_Inst_ff_SDE_14_next_state}), .clk (clk), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4174, RoundReg_Inst_ff_SDE_15_next_state}), .clk (clk), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4176, RoundReg_Inst_ff_SDE_16_next_state}), .clk (clk), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4285, RoundReg_Inst_ff_SDE_17_next_state}), .clk (clk), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4178, RoundReg_Inst_ff_SDE_18_next_state}), .clk (clk), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4287, RoundReg_Inst_ff_SDE_19_next_state}), .clk (clk), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4289, RoundReg_Inst_ff_SDE_20_next_state}), .clk (clk), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4180, RoundReg_Inst_ff_SDE_21_next_state}), .clk (clk), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4182, RoundReg_Inst_ff_SDE_22_next_state}), .clk (clk), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4184, RoundReg_Inst_ff_SDE_23_next_state}), .clk (clk), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4186, RoundReg_Inst_ff_SDE_24_next_state}), .clk (clk), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4291, RoundReg_Inst_ff_SDE_25_next_state}), .clk (clk), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4188, RoundReg_Inst_ff_SDE_26_next_state}), .clk (clk), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4293, RoundReg_Inst_ff_SDE_27_next_state}), .clk (clk), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4295, RoundReg_Inst_ff_SDE_28_next_state}), .clk (clk), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4190, RoundReg_Inst_ff_SDE_29_next_state}), .clk (clk), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4192, RoundReg_Inst_ff_SDE_30_next_state}), .clk (clk), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4194, RoundReg_Inst_ff_SDE_31_next_state}), .clk (clk), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7781, new_AGEMA_signal_7777}), .clk (clk), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7789, new_AGEMA_signal_7785}), .clk (clk), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7797, new_AGEMA_signal_7793}), .clk (clk), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7805, new_AGEMA_signal_7801}), .clk (clk), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7813, new_AGEMA_signal_7809}), .clk (clk), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7821, new_AGEMA_signal_7817}), .clk (clk), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7829, new_AGEMA_signal_7825}), .clk (clk), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7837, new_AGEMA_signal_7833}), .clk (clk), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7845, new_AGEMA_signal_7841}), .clk (clk), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7853, new_AGEMA_signal_7849}), .clk (clk), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7861, new_AGEMA_signal_7857}), .clk (clk), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7869, new_AGEMA_signal_7865}), .clk (clk), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7877, new_AGEMA_signal_7873}), .clk (clk), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7885, new_AGEMA_signal_7881}), .clk (clk), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7893, new_AGEMA_signal_7889}), .clk (clk), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7901, new_AGEMA_signal_7897}), .clk (clk), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7909, new_AGEMA_signal_7905}), .clk (clk), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7917, new_AGEMA_signal_7913}), .clk (clk), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7925, new_AGEMA_signal_7921}), .clk (clk), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7933, new_AGEMA_signal_7929}), .clk (clk), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7941, new_AGEMA_signal_7937}), .clk (clk), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7949, new_AGEMA_signal_7945}), .clk (clk), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7957, new_AGEMA_signal_7953}), .clk (clk), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7965, new_AGEMA_signal_7961}), .clk (clk), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7973, new_AGEMA_signal_7969}), .clk (clk), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7981, new_AGEMA_signal_7977}), .clk (clk), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7989, new_AGEMA_signal_7985}), .clk (clk), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_7997, new_AGEMA_signal_7993}), .clk (clk), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8005, new_AGEMA_signal_8001}), .clk (clk), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8013, new_AGEMA_signal_8009}), .clk (clk), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8021, new_AGEMA_signal_8017}), .clk (clk), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8029, new_AGEMA_signal_8025}), .clk (clk), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8037, new_AGEMA_signal_8033}), .clk (clk), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8045, new_AGEMA_signal_8041}), .clk (clk), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8053, new_AGEMA_signal_8049}), .clk (clk), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8061, new_AGEMA_signal_8057}), .clk (clk), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8069, new_AGEMA_signal_8065}), .clk (clk), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8077, new_AGEMA_signal_8073}), .clk (clk), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8085, new_AGEMA_signal_8081}), .clk (clk), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8093, new_AGEMA_signal_8089}), .clk (clk), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8101, new_AGEMA_signal_8097}), .clk (clk), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8109, new_AGEMA_signal_8105}), .clk (clk), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8117, new_AGEMA_signal_8113}), .clk (clk), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8125, new_AGEMA_signal_8121}), .clk (clk), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8133, new_AGEMA_signal_8129}), .clk (clk), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8141, new_AGEMA_signal_8137}), .clk (clk), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8149, new_AGEMA_signal_8145}), .clk (clk), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8157, new_AGEMA_signal_8153}), .clk (clk), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8165, new_AGEMA_signal_8161}), .clk (clk), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8173, new_AGEMA_signal_8169}), .clk (clk), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8181, new_AGEMA_signal_8177}), .clk (clk), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8189, new_AGEMA_signal_8185}), .clk (clk), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8197, new_AGEMA_signal_8193}), .clk (clk), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8205, new_AGEMA_signal_8201}), .clk (clk), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8213, new_AGEMA_signal_8209}), .clk (clk), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8221, new_AGEMA_signal_8217}), .clk (clk), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8229, new_AGEMA_signal_8225}), .clk (clk), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8237, new_AGEMA_signal_8233}), .clk (clk), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8245, new_AGEMA_signal_8241}), .clk (clk), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8253, new_AGEMA_signal_8249}), .clk (clk), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8261, new_AGEMA_signal_8257}), .clk (clk), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8269, new_AGEMA_signal_8265}), .clk (clk), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8277, new_AGEMA_signal_8273}), .clk (clk), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8285, new_AGEMA_signal_8281}), .clk (clk), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8293, new_AGEMA_signal_8289}), .clk (clk), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8301, new_AGEMA_signal_8297}), .clk (clk), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8309, new_AGEMA_signal_8305}), .clk (clk), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8317, new_AGEMA_signal_8313}), .clk (clk), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8325, new_AGEMA_signal_8321}), .clk (clk), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8333, new_AGEMA_signal_8329}), .clk (clk), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8341, new_AGEMA_signal_8337}), .clk (clk), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8349, new_AGEMA_signal_8345}), .clk (clk), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8357, new_AGEMA_signal_8353}), .clk (clk), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8365, new_AGEMA_signal_8361}), .clk (clk), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8373, new_AGEMA_signal_8369}), .clk (clk), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8381, new_AGEMA_signal_8377}), .clk (clk), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8389, new_AGEMA_signal_8385}), .clk (clk), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8397, new_AGEMA_signal_8393}), .clk (clk), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8405, new_AGEMA_signal_8401}), .clk (clk), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8413, new_AGEMA_signal_8409}), .clk (clk), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8421, new_AGEMA_signal_8417}), .clk (clk), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8429, new_AGEMA_signal_8425}), .clk (clk), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8437, new_AGEMA_signal_8433}), .clk (clk), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8445, new_AGEMA_signal_8441}), .clk (clk), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8453, new_AGEMA_signal_8449}), .clk (clk), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8461, new_AGEMA_signal_8457}), .clk (clk), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8469, new_AGEMA_signal_8465}), .clk (clk), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8477, new_AGEMA_signal_8473}), .clk (clk), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8485, new_AGEMA_signal_8481}), .clk (clk), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8493, new_AGEMA_signal_8489}), .clk (clk), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8501, new_AGEMA_signal_8497}), .clk (clk), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8509, new_AGEMA_signal_8505}), .clk (clk), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8517, new_AGEMA_signal_8513}), .clk (clk), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8525, new_AGEMA_signal_8521}), .clk (clk), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8533, new_AGEMA_signal_8529}), .clk (clk), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_8541, new_AGEMA_signal_8537}), .clk (clk), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4056, KeyReg_Inst_ff_SDE_0_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2339, KSSubBytesInput[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4208, KeyReg_Inst_ff_SDE_1_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2456, KSSubBytesInput[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4210, KeyReg_Inst_ff_SDE_2_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2489, KSSubBytesInput[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4212, KeyReg_Inst_ff_SDE_3_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2522, KSSubBytesInput[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4214, KeyReg_Inst_ff_SDE_4_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2555, KSSubBytesInput[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4216, KeyReg_Inst_ff_SDE_5_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2588, KSSubBytesInput[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4218, KeyReg_Inst_ff_SDE_6_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2621, KSSubBytesInput[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4220, KeyReg_Inst_ff_SDE_7_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2654, KSSubBytesInput[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4058, KeyReg_Inst_ff_SDE_8_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2687, KSSubBytesInput[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4222, KeyReg_Inst_ff_SDE_9_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2720, KSSubBytesInput[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4224, KeyReg_Inst_ff_SDE_10_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2372, KSSubBytesInput[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4226, KeyReg_Inst_ff_SDE_11_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2405, KSSubBytesInput[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4228, KeyReg_Inst_ff_SDE_12_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2432, KSSubBytesInput[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4230, KeyReg_Inst_ff_SDE_13_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2435, KSSubBytesInput[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4232, KeyReg_Inst_ff_SDE_14_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2438, KSSubBytesInput[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4234, KeyReg_Inst_ff_SDE_15_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2441, KSSubBytesInput[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4060, KeyReg_Inst_ff_SDE_16_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2444, KSSubBytesInput[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4236, KeyReg_Inst_ff_SDE_17_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2447, KSSubBytesInput[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4238, KeyReg_Inst_ff_SDE_18_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2450, KSSubBytesInput[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4240, KeyReg_Inst_ff_SDE_19_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2453, KSSubBytesInput[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4242, KeyReg_Inst_ff_SDE_20_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2459, KSSubBytesInput[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4244, KeyReg_Inst_ff_SDE_21_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2462, KSSubBytesInput[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4246, KeyReg_Inst_ff_SDE_22_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2465, KSSubBytesInput[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4248, KeyReg_Inst_ff_SDE_23_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2468, KSSubBytesInput[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4250, KeyReg_Inst_ff_SDE_24_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2471, KSSubBytesInput[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4297, KeyReg_Inst_ff_SDE_25_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2474, KSSubBytesInput[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4299, KeyReg_Inst_ff_SDE_26_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2477, KSSubBytesInput[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4301, KeyReg_Inst_ff_SDE_27_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2480, KSSubBytesInput[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4303, KeyReg_Inst_ff_SDE_28_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2483, KSSubBytesInput[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4305, KeyReg_Inst_ff_SDE_29_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2486, KSSubBytesInput[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4307, KeyReg_Inst_ff_SDE_30_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2492, KSSubBytesInput[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4309, KeyReg_Inst_ff_SDE_31_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2495, KSSubBytesInput[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3899, KeyReg_Inst_ff_SDE_32_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2498, RoundKey[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4062, KeyReg_Inst_ff_SDE_33_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2501, RoundKey[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4064, KeyReg_Inst_ff_SDE_34_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2504, RoundKey[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4066, KeyReg_Inst_ff_SDE_35_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2507, RoundKey[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4068, KeyReg_Inst_ff_SDE_36_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2510, RoundKey[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4070, KeyReg_Inst_ff_SDE_37_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2513, RoundKey[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4072, KeyReg_Inst_ff_SDE_38_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2516, RoundKey[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4074, KeyReg_Inst_ff_SDE_39_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2519, RoundKey[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3901, KeyReg_Inst_ff_SDE_40_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2525, RoundKey[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4076, KeyReg_Inst_ff_SDE_41_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2528, RoundKey[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4078, KeyReg_Inst_ff_SDE_42_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2531, RoundKey[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4080, KeyReg_Inst_ff_SDE_43_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2534, RoundKey[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4082, KeyReg_Inst_ff_SDE_44_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2537, RoundKey[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4084, KeyReg_Inst_ff_SDE_45_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2540, RoundKey[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4086, KeyReg_Inst_ff_SDE_46_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2543, RoundKey[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4088, KeyReg_Inst_ff_SDE_47_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2546, RoundKey[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3903, KeyReg_Inst_ff_SDE_48_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2549, RoundKey[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4090, KeyReg_Inst_ff_SDE_49_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2552, RoundKey[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4092, KeyReg_Inst_ff_SDE_50_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2558, RoundKey[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4094, KeyReg_Inst_ff_SDE_51_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2561, RoundKey[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4096, KeyReg_Inst_ff_SDE_52_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2564, RoundKey[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4098, KeyReg_Inst_ff_SDE_53_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2567, RoundKey[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4100, KeyReg_Inst_ff_SDE_54_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2570, RoundKey[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4102, KeyReg_Inst_ff_SDE_55_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2573, RoundKey[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4104, KeyReg_Inst_ff_SDE_56_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2576, RoundKey[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4252, KeyReg_Inst_ff_SDE_57_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2579, RoundKey[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4254, KeyReg_Inst_ff_SDE_58_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2582, RoundKey[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4256, KeyReg_Inst_ff_SDE_59_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2585, RoundKey[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4258, KeyReg_Inst_ff_SDE_60_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2591, RoundKey[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4260, KeyReg_Inst_ff_SDE_61_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2594, RoundKey[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4262, KeyReg_Inst_ff_SDE_62_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2597, RoundKey[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4264, KeyReg_Inst_ff_SDE_63_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2600, RoundKey[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3753, KeyReg_Inst_ff_SDE_64_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2603, RoundKey[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3905, KeyReg_Inst_ff_SDE_65_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2606, RoundKey[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3907, KeyReg_Inst_ff_SDE_66_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2609, RoundKey[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3909, KeyReg_Inst_ff_SDE_67_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2612, RoundKey[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3911, KeyReg_Inst_ff_SDE_68_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2615, RoundKey[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3913, KeyReg_Inst_ff_SDE_69_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2618, RoundKey[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3915, KeyReg_Inst_ff_SDE_70_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2624, RoundKey[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3917, KeyReg_Inst_ff_SDE_71_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2627, RoundKey[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3755, KeyReg_Inst_ff_SDE_72_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2630, RoundKey[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3919, KeyReg_Inst_ff_SDE_73_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2633, RoundKey[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3921, KeyReg_Inst_ff_SDE_74_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2636, RoundKey[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3923, KeyReg_Inst_ff_SDE_75_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2639, RoundKey[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3925, KeyReg_Inst_ff_SDE_76_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2642, RoundKey[76]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3927, KeyReg_Inst_ff_SDE_77_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2645, RoundKey[77]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3929, KeyReg_Inst_ff_SDE_78_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2648, RoundKey[78]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3931, KeyReg_Inst_ff_SDE_79_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2651, RoundKey[79]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3757, KeyReg_Inst_ff_SDE_80_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2657, RoundKey[80]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3933, KeyReg_Inst_ff_SDE_81_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2660, RoundKey[81]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3935, KeyReg_Inst_ff_SDE_82_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2663, RoundKey[82]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3937, KeyReg_Inst_ff_SDE_83_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2666, RoundKey[83]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3939, KeyReg_Inst_ff_SDE_84_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2669, RoundKey[84]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3941, KeyReg_Inst_ff_SDE_85_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2672, RoundKey[85]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3943, KeyReg_Inst_ff_SDE_86_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2675, RoundKey[86]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3945, KeyReg_Inst_ff_SDE_87_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2678, RoundKey[87]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3947, KeyReg_Inst_ff_SDE_88_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2681, RoundKey[88]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4106, KeyReg_Inst_ff_SDE_89_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2684, RoundKey[89]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4108, KeyReg_Inst_ff_SDE_90_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2690, RoundKey[90]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4110, KeyReg_Inst_ff_SDE_91_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2693, RoundKey[91]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4112, KeyReg_Inst_ff_SDE_92_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2696, RoundKey[92]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4114, KeyReg_Inst_ff_SDE_93_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2699, RoundKey[93]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4116, KeyReg_Inst_ff_SDE_94_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2702, RoundKey[94]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_4118, KeyReg_Inst_ff_SDE_95_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2705, RoundKey[95]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3658, KeyReg_Inst_ff_SDE_96_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2708, RoundKey[96]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3759, KeyReg_Inst_ff_SDE_97_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2711, RoundKey[97]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3761, KeyReg_Inst_ff_SDE_98_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2714, RoundKey[98]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3763, KeyReg_Inst_ff_SDE_99_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2717, RoundKey[99]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3765, KeyReg_Inst_ff_SDE_100_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2342, RoundKey[100]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3767, KeyReg_Inst_ff_SDE_101_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2345, RoundKey[101]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3769, KeyReg_Inst_ff_SDE_102_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2348, RoundKey[102]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3771, KeyReg_Inst_ff_SDE_103_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2351, RoundKey[103]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3660, KeyReg_Inst_ff_SDE_104_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2354, RoundKey[104]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3773, KeyReg_Inst_ff_SDE_105_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2357, RoundKey[105]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3775, KeyReg_Inst_ff_SDE_106_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2360, RoundKey[106]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3777, KeyReg_Inst_ff_SDE_107_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2363, RoundKey[107]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3779, KeyReg_Inst_ff_SDE_108_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2366, RoundKey[108]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3781, KeyReg_Inst_ff_SDE_109_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2369, RoundKey[109]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3783, KeyReg_Inst_ff_SDE_110_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2375, RoundKey[110]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3785, KeyReg_Inst_ff_SDE_111_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2378, RoundKey[111]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3662, KeyReg_Inst_ff_SDE_112_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2381, RoundKey[112]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3787, KeyReg_Inst_ff_SDE_113_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2384, RoundKey[113]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3789, KeyReg_Inst_ff_SDE_114_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2387, RoundKey[114]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3791, KeyReg_Inst_ff_SDE_115_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2390, RoundKey[115]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3793, KeyReg_Inst_ff_SDE_116_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2393, RoundKey[116]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3795, KeyReg_Inst_ff_SDE_117_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2396, RoundKey[117]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3797, KeyReg_Inst_ff_SDE_118_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2399, RoundKey[118]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3799, KeyReg_Inst_ff_SDE_119_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2402, RoundKey[119]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3801, KeyReg_Inst_ff_SDE_120_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2408, RoundKey[120]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3949, KeyReg_Inst_ff_SDE_121_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2411, RoundKey[121]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3951, KeyReg_Inst_ff_SDE_122_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2414, RoundKey[122]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3953, KeyReg_Inst_ff_SDE_123_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2417, RoundKey[123]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3955, KeyReg_Inst_ff_SDE_124_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2420, RoundKey[124]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3957, KeyReg_Inst_ff_SDE_125_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2423, RoundKey[125]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3959, KeyReg_Inst_ff_SDE_126_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2426, RoundKey[126]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .D ({new_AGEMA_signal_3961, KeyReg_Inst_ff_SDE_127_next_state}), .clk (clk), .Q ({new_AGEMA_signal_2429, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .D (new_AGEMA_signal_8545), .CK (clk), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .D (new_AGEMA_signal_8549), .CK (clk), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .D (new_AGEMA_signal_8553), .CK (clk), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .D (new_AGEMA_signal_8557), .CK (clk), .Q (RoundCounter[3]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_0__FF_FF ( .D (new_AGEMA_signal_8561), .CK (clk), .Q (InRoundCounter[0]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_1__FF_FF ( .D (new_AGEMA_signal_8565), .CK (clk), .Q (InRoundCounter[1]), .QN () ) ;
    DFF_X1 InRoundCounterIns_count_reg_2__FF_FF ( .D (new_AGEMA_signal_8569), .CK (clk), .Q (InRoundCounter[2]), .QN () ) ;
endmodule
