/* modified netlist. Source: module AES in file /AES_round-based/AGEMA/AES.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module AES_HPC2_ClockGating_d3 (plaintext_s0, key_s0, clk, reset, key_s1, key_s2, key_s3, plaintext_s1, plaintext_s2, plaintext_s3, Fresh, ciphertext_s0, done, ciphertext_s1, ciphertext_s2, ciphertext_s3, Synch);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] key_s1 ;
    input [127:0] key_s2 ;
    input [127:0] key_s3 ;
    input [127:0] plaintext_s1 ;
    input [127:0] plaintext_s2 ;
    input [127:0] plaintext_s3 ;
    input [4079:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    output [127:0] ciphertext_s2 ;
    output [127:0] ciphertext_s3 ;
    output Synch ;
    wire n283 ;
    wire n285 ;
    wire n314 ;
    wire n315 ;
    wire n316 ;
    wire n317 ;
    wire n318 ;
    wire n319 ;
    wire n320 ;
    wire n321 ;
    wire n322 ;
    wire n323 ;
    wire n324 ;
    wire n325 ;
    wire n326 ;
    wire n327 ;
    wire n328 ;
    wire n329 ;
    wire n330 ;
    wire n331 ;
    wire n332 ;
    wire n333 ;
    wire n334 ;
    wire n335 ;
    wire n336 ;
    wire n337 ;
    wire n338 ;
    wire n339 ;
    wire RoundReg_Inst_ff_SDE_0_next_state ;
    wire RoundReg_Inst_ff_SDE_1_next_state ;
    wire RoundReg_Inst_ff_SDE_2_next_state ;
    wire RoundReg_Inst_ff_SDE_3_next_state ;
    wire RoundReg_Inst_ff_SDE_4_next_state ;
    wire RoundReg_Inst_ff_SDE_5_next_state ;
    wire RoundReg_Inst_ff_SDE_6_next_state ;
    wire RoundReg_Inst_ff_SDE_7_next_state ;
    wire RoundReg_Inst_ff_SDE_8_next_state ;
    wire RoundReg_Inst_ff_SDE_9_next_state ;
    wire RoundReg_Inst_ff_SDE_10_next_state ;
    wire RoundReg_Inst_ff_SDE_11_next_state ;
    wire RoundReg_Inst_ff_SDE_12_next_state ;
    wire RoundReg_Inst_ff_SDE_13_next_state ;
    wire RoundReg_Inst_ff_SDE_14_next_state ;
    wire RoundReg_Inst_ff_SDE_15_next_state ;
    wire RoundReg_Inst_ff_SDE_16_next_state ;
    wire RoundReg_Inst_ff_SDE_17_next_state ;
    wire RoundReg_Inst_ff_SDE_18_next_state ;
    wire RoundReg_Inst_ff_SDE_19_next_state ;
    wire RoundReg_Inst_ff_SDE_20_next_state ;
    wire RoundReg_Inst_ff_SDE_21_next_state ;
    wire RoundReg_Inst_ff_SDE_22_next_state ;
    wire RoundReg_Inst_ff_SDE_23_next_state ;
    wire RoundReg_Inst_ff_SDE_24_next_state ;
    wire RoundReg_Inst_ff_SDE_25_next_state ;
    wire RoundReg_Inst_ff_SDE_26_next_state ;
    wire RoundReg_Inst_ff_SDE_27_next_state ;
    wire RoundReg_Inst_ff_SDE_28_next_state ;
    wire RoundReg_Inst_ff_SDE_29_next_state ;
    wire RoundReg_Inst_ff_SDE_30_next_state ;
    wire RoundReg_Inst_ff_SDE_31_next_state ;
    wire RoundReg_Inst_ff_SDE_32_next_state ;
    wire RoundReg_Inst_ff_SDE_33_next_state ;
    wire RoundReg_Inst_ff_SDE_34_next_state ;
    wire RoundReg_Inst_ff_SDE_35_next_state ;
    wire RoundReg_Inst_ff_SDE_36_next_state ;
    wire RoundReg_Inst_ff_SDE_37_next_state ;
    wire RoundReg_Inst_ff_SDE_38_next_state ;
    wire RoundReg_Inst_ff_SDE_39_next_state ;
    wire RoundReg_Inst_ff_SDE_40_next_state ;
    wire RoundReg_Inst_ff_SDE_41_next_state ;
    wire RoundReg_Inst_ff_SDE_42_next_state ;
    wire RoundReg_Inst_ff_SDE_43_next_state ;
    wire RoundReg_Inst_ff_SDE_44_next_state ;
    wire RoundReg_Inst_ff_SDE_45_next_state ;
    wire RoundReg_Inst_ff_SDE_46_next_state ;
    wire RoundReg_Inst_ff_SDE_47_next_state ;
    wire RoundReg_Inst_ff_SDE_48_next_state ;
    wire RoundReg_Inst_ff_SDE_49_next_state ;
    wire RoundReg_Inst_ff_SDE_50_next_state ;
    wire RoundReg_Inst_ff_SDE_51_next_state ;
    wire RoundReg_Inst_ff_SDE_52_next_state ;
    wire RoundReg_Inst_ff_SDE_53_next_state ;
    wire RoundReg_Inst_ff_SDE_54_next_state ;
    wire RoundReg_Inst_ff_SDE_55_next_state ;
    wire RoundReg_Inst_ff_SDE_56_next_state ;
    wire RoundReg_Inst_ff_SDE_57_next_state ;
    wire RoundReg_Inst_ff_SDE_58_next_state ;
    wire RoundReg_Inst_ff_SDE_59_next_state ;
    wire RoundReg_Inst_ff_SDE_60_next_state ;
    wire RoundReg_Inst_ff_SDE_61_next_state ;
    wire RoundReg_Inst_ff_SDE_62_next_state ;
    wire RoundReg_Inst_ff_SDE_63_next_state ;
    wire RoundReg_Inst_ff_SDE_64_next_state ;
    wire RoundReg_Inst_ff_SDE_65_next_state ;
    wire RoundReg_Inst_ff_SDE_66_next_state ;
    wire RoundReg_Inst_ff_SDE_67_next_state ;
    wire RoundReg_Inst_ff_SDE_68_next_state ;
    wire RoundReg_Inst_ff_SDE_69_next_state ;
    wire RoundReg_Inst_ff_SDE_70_next_state ;
    wire RoundReg_Inst_ff_SDE_71_next_state ;
    wire RoundReg_Inst_ff_SDE_72_next_state ;
    wire RoundReg_Inst_ff_SDE_73_next_state ;
    wire RoundReg_Inst_ff_SDE_74_next_state ;
    wire RoundReg_Inst_ff_SDE_75_next_state ;
    wire RoundReg_Inst_ff_SDE_76_next_state ;
    wire RoundReg_Inst_ff_SDE_77_next_state ;
    wire RoundReg_Inst_ff_SDE_78_next_state ;
    wire RoundReg_Inst_ff_SDE_79_next_state ;
    wire RoundReg_Inst_ff_SDE_80_next_state ;
    wire RoundReg_Inst_ff_SDE_81_next_state ;
    wire RoundReg_Inst_ff_SDE_82_next_state ;
    wire RoundReg_Inst_ff_SDE_83_next_state ;
    wire RoundReg_Inst_ff_SDE_84_next_state ;
    wire RoundReg_Inst_ff_SDE_85_next_state ;
    wire RoundReg_Inst_ff_SDE_86_next_state ;
    wire RoundReg_Inst_ff_SDE_87_next_state ;
    wire RoundReg_Inst_ff_SDE_88_next_state ;
    wire RoundReg_Inst_ff_SDE_89_next_state ;
    wire RoundReg_Inst_ff_SDE_90_next_state ;
    wire RoundReg_Inst_ff_SDE_91_next_state ;
    wire RoundReg_Inst_ff_SDE_92_next_state ;
    wire RoundReg_Inst_ff_SDE_93_next_state ;
    wire RoundReg_Inst_ff_SDE_94_next_state ;
    wire RoundReg_Inst_ff_SDE_95_next_state ;
    wire RoundReg_Inst_ff_SDE_96_next_state ;
    wire RoundReg_Inst_ff_SDE_97_next_state ;
    wire RoundReg_Inst_ff_SDE_98_next_state ;
    wire RoundReg_Inst_ff_SDE_99_next_state ;
    wire RoundReg_Inst_ff_SDE_100_next_state ;
    wire RoundReg_Inst_ff_SDE_101_next_state ;
    wire RoundReg_Inst_ff_SDE_102_next_state ;
    wire RoundReg_Inst_ff_SDE_103_next_state ;
    wire RoundReg_Inst_ff_SDE_104_next_state ;
    wire RoundReg_Inst_ff_SDE_105_next_state ;
    wire RoundReg_Inst_ff_SDE_106_next_state ;
    wire RoundReg_Inst_ff_SDE_107_next_state ;
    wire RoundReg_Inst_ff_SDE_108_next_state ;
    wire RoundReg_Inst_ff_SDE_109_next_state ;
    wire RoundReg_Inst_ff_SDE_110_next_state ;
    wire RoundReg_Inst_ff_SDE_111_next_state ;
    wire RoundReg_Inst_ff_SDE_112_next_state ;
    wire RoundReg_Inst_ff_SDE_113_next_state ;
    wire RoundReg_Inst_ff_SDE_114_next_state ;
    wire RoundReg_Inst_ff_SDE_115_next_state ;
    wire RoundReg_Inst_ff_SDE_116_next_state ;
    wire RoundReg_Inst_ff_SDE_117_next_state ;
    wire RoundReg_Inst_ff_SDE_118_next_state ;
    wire RoundReg_Inst_ff_SDE_119_next_state ;
    wire RoundReg_Inst_ff_SDE_120_next_state ;
    wire RoundReg_Inst_ff_SDE_121_next_state ;
    wire RoundReg_Inst_ff_SDE_122_next_state ;
    wire RoundReg_Inst_ff_SDE_123_next_state ;
    wire RoundReg_Inst_ff_SDE_124_next_state ;
    wire RoundReg_Inst_ff_SDE_125_next_state ;
    wire RoundReg_Inst_ff_SDE_126_next_state ;
    wire RoundReg_Inst_ff_SDE_127_next_state ;
    wire SubBytesIns_Inst_Sbox_0_L29 ;
    wire SubBytesIns_Inst_Sbox_0_L28 ;
    wire SubBytesIns_Inst_Sbox_0_L27 ;
    wire SubBytesIns_Inst_Sbox_0_L26 ;
    wire SubBytesIns_Inst_Sbox_0_L25 ;
    wire SubBytesIns_Inst_Sbox_0_L24 ;
    wire SubBytesIns_Inst_Sbox_0_L23 ;
    wire SubBytesIns_Inst_Sbox_0_L22 ;
    wire SubBytesIns_Inst_Sbox_0_L21 ;
    wire SubBytesIns_Inst_Sbox_0_L20 ;
    wire SubBytesIns_Inst_Sbox_0_L19 ;
    wire SubBytesIns_Inst_Sbox_0_L18 ;
    wire SubBytesIns_Inst_Sbox_0_L17 ;
    wire SubBytesIns_Inst_Sbox_0_L16 ;
    wire SubBytesIns_Inst_Sbox_0_L15 ;
    wire SubBytesIns_Inst_Sbox_0_L14 ;
    wire SubBytesIns_Inst_Sbox_0_L13 ;
    wire SubBytesIns_Inst_Sbox_0_L12 ;
    wire SubBytesIns_Inst_Sbox_0_L11 ;
    wire SubBytesIns_Inst_Sbox_0_L10 ;
    wire SubBytesIns_Inst_Sbox_0_L9 ;
    wire SubBytesIns_Inst_Sbox_0_L8 ;
    wire SubBytesIns_Inst_Sbox_0_L7 ;
    wire SubBytesIns_Inst_Sbox_0_L6 ;
    wire SubBytesIns_Inst_Sbox_0_L5 ;
    wire SubBytesIns_Inst_Sbox_0_L4 ;
    wire SubBytesIns_Inst_Sbox_0_L3 ;
    wire SubBytesIns_Inst_Sbox_0_L2 ;
    wire SubBytesIns_Inst_Sbox_0_L1 ;
    wire SubBytesIns_Inst_Sbox_0_L0 ;
    wire SubBytesIns_Inst_Sbox_0_M63 ;
    wire SubBytesIns_Inst_Sbox_0_M62 ;
    wire SubBytesIns_Inst_Sbox_0_M61 ;
    wire SubBytesIns_Inst_Sbox_0_M60 ;
    wire SubBytesIns_Inst_Sbox_0_M59 ;
    wire SubBytesIns_Inst_Sbox_0_M58 ;
    wire SubBytesIns_Inst_Sbox_0_M57 ;
    wire SubBytesIns_Inst_Sbox_0_M56 ;
    wire SubBytesIns_Inst_Sbox_0_M55 ;
    wire SubBytesIns_Inst_Sbox_0_M54 ;
    wire SubBytesIns_Inst_Sbox_0_M53 ;
    wire SubBytesIns_Inst_Sbox_0_M52 ;
    wire SubBytesIns_Inst_Sbox_0_M51 ;
    wire SubBytesIns_Inst_Sbox_0_M50 ;
    wire SubBytesIns_Inst_Sbox_0_M49 ;
    wire SubBytesIns_Inst_Sbox_0_M48 ;
    wire SubBytesIns_Inst_Sbox_0_M47 ;
    wire SubBytesIns_Inst_Sbox_0_M46 ;
    wire SubBytesIns_Inst_Sbox_0_M45 ;
    wire SubBytesIns_Inst_Sbox_0_M44 ;
    wire SubBytesIns_Inst_Sbox_0_M43 ;
    wire SubBytesIns_Inst_Sbox_0_M42 ;
    wire SubBytesIns_Inst_Sbox_0_M41 ;
    wire SubBytesIns_Inst_Sbox_0_M40 ;
    wire SubBytesIns_Inst_Sbox_0_M39 ;
    wire SubBytesIns_Inst_Sbox_0_M38 ;
    wire SubBytesIns_Inst_Sbox_0_M37 ;
    wire SubBytesIns_Inst_Sbox_0_M36 ;
    wire SubBytesIns_Inst_Sbox_0_M35 ;
    wire SubBytesIns_Inst_Sbox_0_M34 ;
    wire SubBytesIns_Inst_Sbox_0_M33 ;
    wire SubBytesIns_Inst_Sbox_0_M32 ;
    wire SubBytesIns_Inst_Sbox_0_M31 ;
    wire SubBytesIns_Inst_Sbox_0_M30 ;
    wire SubBytesIns_Inst_Sbox_0_M29 ;
    wire SubBytesIns_Inst_Sbox_0_M28 ;
    wire SubBytesIns_Inst_Sbox_0_M27 ;
    wire SubBytesIns_Inst_Sbox_0_M26 ;
    wire SubBytesIns_Inst_Sbox_0_M25 ;
    wire SubBytesIns_Inst_Sbox_0_M24 ;
    wire SubBytesIns_Inst_Sbox_0_M23 ;
    wire SubBytesIns_Inst_Sbox_0_M22 ;
    wire SubBytesIns_Inst_Sbox_0_M21 ;
    wire SubBytesIns_Inst_Sbox_0_M20 ;
    wire SubBytesIns_Inst_Sbox_0_M19 ;
    wire SubBytesIns_Inst_Sbox_0_M18 ;
    wire SubBytesIns_Inst_Sbox_0_M17 ;
    wire SubBytesIns_Inst_Sbox_0_M16 ;
    wire SubBytesIns_Inst_Sbox_0_M15 ;
    wire SubBytesIns_Inst_Sbox_0_M14 ;
    wire SubBytesIns_Inst_Sbox_0_M13 ;
    wire SubBytesIns_Inst_Sbox_0_M12 ;
    wire SubBytesIns_Inst_Sbox_0_M11 ;
    wire SubBytesIns_Inst_Sbox_0_M10 ;
    wire SubBytesIns_Inst_Sbox_0_M9 ;
    wire SubBytesIns_Inst_Sbox_0_M8 ;
    wire SubBytesIns_Inst_Sbox_0_M7 ;
    wire SubBytesIns_Inst_Sbox_0_M6 ;
    wire SubBytesIns_Inst_Sbox_0_M5 ;
    wire SubBytesIns_Inst_Sbox_0_M4 ;
    wire SubBytesIns_Inst_Sbox_0_M3 ;
    wire SubBytesIns_Inst_Sbox_0_M2 ;
    wire SubBytesIns_Inst_Sbox_0_M1 ;
    wire SubBytesIns_Inst_Sbox_0_T27 ;
    wire SubBytesIns_Inst_Sbox_0_T26 ;
    wire SubBytesIns_Inst_Sbox_0_T25 ;
    wire SubBytesIns_Inst_Sbox_0_T24 ;
    wire SubBytesIns_Inst_Sbox_0_T23 ;
    wire SubBytesIns_Inst_Sbox_0_T22 ;
    wire SubBytesIns_Inst_Sbox_0_T21 ;
    wire SubBytesIns_Inst_Sbox_0_T20 ;
    wire SubBytesIns_Inst_Sbox_0_T19 ;
    wire SubBytesIns_Inst_Sbox_0_T18 ;
    wire SubBytesIns_Inst_Sbox_0_T17 ;
    wire SubBytesIns_Inst_Sbox_0_T16 ;
    wire SubBytesIns_Inst_Sbox_0_T15 ;
    wire SubBytesIns_Inst_Sbox_0_T14 ;
    wire SubBytesIns_Inst_Sbox_0_T13 ;
    wire SubBytesIns_Inst_Sbox_0_T12 ;
    wire SubBytesIns_Inst_Sbox_0_T11 ;
    wire SubBytesIns_Inst_Sbox_0_T10 ;
    wire SubBytesIns_Inst_Sbox_0_T9 ;
    wire SubBytesIns_Inst_Sbox_0_T8 ;
    wire SubBytesIns_Inst_Sbox_0_T7 ;
    wire SubBytesIns_Inst_Sbox_0_T6 ;
    wire SubBytesIns_Inst_Sbox_0_T5 ;
    wire SubBytesIns_Inst_Sbox_0_T4 ;
    wire SubBytesIns_Inst_Sbox_0_T3 ;
    wire SubBytesIns_Inst_Sbox_0_T2 ;
    wire SubBytesIns_Inst_Sbox_0_T1 ;
    wire SubBytesIns_Inst_Sbox_1_L29 ;
    wire SubBytesIns_Inst_Sbox_1_L28 ;
    wire SubBytesIns_Inst_Sbox_1_L27 ;
    wire SubBytesIns_Inst_Sbox_1_L26 ;
    wire SubBytesIns_Inst_Sbox_1_L25 ;
    wire SubBytesIns_Inst_Sbox_1_L24 ;
    wire SubBytesIns_Inst_Sbox_1_L23 ;
    wire SubBytesIns_Inst_Sbox_1_L22 ;
    wire SubBytesIns_Inst_Sbox_1_L21 ;
    wire SubBytesIns_Inst_Sbox_1_L20 ;
    wire SubBytesIns_Inst_Sbox_1_L19 ;
    wire SubBytesIns_Inst_Sbox_1_L18 ;
    wire SubBytesIns_Inst_Sbox_1_L17 ;
    wire SubBytesIns_Inst_Sbox_1_L16 ;
    wire SubBytesIns_Inst_Sbox_1_L15 ;
    wire SubBytesIns_Inst_Sbox_1_L14 ;
    wire SubBytesIns_Inst_Sbox_1_L13 ;
    wire SubBytesIns_Inst_Sbox_1_L12 ;
    wire SubBytesIns_Inst_Sbox_1_L11 ;
    wire SubBytesIns_Inst_Sbox_1_L10 ;
    wire SubBytesIns_Inst_Sbox_1_L9 ;
    wire SubBytesIns_Inst_Sbox_1_L8 ;
    wire SubBytesIns_Inst_Sbox_1_L7 ;
    wire SubBytesIns_Inst_Sbox_1_L6 ;
    wire SubBytesIns_Inst_Sbox_1_L5 ;
    wire SubBytesIns_Inst_Sbox_1_L4 ;
    wire SubBytesIns_Inst_Sbox_1_L3 ;
    wire SubBytesIns_Inst_Sbox_1_L2 ;
    wire SubBytesIns_Inst_Sbox_1_L1 ;
    wire SubBytesIns_Inst_Sbox_1_L0 ;
    wire SubBytesIns_Inst_Sbox_1_M63 ;
    wire SubBytesIns_Inst_Sbox_1_M62 ;
    wire SubBytesIns_Inst_Sbox_1_M61 ;
    wire SubBytesIns_Inst_Sbox_1_M60 ;
    wire SubBytesIns_Inst_Sbox_1_M59 ;
    wire SubBytesIns_Inst_Sbox_1_M58 ;
    wire SubBytesIns_Inst_Sbox_1_M57 ;
    wire SubBytesIns_Inst_Sbox_1_M56 ;
    wire SubBytesIns_Inst_Sbox_1_M55 ;
    wire SubBytesIns_Inst_Sbox_1_M54 ;
    wire SubBytesIns_Inst_Sbox_1_M53 ;
    wire SubBytesIns_Inst_Sbox_1_M52 ;
    wire SubBytesIns_Inst_Sbox_1_M51 ;
    wire SubBytesIns_Inst_Sbox_1_M50 ;
    wire SubBytesIns_Inst_Sbox_1_M49 ;
    wire SubBytesIns_Inst_Sbox_1_M48 ;
    wire SubBytesIns_Inst_Sbox_1_M47 ;
    wire SubBytesIns_Inst_Sbox_1_M46 ;
    wire SubBytesIns_Inst_Sbox_1_M45 ;
    wire SubBytesIns_Inst_Sbox_1_M44 ;
    wire SubBytesIns_Inst_Sbox_1_M43 ;
    wire SubBytesIns_Inst_Sbox_1_M42 ;
    wire SubBytesIns_Inst_Sbox_1_M41 ;
    wire SubBytesIns_Inst_Sbox_1_M40 ;
    wire SubBytesIns_Inst_Sbox_1_M39 ;
    wire SubBytesIns_Inst_Sbox_1_M38 ;
    wire SubBytesIns_Inst_Sbox_1_M37 ;
    wire SubBytesIns_Inst_Sbox_1_M36 ;
    wire SubBytesIns_Inst_Sbox_1_M35 ;
    wire SubBytesIns_Inst_Sbox_1_M34 ;
    wire SubBytesIns_Inst_Sbox_1_M33 ;
    wire SubBytesIns_Inst_Sbox_1_M32 ;
    wire SubBytesIns_Inst_Sbox_1_M31 ;
    wire SubBytesIns_Inst_Sbox_1_M30 ;
    wire SubBytesIns_Inst_Sbox_1_M29 ;
    wire SubBytesIns_Inst_Sbox_1_M28 ;
    wire SubBytesIns_Inst_Sbox_1_M27 ;
    wire SubBytesIns_Inst_Sbox_1_M26 ;
    wire SubBytesIns_Inst_Sbox_1_M25 ;
    wire SubBytesIns_Inst_Sbox_1_M24 ;
    wire SubBytesIns_Inst_Sbox_1_M23 ;
    wire SubBytesIns_Inst_Sbox_1_M22 ;
    wire SubBytesIns_Inst_Sbox_1_M21 ;
    wire SubBytesIns_Inst_Sbox_1_M20 ;
    wire SubBytesIns_Inst_Sbox_1_M19 ;
    wire SubBytesIns_Inst_Sbox_1_M18 ;
    wire SubBytesIns_Inst_Sbox_1_M17 ;
    wire SubBytesIns_Inst_Sbox_1_M16 ;
    wire SubBytesIns_Inst_Sbox_1_M15 ;
    wire SubBytesIns_Inst_Sbox_1_M14 ;
    wire SubBytesIns_Inst_Sbox_1_M13 ;
    wire SubBytesIns_Inst_Sbox_1_M12 ;
    wire SubBytesIns_Inst_Sbox_1_M11 ;
    wire SubBytesIns_Inst_Sbox_1_M10 ;
    wire SubBytesIns_Inst_Sbox_1_M9 ;
    wire SubBytesIns_Inst_Sbox_1_M8 ;
    wire SubBytesIns_Inst_Sbox_1_M7 ;
    wire SubBytesIns_Inst_Sbox_1_M6 ;
    wire SubBytesIns_Inst_Sbox_1_M5 ;
    wire SubBytesIns_Inst_Sbox_1_M4 ;
    wire SubBytesIns_Inst_Sbox_1_M3 ;
    wire SubBytesIns_Inst_Sbox_1_M2 ;
    wire SubBytesIns_Inst_Sbox_1_M1 ;
    wire SubBytesIns_Inst_Sbox_1_T27 ;
    wire SubBytesIns_Inst_Sbox_1_T26 ;
    wire SubBytesIns_Inst_Sbox_1_T25 ;
    wire SubBytesIns_Inst_Sbox_1_T24 ;
    wire SubBytesIns_Inst_Sbox_1_T23 ;
    wire SubBytesIns_Inst_Sbox_1_T22 ;
    wire SubBytesIns_Inst_Sbox_1_T21 ;
    wire SubBytesIns_Inst_Sbox_1_T20 ;
    wire SubBytesIns_Inst_Sbox_1_T19 ;
    wire SubBytesIns_Inst_Sbox_1_T18 ;
    wire SubBytesIns_Inst_Sbox_1_T17 ;
    wire SubBytesIns_Inst_Sbox_1_T16 ;
    wire SubBytesIns_Inst_Sbox_1_T15 ;
    wire SubBytesIns_Inst_Sbox_1_T14 ;
    wire SubBytesIns_Inst_Sbox_1_T13 ;
    wire SubBytesIns_Inst_Sbox_1_T12 ;
    wire SubBytesIns_Inst_Sbox_1_T11 ;
    wire SubBytesIns_Inst_Sbox_1_T10 ;
    wire SubBytesIns_Inst_Sbox_1_T9 ;
    wire SubBytesIns_Inst_Sbox_1_T8 ;
    wire SubBytesIns_Inst_Sbox_1_T7 ;
    wire SubBytesIns_Inst_Sbox_1_T6 ;
    wire SubBytesIns_Inst_Sbox_1_T5 ;
    wire SubBytesIns_Inst_Sbox_1_T4 ;
    wire SubBytesIns_Inst_Sbox_1_T3 ;
    wire SubBytesIns_Inst_Sbox_1_T2 ;
    wire SubBytesIns_Inst_Sbox_1_T1 ;
    wire SubBytesIns_Inst_Sbox_2_L29 ;
    wire SubBytesIns_Inst_Sbox_2_L28 ;
    wire SubBytesIns_Inst_Sbox_2_L27 ;
    wire SubBytesIns_Inst_Sbox_2_L26 ;
    wire SubBytesIns_Inst_Sbox_2_L25 ;
    wire SubBytesIns_Inst_Sbox_2_L24 ;
    wire SubBytesIns_Inst_Sbox_2_L23 ;
    wire SubBytesIns_Inst_Sbox_2_L22 ;
    wire SubBytesIns_Inst_Sbox_2_L21 ;
    wire SubBytesIns_Inst_Sbox_2_L20 ;
    wire SubBytesIns_Inst_Sbox_2_L19 ;
    wire SubBytesIns_Inst_Sbox_2_L18 ;
    wire SubBytesIns_Inst_Sbox_2_L17 ;
    wire SubBytesIns_Inst_Sbox_2_L16 ;
    wire SubBytesIns_Inst_Sbox_2_L15 ;
    wire SubBytesIns_Inst_Sbox_2_L14 ;
    wire SubBytesIns_Inst_Sbox_2_L13 ;
    wire SubBytesIns_Inst_Sbox_2_L12 ;
    wire SubBytesIns_Inst_Sbox_2_L11 ;
    wire SubBytesIns_Inst_Sbox_2_L10 ;
    wire SubBytesIns_Inst_Sbox_2_L9 ;
    wire SubBytesIns_Inst_Sbox_2_L8 ;
    wire SubBytesIns_Inst_Sbox_2_L7 ;
    wire SubBytesIns_Inst_Sbox_2_L6 ;
    wire SubBytesIns_Inst_Sbox_2_L5 ;
    wire SubBytesIns_Inst_Sbox_2_L4 ;
    wire SubBytesIns_Inst_Sbox_2_L3 ;
    wire SubBytesIns_Inst_Sbox_2_L2 ;
    wire SubBytesIns_Inst_Sbox_2_L1 ;
    wire SubBytesIns_Inst_Sbox_2_L0 ;
    wire SubBytesIns_Inst_Sbox_2_M63 ;
    wire SubBytesIns_Inst_Sbox_2_M62 ;
    wire SubBytesIns_Inst_Sbox_2_M61 ;
    wire SubBytesIns_Inst_Sbox_2_M60 ;
    wire SubBytesIns_Inst_Sbox_2_M59 ;
    wire SubBytesIns_Inst_Sbox_2_M58 ;
    wire SubBytesIns_Inst_Sbox_2_M57 ;
    wire SubBytesIns_Inst_Sbox_2_M56 ;
    wire SubBytesIns_Inst_Sbox_2_M55 ;
    wire SubBytesIns_Inst_Sbox_2_M54 ;
    wire SubBytesIns_Inst_Sbox_2_M53 ;
    wire SubBytesIns_Inst_Sbox_2_M52 ;
    wire SubBytesIns_Inst_Sbox_2_M51 ;
    wire SubBytesIns_Inst_Sbox_2_M50 ;
    wire SubBytesIns_Inst_Sbox_2_M49 ;
    wire SubBytesIns_Inst_Sbox_2_M48 ;
    wire SubBytesIns_Inst_Sbox_2_M47 ;
    wire SubBytesIns_Inst_Sbox_2_M46 ;
    wire SubBytesIns_Inst_Sbox_2_M45 ;
    wire SubBytesIns_Inst_Sbox_2_M44 ;
    wire SubBytesIns_Inst_Sbox_2_M43 ;
    wire SubBytesIns_Inst_Sbox_2_M42 ;
    wire SubBytesIns_Inst_Sbox_2_M41 ;
    wire SubBytesIns_Inst_Sbox_2_M40 ;
    wire SubBytesIns_Inst_Sbox_2_M39 ;
    wire SubBytesIns_Inst_Sbox_2_M38 ;
    wire SubBytesIns_Inst_Sbox_2_M37 ;
    wire SubBytesIns_Inst_Sbox_2_M36 ;
    wire SubBytesIns_Inst_Sbox_2_M35 ;
    wire SubBytesIns_Inst_Sbox_2_M34 ;
    wire SubBytesIns_Inst_Sbox_2_M33 ;
    wire SubBytesIns_Inst_Sbox_2_M32 ;
    wire SubBytesIns_Inst_Sbox_2_M31 ;
    wire SubBytesIns_Inst_Sbox_2_M30 ;
    wire SubBytesIns_Inst_Sbox_2_M29 ;
    wire SubBytesIns_Inst_Sbox_2_M28 ;
    wire SubBytesIns_Inst_Sbox_2_M27 ;
    wire SubBytesIns_Inst_Sbox_2_M26 ;
    wire SubBytesIns_Inst_Sbox_2_M25 ;
    wire SubBytesIns_Inst_Sbox_2_M24 ;
    wire SubBytesIns_Inst_Sbox_2_M23 ;
    wire SubBytesIns_Inst_Sbox_2_M22 ;
    wire SubBytesIns_Inst_Sbox_2_M21 ;
    wire SubBytesIns_Inst_Sbox_2_M20 ;
    wire SubBytesIns_Inst_Sbox_2_M19 ;
    wire SubBytesIns_Inst_Sbox_2_M18 ;
    wire SubBytesIns_Inst_Sbox_2_M17 ;
    wire SubBytesIns_Inst_Sbox_2_M16 ;
    wire SubBytesIns_Inst_Sbox_2_M15 ;
    wire SubBytesIns_Inst_Sbox_2_M14 ;
    wire SubBytesIns_Inst_Sbox_2_M13 ;
    wire SubBytesIns_Inst_Sbox_2_M12 ;
    wire SubBytesIns_Inst_Sbox_2_M11 ;
    wire SubBytesIns_Inst_Sbox_2_M10 ;
    wire SubBytesIns_Inst_Sbox_2_M9 ;
    wire SubBytesIns_Inst_Sbox_2_M8 ;
    wire SubBytesIns_Inst_Sbox_2_M7 ;
    wire SubBytesIns_Inst_Sbox_2_M6 ;
    wire SubBytesIns_Inst_Sbox_2_M5 ;
    wire SubBytesIns_Inst_Sbox_2_M4 ;
    wire SubBytesIns_Inst_Sbox_2_M3 ;
    wire SubBytesIns_Inst_Sbox_2_M2 ;
    wire SubBytesIns_Inst_Sbox_2_M1 ;
    wire SubBytesIns_Inst_Sbox_2_T27 ;
    wire SubBytesIns_Inst_Sbox_2_T26 ;
    wire SubBytesIns_Inst_Sbox_2_T25 ;
    wire SubBytesIns_Inst_Sbox_2_T24 ;
    wire SubBytesIns_Inst_Sbox_2_T23 ;
    wire SubBytesIns_Inst_Sbox_2_T22 ;
    wire SubBytesIns_Inst_Sbox_2_T21 ;
    wire SubBytesIns_Inst_Sbox_2_T20 ;
    wire SubBytesIns_Inst_Sbox_2_T19 ;
    wire SubBytesIns_Inst_Sbox_2_T18 ;
    wire SubBytesIns_Inst_Sbox_2_T17 ;
    wire SubBytesIns_Inst_Sbox_2_T16 ;
    wire SubBytesIns_Inst_Sbox_2_T15 ;
    wire SubBytesIns_Inst_Sbox_2_T14 ;
    wire SubBytesIns_Inst_Sbox_2_T13 ;
    wire SubBytesIns_Inst_Sbox_2_T12 ;
    wire SubBytesIns_Inst_Sbox_2_T11 ;
    wire SubBytesIns_Inst_Sbox_2_T10 ;
    wire SubBytesIns_Inst_Sbox_2_T9 ;
    wire SubBytesIns_Inst_Sbox_2_T8 ;
    wire SubBytesIns_Inst_Sbox_2_T7 ;
    wire SubBytesIns_Inst_Sbox_2_T6 ;
    wire SubBytesIns_Inst_Sbox_2_T5 ;
    wire SubBytesIns_Inst_Sbox_2_T4 ;
    wire SubBytesIns_Inst_Sbox_2_T3 ;
    wire SubBytesIns_Inst_Sbox_2_T2 ;
    wire SubBytesIns_Inst_Sbox_2_T1 ;
    wire SubBytesIns_Inst_Sbox_3_L29 ;
    wire SubBytesIns_Inst_Sbox_3_L28 ;
    wire SubBytesIns_Inst_Sbox_3_L27 ;
    wire SubBytesIns_Inst_Sbox_3_L26 ;
    wire SubBytesIns_Inst_Sbox_3_L25 ;
    wire SubBytesIns_Inst_Sbox_3_L24 ;
    wire SubBytesIns_Inst_Sbox_3_L23 ;
    wire SubBytesIns_Inst_Sbox_3_L22 ;
    wire SubBytesIns_Inst_Sbox_3_L21 ;
    wire SubBytesIns_Inst_Sbox_3_L20 ;
    wire SubBytesIns_Inst_Sbox_3_L19 ;
    wire SubBytesIns_Inst_Sbox_3_L18 ;
    wire SubBytesIns_Inst_Sbox_3_L17 ;
    wire SubBytesIns_Inst_Sbox_3_L16 ;
    wire SubBytesIns_Inst_Sbox_3_L15 ;
    wire SubBytesIns_Inst_Sbox_3_L14 ;
    wire SubBytesIns_Inst_Sbox_3_L13 ;
    wire SubBytesIns_Inst_Sbox_3_L12 ;
    wire SubBytesIns_Inst_Sbox_3_L11 ;
    wire SubBytesIns_Inst_Sbox_3_L10 ;
    wire SubBytesIns_Inst_Sbox_3_L9 ;
    wire SubBytesIns_Inst_Sbox_3_L8 ;
    wire SubBytesIns_Inst_Sbox_3_L7 ;
    wire SubBytesIns_Inst_Sbox_3_L6 ;
    wire SubBytesIns_Inst_Sbox_3_L5 ;
    wire SubBytesIns_Inst_Sbox_3_L4 ;
    wire SubBytesIns_Inst_Sbox_3_L3 ;
    wire SubBytesIns_Inst_Sbox_3_L2 ;
    wire SubBytesIns_Inst_Sbox_3_L1 ;
    wire SubBytesIns_Inst_Sbox_3_L0 ;
    wire SubBytesIns_Inst_Sbox_3_M63 ;
    wire SubBytesIns_Inst_Sbox_3_M62 ;
    wire SubBytesIns_Inst_Sbox_3_M61 ;
    wire SubBytesIns_Inst_Sbox_3_M60 ;
    wire SubBytesIns_Inst_Sbox_3_M59 ;
    wire SubBytesIns_Inst_Sbox_3_M58 ;
    wire SubBytesIns_Inst_Sbox_3_M57 ;
    wire SubBytesIns_Inst_Sbox_3_M56 ;
    wire SubBytesIns_Inst_Sbox_3_M55 ;
    wire SubBytesIns_Inst_Sbox_3_M54 ;
    wire SubBytesIns_Inst_Sbox_3_M53 ;
    wire SubBytesIns_Inst_Sbox_3_M52 ;
    wire SubBytesIns_Inst_Sbox_3_M51 ;
    wire SubBytesIns_Inst_Sbox_3_M50 ;
    wire SubBytesIns_Inst_Sbox_3_M49 ;
    wire SubBytesIns_Inst_Sbox_3_M48 ;
    wire SubBytesIns_Inst_Sbox_3_M47 ;
    wire SubBytesIns_Inst_Sbox_3_M46 ;
    wire SubBytesIns_Inst_Sbox_3_M45 ;
    wire SubBytesIns_Inst_Sbox_3_M44 ;
    wire SubBytesIns_Inst_Sbox_3_M43 ;
    wire SubBytesIns_Inst_Sbox_3_M42 ;
    wire SubBytesIns_Inst_Sbox_3_M41 ;
    wire SubBytesIns_Inst_Sbox_3_M40 ;
    wire SubBytesIns_Inst_Sbox_3_M39 ;
    wire SubBytesIns_Inst_Sbox_3_M38 ;
    wire SubBytesIns_Inst_Sbox_3_M37 ;
    wire SubBytesIns_Inst_Sbox_3_M36 ;
    wire SubBytesIns_Inst_Sbox_3_M35 ;
    wire SubBytesIns_Inst_Sbox_3_M34 ;
    wire SubBytesIns_Inst_Sbox_3_M33 ;
    wire SubBytesIns_Inst_Sbox_3_M32 ;
    wire SubBytesIns_Inst_Sbox_3_M31 ;
    wire SubBytesIns_Inst_Sbox_3_M30 ;
    wire SubBytesIns_Inst_Sbox_3_M29 ;
    wire SubBytesIns_Inst_Sbox_3_M28 ;
    wire SubBytesIns_Inst_Sbox_3_M27 ;
    wire SubBytesIns_Inst_Sbox_3_M26 ;
    wire SubBytesIns_Inst_Sbox_3_M25 ;
    wire SubBytesIns_Inst_Sbox_3_M24 ;
    wire SubBytesIns_Inst_Sbox_3_M23 ;
    wire SubBytesIns_Inst_Sbox_3_M22 ;
    wire SubBytesIns_Inst_Sbox_3_M21 ;
    wire SubBytesIns_Inst_Sbox_3_M20 ;
    wire SubBytesIns_Inst_Sbox_3_M19 ;
    wire SubBytesIns_Inst_Sbox_3_M18 ;
    wire SubBytesIns_Inst_Sbox_3_M17 ;
    wire SubBytesIns_Inst_Sbox_3_M16 ;
    wire SubBytesIns_Inst_Sbox_3_M15 ;
    wire SubBytesIns_Inst_Sbox_3_M14 ;
    wire SubBytesIns_Inst_Sbox_3_M13 ;
    wire SubBytesIns_Inst_Sbox_3_M12 ;
    wire SubBytesIns_Inst_Sbox_3_M11 ;
    wire SubBytesIns_Inst_Sbox_3_M10 ;
    wire SubBytesIns_Inst_Sbox_3_M9 ;
    wire SubBytesIns_Inst_Sbox_3_M8 ;
    wire SubBytesIns_Inst_Sbox_3_M7 ;
    wire SubBytesIns_Inst_Sbox_3_M6 ;
    wire SubBytesIns_Inst_Sbox_3_M5 ;
    wire SubBytesIns_Inst_Sbox_3_M4 ;
    wire SubBytesIns_Inst_Sbox_3_M3 ;
    wire SubBytesIns_Inst_Sbox_3_M2 ;
    wire SubBytesIns_Inst_Sbox_3_M1 ;
    wire SubBytesIns_Inst_Sbox_3_T27 ;
    wire SubBytesIns_Inst_Sbox_3_T26 ;
    wire SubBytesIns_Inst_Sbox_3_T25 ;
    wire SubBytesIns_Inst_Sbox_3_T24 ;
    wire SubBytesIns_Inst_Sbox_3_T23 ;
    wire SubBytesIns_Inst_Sbox_3_T22 ;
    wire SubBytesIns_Inst_Sbox_3_T21 ;
    wire SubBytesIns_Inst_Sbox_3_T20 ;
    wire SubBytesIns_Inst_Sbox_3_T19 ;
    wire SubBytesIns_Inst_Sbox_3_T18 ;
    wire SubBytesIns_Inst_Sbox_3_T17 ;
    wire SubBytesIns_Inst_Sbox_3_T16 ;
    wire SubBytesIns_Inst_Sbox_3_T15 ;
    wire SubBytesIns_Inst_Sbox_3_T14 ;
    wire SubBytesIns_Inst_Sbox_3_T13 ;
    wire SubBytesIns_Inst_Sbox_3_T12 ;
    wire SubBytesIns_Inst_Sbox_3_T11 ;
    wire SubBytesIns_Inst_Sbox_3_T10 ;
    wire SubBytesIns_Inst_Sbox_3_T9 ;
    wire SubBytesIns_Inst_Sbox_3_T8 ;
    wire SubBytesIns_Inst_Sbox_3_T7 ;
    wire SubBytesIns_Inst_Sbox_3_T6 ;
    wire SubBytesIns_Inst_Sbox_3_T5 ;
    wire SubBytesIns_Inst_Sbox_3_T4 ;
    wire SubBytesIns_Inst_Sbox_3_T3 ;
    wire SubBytesIns_Inst_Sbox_3_T2 ;
    wire SubBytesIns_Inst_Sbox_3_T1 ;
    wire SubBytesIns_Inst_Sbox_4_L29 ;
    wire SubBytesIns_Inst_Sbox_4_L28 ;
    wire SubBytesIns_Inst_Sbox_4_L27 ;
    wire SubBytesIns_Inst_Sbox_4_L26 ;
    wire SubBytesIns_Inst_Sbox_4_L25 ;
    wire SubBytesIns_Inst_Sbox_4_L24 ;
    wire SubBytesIns_Inst_Sbox_4_L23 ;
    wire SubBytesIns_Inst_Sbox_4_L22 ;
    wire SubBytesIns_Inst_Sbox_4_L21 ;
    wire SubBytesIns_Inst_Sbox_4_L20 ;
    wire SubBytesIns_Inst_Sbox_4_L19 ;
    wire SubBytesIns_Inst_Sbox_4_L18 ;
    wire SubBytesIns_Inst_Sbox_4_L17 ;
    wire SubBytesIns_Inst_Sbox_4_L16 ;
    wire SubBytesIns_Inst_Sbox_4_L15 ;
    wire SubBytesIns_Inst_Sbox_4_L14 ;
    wire SubBytesIns_Inst_Sbox_4_L13 ;
    wire SubBytesIns_Inst_Sbox_4_L12 ;
    wire SubBytesIns_Inst_Sbox_4_L11 ;
    wire SubBytesIns_Inst_Sbox_4_L10 ;
    wire SubBytesIns_Inst_Sbox_4_L9 ;
    wire SubBytesIns_Inst_Sbox_4_L8 ;
    wire SubBytesIns_Inst_Sbox_4_L7 ;
    wire SubBytesIns_Inst_Sbox_4_L6 ;
    wire SubBytesIns_Inst_Sbox_4_L5 ;
    wire SubBytesIns_Inst_Sbox_4_L4 ;
    wire SubBytesIns_Inst_Sbox_4_L3 ;
    wire SubBytesIns_Inst_Sbox_4_L2 ;
    wire SubBytesIns_Inst_Sbox_4_L1 ;
    wire SubBytesIns_Inst_Sbox_4_L0 ;
    wire SubBytesIns_Inst_Sbox_4_M63 ;
    wire SubBytesIns_Inst_Sbox_4_M62 ;
    wire SubBytesIns_Inst_Sbox_4_M61 ;
    wire SubBytesIns_Inst_Sbox_4_M60 ;
    wire SubBytesIns_Inst_Sbox_4_M59 ;
    wire SubBytesIns_Inst_Sbox_4_M58 ;
    wire SubBytesIns_Inst_Sbox_4_M57 ;
    wire SubBytesIns_Inst_Sbox_4_M56 ;
    wire SubBytesIns_Inst_Sbox_4_M55 ;
    wire SubBytesIns_Inst_Sbox_4_M54 ;
    wire SubBytesIns_Inst_Sbox_4_M53 ;
    wire SubBytesIns_Inst_Sbox_4_M52 ;
    wire SubBytesIns_Inst_Sbox_4_M51 ;
    wire SubBytesIns_Inst_Sbox_4_M50 ;
    wire SubBytesIns_Inst_Sbox_4_M49 ;
    wire SubBytesIns_Inst_Sbox_4_M48 ;
    wire SubBytesIns_Inst_Sbox_4_M47 ;
    wire SubBytesIns_Inst_Sbox_4_M46 ;
    wire SubBytesIns_Inst_Sbox_4_M45 ;
    wire SubBytesIns_Inst_Sbox_4_M44 ;
    wire SubBytesIns_Inst_Sbox_4_M43 ;
    wire SubBytesIns_Inst_Sbox_4_M42 ;
    wire SubBytesIns_Inst_Sbox_4_M41 ;
    wire SubBytesIns_Inst_Sbox_4_M40 ;
    wire SubBytesIns_Inst_Sbox_4_M39 ;
    wire SubBytesIns_Inst_Sbox_4_M38 ;
    wire SubBytesIns_Inst_Sbox_4_M37 ;
    wire SubBytesIns_Inst_Sbox_4_M36 ;
    wire SubBytesIns_Inst_Sbox_4_M35 ;
    wire SubBytesIns_Inst_Sbox_4_M34 ;
    wire SubBytesIns_Inst_Sbox_4_M33 ;
    wire SubBytesIns_Inst_Sbox_4_M32 ;
    wire SubBytesIns_Inst_Sbox_4_M31 ;
    wire SubBytesIns_Inst_Sbox_4_M30 ;
    wire SubBytesIns_Inst_Sbox_4_M29 ;
    wire SubBytesIns_Inst_Sbox_4_M28 ;
    wire SubBytesIns_Inst_Sbox_4_M27 ;
    wire SubBytesIns_Inst_Sbox_4_M26 ;
    wire SubBytesIns_Inst_Sbox_4_M25 ;
    wire SubBytesIns_Inst_Sbox_4_M24 ;
    wire SubBytesIns_Inst_Sbox_4_M23 ;
    wire SubBytesIns_Inst_Sbox_4_M22 ;
    wire SubBytesIns_Inst_Sbox_4_M21 ;
    wire SubBytesIns_Inst_Sbox_4_M20 ;
    wire SubBytesIns_Inst_Sbox_4_M19 ;
    wire SubBytesIns_Inst_Sbox_4_M18 ;
    wire SubBytesIns_Inst_Sbox_4_M17 ;
    wire SubBytesIns_Inst_Sbox_4_M16 ;
    wire SubBytesIns_Inst_Sbox_4_M15 ;
    wire SubBytesIns_Inst_Sbox_4_M14 ;
    wire SubBytesIns_Inst_Sbox_4_M13 ;
    wire SubBytesIns_Inst_Sbox_4_M12 ;
    wire SubBytesIns_Inst_Sbox_4_M11 ;
    wire SubBytesIns_Inst_Sbox_4_M10 ;
    wire SubBytesIns_Inst_Sbox_4_M9 ;
    wire SubBytesIns_Inst_Sbox_4_M8 ;
    wire SubBytesIns_Inst_Sbox_4_M7 ;
    wire SubBytesIns_Inst_Sbox_4_M6 ;
    wire SubBytesIns_Inst_Sbox_4_M5 ;
    wire SubBytesIns_Inst_Sbox_4_M4 ;
    wire SubBytesIns_Inst_Sbox_4_M3 ;
    wire SubBytesIns_Inst_Sbox_4_M2 ;
    wire SubBytesIns_Inst_Sbox_4_M1 ;
    wire SubBytesIns_Inst_Sbox_4_T27 ;
    wire SubBytesIns_Inst_Sbox_4_T26 ;
    wire SubBytesIns_Inst_Sbox_4_T25 ;
    wire SubBytesIns_Inst_Sbox_4_T24 ;
    wire SubBytesIns_Inst_Sbox_4_T23 ;
    wire SubBytesIns_Inst_Sbox_4_T22 ;
    wire SubBytesIns_Inst_Sbox_4_T21 ;
    wire SubBytesIns_Inst_Sbox_4_T20 ;
    wire SubBytesIns_Inst_Sbox_4_T19 ;
    wire SubBytesIns_Inst_Sbox_4_T18 ;
    wire SubBytesIns_Inst_Sbox_4_T17 ;
    wire SubBytesIns_Inst_Sbox_4_T16 ;
    wire SubBytesIns_Inst_Sbox_4_T15 ;
    wire SubBytesIns_Inst_Sbox_4_T14 ;
    wire SubBytesIns_Inst_Sbox_4_T13 ;
    wire SubBytesIns_Inst_Sbox_4_T12 ;
    wire SubBytesIns_Inst_Sbox_4_T11 ;
    wire SubBytesIns_Inst_Sbox_4_T10 ;
    wire SubBytesIns_Inst_Sbox_4_T9 ;
    wire SubBytesIns_Inst_Sbox_4_T8 ;
    wire SubBytesIns_Inst_Sbox_4_T7 ;
    wire SubBytesIns_Inst_Sbox_4_T6 ;
    wire SubBytesIns_Inst_Sbox_4_T5 ;
    wire SubBytesIns_Inst_Sbox_4_T4 ;
    wire SubBytesIns_Inst_Sbox_4_T3 ;
    wire SubBytesIns_Inst_Sbox_4_T2 ;
    wire SubBytesIns_Inst_Sbox_4_T1 ;
    wire SubBytesIns_Inst_Sbox_5_L29 ;
    wire SubBytesIns_Inst_Sbox_5_L28 ;
    wire SubBytesIns_Inst_Sbox_5_L27 ;
    wire SubBytesIns_Inst_Sbox_5_L26 ;
    wire SubBytesIns_Inst_Sbox_5_L25 ;
    wire SubBytesIns_Inst_Sbox_5_L24 ;
    wire SubBytesIns_Inst_Sbox_5_L23 ;
    wire SubBytesIns_Inst_Sbox_5_L22 ;
    wire SubBytesIns_Inst_Sbox_5_L21 ;
    wire SubBytesIns_Inst_Sbox_5_L20 ;
    wire SubBytesIns_Inst_Sbox_5_L19 ;
    wire SubBytesIns_Inst_Sbox_5_L18 ;
    wire SubBytesIns_Inst_Sbox_5_L17 ;
    wire SubBytesIns_Inst_Sbox_5_L16 ;
    wire SubBytesIns_Inst_Sbox_5_L15 ;
    wire SubBytesIns_Inst_Sbox_5_L14 ;
    wire SubBytesIns_Inst_Sbox_5_L13 ;
    wire SubBytesIns_Inst_Sbox_5_L12 ;
    wire SubBytesIns_Inst_Sbox_5_L11 ;
    wire SubBytesIns_Inst_Sbox_5_L10 ;
    wire SubBytesIns_Inst_Sbox_5_L9 ;
    wire SubBytesIns_Inst_Sbox_5_L8 ;
    wire SubBytesIns_Inst_Sbox_5_L7 ;
    wire SubBytesIns_Inst_Sbox_5_L6 ;
    wire SubBytesIns_Inst_Sbox_5_L5 ;
    wire SubBytesIns_Inst_Sbox_5_L4 ;
    wire SubBytesIns_Inst_Sbox_5_L3 ;
    wire SubBytesIns_Inst_Sbox_5_L2 ;
    wire SubBytesIns_Inst_Sbox_5_L1 ;
    wire SubBytesIns_Inst_Sbox_5_L0 ;
    wire SubBytesIns_Inst_Sbox_5_M63 ;
    wire SubBytesIns_Inst_Sbox_5_M62 ;
    wire SubBytesIns_Inst_Sbox_5_M61 ;
    wire SubBytesIns_Inst_Sbox_5_M60 ;
    wire SubBytesIns_Inst_Sbox_5_M59 ;
    wire SubBytesIns_Inst_Sbox_5_M58 ;
    wire SubBytesIns_Inst_Sbox_5_M57 ;
    wire SubBytesIns_Inst_Sbox_5_M56 ;
    wire SubBytesIns_Inst_Sbox_5_M55 ;
    wire SubBytesIns_Inst_Sbox_5_M54 ;
    wire SubBytesIns_Inst_Sbox_5_M53 ;
    wire SubBytesIns_Inst_Sbox_5_M52 ;
    wire SubBytesIns_Inst_Sbox_5_M51 ;
    wire SubBytesIns_Inst_Sbox_5_M50 ;
    wire SubBytesIns_Inst_Sbox_5_M49 ;
    wire SubBytesIns_Inst_Sbox_5_M48 ;
    wire SubBytesIns_Inst_Sbox_5_M47 ;
    wire SubBytesIns_Inst_Sbox_5_M46 ;
    wire SubBytesIns_Inst_Sbox_5_M45 ;
    wire SubBytesIns_Inst_Sbox_5_M44 ;
    wire SubBytesIns_Inst_Sbox_5_M43 ;
    wire SubBytesIns_Inst_Sbox_5_M42 ;
    wire SubBytesIns_Inst_Sbox_5_M41 ;
    wire SubBytesIns_Inst_Sbox_5_M40 ;
    wire SubBytesIns_Inst_Sbox_5_M39 ;
    wire SubBytesIns_Inst_Sbox_5_M38 ;
    wire SubBytesIns_Inst_Sbox_5_M37 ;
    wire SubBytesIns_Inst_Sbox_5_M36 ;
    wire SubBytesIns_Inst_Sbox_5_M35 ;
    wire SubBytesIns_Inst_Sbox_5_M34 ;
    wire SubBytesIns_Inst_Sbox_5_M33 ;
    wire SubBytesIns_Inst_Sbox_5_M32 ;
    wire SubBytesIns_Inst_Sbox_5_M31 ;
    wire SubBytesIns_Inst_Sbox_5_M30 ;
    wire SubBytesIns_Inst_Sbox_5_M29 ;
    wire SubBytesIns_Inst_Sbox_5_M28 ;
    wire SubBytesIns_Inst_Sbox_5_M27 ;
    wire SubBytesIns_Inst_Sbox_5_M26 ;
    wire SubBytesIns_Inst_Sbox_5_M25 ;
    wire SubBytesIns_Inst_Sbox_5_M24 ;
    wire SubBytesIns_Inst_Sbox_5_M23 ;
    wire SubBytesIns_Inst_Sbox_5_M22 ;
    wire SubBytesIns_Inst_Sbox_5_M21 ;
    wire SubBytesIns_Inst_Sbox_5_M20 ;
    wire SubBytesIns_Inst_Sbox_5_M19 ;
    wire SubBytesIns_Inst_Sbox_5_M18 ;
    wire SubBytesIns_Inst_Sbox_5_M17 ;
    wire SubBytesIns_Inst_Sbox_5_M16 ;
    wire SubBytesIns_Inst_Sbox_5_M15 ;
    wire SubBytesIns_Inst_Sbox_5_M14 ;
    wire SubBytesIns_Inst_Sbox_5_M13 ;
    wire SubBytesIns_Inst_Sbox_5_M12 ;
    wire SubBytesIns_Inst_Sbox_5_M11 ;
    wire SubBytesIns_Inst_Sbox_5_M10 ;
    wire SubBytesIns_Inst_Sbox_5_M9 ;
    wire SubBytesIns_Inst_Sbox_5_M8 ;
    wire SubBytesIns_Inst_Sbox_5_M7 ;
    wire SubBytesIns_Inst_Sbox_5_M6 ;
    wire SubBytesIns_Inst_Sbox_5_M5 ;
    wire SubBytesIns_Inst_Sbox_5_M4 ;
    wire SubBytesIns_Inst_Sbox_5_M3 ;
    wire SubBytesIns_Inst_Sbox_5_M2 ;
    wire SubBytesIns_Inst_Sbox_5_M1 ;
    wire SubBytesIns_Inst_Sbox_5_T27 ;
    wire SubBytesIns_Inst_Sbox_5_T26 ;
    wire SubBytesIns_Inst_Sbox_5_T25 ;
    wire SubBytesIns_Inst_Sbox_5_T24 ;
    wire SubBytesIns_Inst_Sbox_5_T23 ;
    wire SubBytesIns_Inst_Sbox_5_T22 ;
    wire SubBytesIns_Inst_Sbox_5_T21 ;
    wire SubBytesIns_Inst_Sbox_5_T20 ;
    wire SubBytesIns_Inst_Sbox_5_T19 ;
    wire SubBytesIns_Inst_Sbox_5_T18 ;
    wire SubBytesIns_Inst_Sbox_5_T17 ;
    wire SubBytesIns_Inst_Sbox_5_T16 ;
    wire SubBytesIns_Inst_Sbox_5_T15 ;
    wire SubBytesIns_Inst_Sbox_5_T14 ;
    wire SubBytesIns_Inst_Sbox_5_T13 ;
    wire SubBytesIns_Inst_Sbox_5_T12 ;
    wire SubBytesIns_Inst_Sbox_5_T11 ;
    wire SubBytesIns_Inst_Sbox_5_T10 ;
    wire SubBytesIns_Inst_Sbox_5_T9 ;
    wire SubBytesIns_Inst_Sbox_5_T8 ;
    wire SubBytesIns_Inst_Sbox_5_T7 ;
    wire SubBytesIns_Inst_Sbox_5_T6 ;
    wire SubBytesIns_Inst_Sbox_5_T5 ;
    wire SubBytesIns_Inst_Sbox_5_T4 ;
    wire SubBytesIns_Inst_Sbox_5_T3 ;
    wire SubBytesIns_Inst_Sbox_5_T2 ;
    wire SubBytesIns_Inst_Sbox_5_T1 ;
    wire SubBytesIns_Inst_Sbox_6_L29 ;
    wire SubBytesIns_Inst_Sbox_6_L28 ;
    wire SubBytesIns_Inst_Sbox_6_L27 ;
    wire SubBytesIns_Inst_Sbox_6_L26 ;
    wire SubBytesIns_Inst_Sbox_6_L25 ;
    wire SubBytesIns_Inst_Sbox_6_L24 ;
    wire SubBytesIns_Inst_Sbox_6_L23 ;
    wire SubBytesIns_Inst_Sbox_6_L22 ;
    wire SubBytesIns_Inst_Sbox_6_L21 ;
    wire SubBytesIns_Inst_Sbox_6_L20 ;
    wire SubBytesIns_Inst_Sbox_6_L19 ;
    wire SubBytesIns_Inst_Sbox_6_L18 ;
    wire SubBytesIns_Inst_Sbox_6_L17 ;
    wire SubBytesIns_Inst_Sbox_6_L16 ;
    wire SubBytesIns_Inst_Sbox_6_L15 ;
    wire SubBytesIns_Inst_Sbox_6_L14 ;
    wire SubBytesIns_Inst_Sbox_6_L13 ;
    wire SubBytesIns_Inst_Sbox_6_L12 ;
    wire SubBytesIns_Inst_Sbox_6_L11 ;
    wire SubBytesIns_Inst_Sbox_6_L10 ;
    wire SubBytesIns_Inst_Sbox_6_L9 ;
    wire SubBytesIns_Inst_Sbox_6_L8 ;
    wire SubBytesIns_Inst_Sbox_6_L7 ;
    wire SubBytesIns_Inst_Sbox_6_L6 ;
    wire SubBytesIns_Inst_Sbox_6_L5 ;
    wire SubBytesIns_Inst_Sbox_6_L4 ;
    wire SubBytesIns_Inst_Sbox_6_L3 ;
    wire SubBytesIns_Inst_Sbox_6_L2 ;
    wire SubBytesIns_Inst_Sbox_6_L1 ;
    wire SubBytesIns_Inst_Sbox_6_L0 ;
    wire SubBytesIns_Inst_Sbox_6_M63 ;
    wire SubBytesIns_Inst_Sbox_6_M62 ;
    wire SubBytesIns_Inst_Sbox_6_M61 ;
    wire SubBytesIns_Inst_Sbox_6_M60 ;
    wire SubBytesIns_Inst_Sbox_6_M59 ;
    wire SubBytesIns_Inst_Sbox_6_M58 ;
    wire SubBytesIns_Inst_Sbox_6_M57 ;
    wire SubBytesIns_Inst_Sbox_6_M56 ;
    wire SubBytesIns_Inst_Sbox_6_M55 ;
    wire SubBytesIns_Inst_Sbox_6_M54 ;
    wire SubBytesIns_Inst_Sbox_6_M53 ;
    wire SubBytesIns_Inst_Sbox_6_M52 ;
    wire SubBytesIns_Inst_Sbox_6_M51 ;
    wire SubBytesIns_Inst_Sbox_6_M50 ;
    wire SubBytesIns_Inst_Sbox_6_M49 ;
    wire SubBytesIns_Inst_Sbox_6_M48 ;
    wire SubBytesIns_Inst_Sbox_6_M47 ;
    wire SubBytesIns_Inst_Sbox_6_M46 ;
    wire SubBytesIns_Inst_Sbox_6_M45 ;
    wire SubBytesIns_Inst_Sbox_6_M44 ;
    wire SubBytesIns_Inst_Sbox_6_M43 ;
    wire SubBytesIns_Inst_Sbox_6_M42 ;
    wire SubBytesIns_Inst_Sbox_6_M41 ;
    wire SubBytesIns_Inst_Sbox_6_M40 ;
    wire SubBytesIns_Inst_Sbox_6_M39 ;
    wire SubBytesIns_Inst_Sbox_6_M38 ;
    wire SubBytesIns_Inst_Sbox_6_M37 ;
    wire SubBytesIns_Inst_Sbox_6_M36 ;
    wire SubBytesIns_Inst_Sbox_6_M35 ;
    wire SubBytesIns_Inst_Sbox_6_M34 ;
    wire SubBytesIns_Inst_Sbox_6_M33 ;
    wire SubBytesIns_Inst_Sbox_6_M32 ;
    wire SubBytesIns_Inst_Sbox_6_M31 ;
    wire SubBytesIns_Inst_Sbox_6_M30 ;
    wire SubBytesIns_Inst_Sbox_6_M29 ;
    wire SubBytesIns_Inst_Sbox_6_M28 ;
    wire SubBytesIns_Inst_Sbox_6_M27 ;
    wire SubBytesIns_Inst_Sbox_6_M26 ;
    wire SubBytesIns_Inst_Sbox_6_M25 ;
    wire SubBytesIns_Inst_Sbox_6_M24 ;
    wire SubBytesIns_Inst_Sbox_6_M23 ;
    wire SubBytesIns_Inst_Sbox_6_M22 ;
    wire SubBytesIns_Inst_Sbox_6_M21 ;
    wire SubBytesIns_Inst_Sbox_6_M20 ;
    wire SubBytesIns_Inst_Sbox_6_M19 ;
    wire SubBytesIns_Inst_Sbox_6_M18 ;
    wire SubBytesIns_Inst_Sbox_6_M17 ;
    wire SubBytesIns_Inst_Sbox_6_M16 ;
    wire SubBytesIns_Inst_Sbox_6_M15 ;
    wire SubBytesIns_Inst_Sbox_6_M14 ;
    wire SubBytesIns_Inst_Sbox_6_M13 ;
    wire SubBytesIns_Inst_Sbox_6_M12 ;
    wire SubBytesIns_Inst_Sbox_6_M11 ;
    wire SubBytesIns_Inst_Sbox_6_M10 ;
    wire SubBytesIns_Inst_Sbox_6_M9 ;
    wire SubBytesIns_Inst_Sbox_6_M8 ;
    wire SubBytesIns_Inst_Sbox_6_M7 ;
    wire SubBytesIns_Inst_Sbox_6_M6 ;
    wire SubBytesIns_Inst_Sbox_6_M5 ;
    wire SubBytesIns_Inst_Sbox_6_M4 ;
    wire SubBytesIns_Inst_Sbox_6_M3 ;
    wire SubBytesIns_Inst_Sbox_6_M2 ;
    wire SubBytesIns_Inst_Sbox_6_M1 ;
    wire SubBytesIns_Inst_Sbox_6_T27 ;
    wire SubBytesIns_Inst_Sbox_6_T26 ;
    wire SubBytesIns_Inst_Sbox_6_T25 ;
    wire SubBytesIns_Inst_Sbox_6_T24 ;
    wire SubBytesIns_Inst_Sbox_6_T23 ;
    wire SubBytesIns_Inst_Sbox_6_T22 ;
    wire SubBytesIns_Inst_Sbox_6_T21 ;
    wire SubBytesIns_Inst_Sbox_6_T20 ;
    wire SubBytesIns_Inst_Sbox_6_T19 ;
    wire SubBytesIns_Inst_Sbox_6_T18 ;
    wire SubBytesIns_Inst_Sbox_6_T17 ;
    wire SubBytesIns_Inst_Sbox_6_T16 ;
    wire SubBytesIns_Inst_Sbox_6_T15 ;
    wire SubBytesIns_Inst_Sbox_6_T14 ;
    wire SubBytesIns_Inst_Sbox_6_T13 ;
    wire SubBytesIns_Inst_Sbox_6_T12 ;
    wire SubBytesIns_Inst_Sbox_6_T11 ;
    wire SubBytesIns_Inst_Sbox_6_T10 ;
    wire SubBytesIns_Inst_Sbox_6_T9 ;
    wire SubBytesIns_Inst_Sbox_6_T8 ;
    wire SubBytesIns_Inst_Sbox_6_T7 ;
    wire SubBytesIns_Inst_Sbox_6_T6 ;
    wire SubBytesIns_Inst_Sbox_6_T5 ;
    wire SubBytesIns_Inst_Sbox_6_T4 ;
    wire SubBytesIns_Inst_Sbox_6_T3 ;
    wire SubBytesIns_Inst_Sbox_6_T2 ;
    wire SubBytesIns_Inst_Sbox_6_T1 ;
    wire SubBytesIns_Inst_Sbox_7_L29 ;
    wire SubBytesIns_Inst_Sbox_7_L28 ;
    wire SubBytesIns_Inst_Sbox_7_L27 ;
    wire SubBytesIns_Inst_Sbox_7_L26 ;
    wire SubBytesIns_Inst_Sbox_7_L25 ;
    wire SubBytesIns_Inst_Sbox_7_L24 ;
    wire SubBytesIns_Inst_Sbox_7_L23 ;
    wire SubBytesIns_Inst_Sbox_7_L22 ;
    wire SubBytesIns_Inst_Sbox_7_L21 ;
    wire SubBytesIns_Inst_Sbox_7_L20 ;
    wire SubBytesIns_Inst_Sbox_7_L19 ;
    wire SubBytesIns_Inst_Sbox_7_L18 ;
    wire SubBytesIns_Inst_Sbox_7_L17 ;
    wire SubBytesIns_Inst_Sbox_7_L16 ;
    wire SubBytesIns_Inst_Sbox_7_L15 ;
    wire SubBytesIns_Inst_Sbox_7_L14 ;
    wire SubBytesIns_Inst_Sbox_7_L13 ;
    wire SubBytesIns_Inst_Sbox_7_L12 ;
    wire SubBytesIns_Inst_Sbox_7_L11 ;
    wire SubBytesIns_Inst_Sbox_7_L10 ;
    wire SubBytesIns_Inst_Sbox_7_L9 ;
    wire SubBytesIns_Inst_Sbox_7_L8 ;
    wire SubBytesIns_Inst_Sbox_7_L7 ;
    wire SubBytesIns_Inst_Sbox_7_L6 ;
    wire SubBytesIns_Inst_Sbox_7_L5 ;
    wire SubBytesIns_Inst_Sbox_7_L4 ;
    wire SubBytesIns_Inst_Sbox_7_L3 ;
    wire SubBytesIns_Inst_Sbox_7_L2 ;
    wire SubBytesIns_Inst_Sbox_7_L1 ;
    wire SubBytesIns_Inst_Sbox_7_L0 ;
    wire SubBytesIns_Inst_Sbox_7_M63 ;
    wire SubBytesIns_Inst_Sbox_7_M62 ;
    wire SubBytesIns_Inst_Sbox_7_M61 ;
    wire SubBytesIns_Inst_Sbox_7_M60 ;
    wire SubBytesIns_Inst_Sbox_7_M59 ;
    wire SubBytesIns_Inst_Sbox_7_M58 ;
    wire SubBytesIns_Inst_Sbox_7_M57 ;
    wire SubBytesIns_Inst_Sbox_7_M56 ;
    wire SubBytesIns_Inst_Sbox_7_M55 ;
    wire SubBytesIns_Inst_Sbox_7_M54 ;
    wire SubBytesIns_Inst_Sbox_7_M53 ;
    wire SubBytesIns_Inst_Sbox_7_M52 ;
    wire SubBytesIns_Inst_Sbox_7_M51 ;
    wire SubBytesIns_Inst_Sbox_7_M50 ;
    wire SubBytesIns_Inst_Sbox_7_M49 ;
    wire SubBytesIns_Inst_Sbox_7_M48 ;
    wire SubBytesIns_Inst_Sbox_7_M47 ;
    wire SubBytesIns_Inst_Sbox_7_M46 ;
    wire SubBytesIns_Inst_Sbox_7_M45 ;
    wire SubBytesIns_Inst_Sbox_7_M44 ;
    wire SubBytesIns_Inst_Sbox_7_M43 ;
    wire SubBytesIns_Inst_Sbox_7_M42 ;
    wire SubBytesIns_Inst_Sbox_7_M41 ;
    wire SubBytesIns_Inst_Sbox_7_M40 ;
    wire SubBytesIns_Inst_Sbox_7_M39 ;
    wire SubBytesIns_Inst_Sbox_7_M38 ;
    wire SubBytesIns_Inst_Sbox_7_M37 ;
    wire SubBytesIns_Inst_Sbox_7_M36 ;
    wire SubBytesIns_Inst_Sbox_7_M35 ;
    wire SubBytesIns_Inst_Sbox_7_M34 ;
    wire SubBytesIns_Inst_Sbox_7_M33 ;
    wire SubBytesIns_Inst_Sbox_7_M32 ;
    wire SubBytesIns_Inst_Sbox_7_M31 ;
    wire SubBytesIns_Inst_Sbox_7_M30 ;
    wire SubBytesIns_Inst_Sbox_7_M29 ;
    wire SubBytesIns_Inst_Sbox_7_M28 ;
    wire SubBytesIns_Inst_Sbox_7_M27 ;
    wire SubBytesIns_Inst_Sbox_7_M26 ;
    wire SubBytesIns_Inst_Sbox_7_M25 ;
    wire SubBytesIns_Inst_Sbox_7_M24 ;
    wire SubBytesIns_Inst_Sbox_7_M23 ;
    wire SubBytesIns_Inst_Sbox_7_M22 ;
    wire SubBytesIns_Inst_Sbox_7_M21 ;
    wire SubBytesIns_Inst_Sbox_7_M20 ;
    wire SubBytesIns_Inst_Sbox_7_M19 ;
    wire SubBytesIns_Inst_Sbox_7_M18 ;
    wire SubBytesIns_Inst_Sbox_7_M17 ;
    wire SubBytesIns_Inst_Sbox_7_M16 ;
    wire SubBytesIns_Inst_Sbox_7_M15 ;
    wire SubBytesIns_Inst_Sbox_7_M14 ;
    wire SubBytesIns_Inst_Sbox_7_M13 ;
    wire SubBytesIns_Inst_Sbox_7_M12 ;
    wire SubBytesIns_Inst_Sbox_7_M11 ;
    wire SubBytesIns_Inst_Sbox_7_M10 ;
    wire SubBytesIns_Inst_Sbox_7_M9 ;
    wire SubBytesIns_Inst_Sbox_7_M8 ;
    wire SubBytesIns_Inst_Sbox_7_M7 ;
    wire SubBytesIns_Inst_Sbox_7_M6 ;
    wire SubBytesIns_Inst_Sbox_7_M5 ;
    wire SubBytesIns_Inst_Sbox_7_M4 ;
    wire SubBytesIns_Inst_Sbox_7_M3 ;
    wire SubBytesIns_Inst_Sbox_7_M2 ;
    wire SubBytesIns_Inst_Sbox_7_M1 ;
    wire SubBytesIns_Inst_Sbox_7_T27 ;
    wire SubBytesIns_Inst_Sbox_7_T26 ;
    wire SubBytesIns_Inst_Sbox_7_T25 ;
    wire SubBytesIns_Inst_Sbox_7_T24 ;
    wire SubBytesIns_Inst_Sbox_7_T23 ;
    wire SubBytesIns_Inst_Sbox_7_T22 ;
    wire SubBytesIns_Inst_Sbox_7_T21 ;
    wire SubBytesIns_Inst_Sbox_7_T20 ;
    wire SubBytesIns_Inst_Sbox_7_T19 ;
    wire SubBytesIns_Inst_Sbox_7_T18 ;
    wire SubBytesIns_Inst_Sbox_7_T17 ;
    wire SubBytesIns_Inst_Sbox_7_T16 ;
    wire SubBytesIns_Inst_Sbox_7_T15 ;
    wire SubBytesIns_Inst_Sbox_7_T14 ;
    wire SubBytesIns_Inst_Sbox_7_T13 ;
    wire SubBytesIns_Inst_Sbox_7_T12 ;
    wire SubBytesIns_Inst_Sbox_7_T11 ;
    wire SubBytesIns_Inst_Sbox_7_T10 ;
    wire SubBytesIns_Inst_Sbox_7_T9 ;
    wire SubBytesIns_Inst_Sbox_7_T8 ;
    wire SubBytesIns_Inst_Sbox_7_T7 ;
    wire SubBytesIns_Inst_Sbox_7_T6 ;
    wire SubBytesIns_Inst_Sbox_7_T5 ;
    wire SubBytesIns_Inst_Sbox_7_T4 ;
    wire SubBytesIns_Inst_Sbox_7_T3 ;
    wire SubBytesIns_Inst_Sbox_7_T2 ;
    wire SubBytesIns_Inst_Sbox_7_T1 ;
    wire SubBytesIns_Inst_Sbox_8_L29 ;
    wire SubBytesIns_Inst_Sbox_8_L28 ;
    wire SubBytesIns_Inst_Sbox_8_L27 ;
    wire SubBytesIns_Inst_Sbox_8_L26 ;
    wire SubBytesIns_Inst_Sbox_8_L25 ;
    wire SubBytesIns_Inst_Sbox_8_L24 ;
    wire SubBytesIns_Inst_Sbox_8_L23 ;
    wire SubBytesIns_Inst_Sbox_8_L22 ;
    wire SubBytesIns_Inst_Sbox_8_L21 ;
    wire SubBytesIns_Inst_Sbox_8_L20 ;
    wire SubBytesIns_Inst_Sbox_8_L19 ;
    wire SubBytesIns_Inst_Sbox_8_L18 ;
    wire SubBytesIns_Inst_Sbox_8_L17 ;
    wire SubBytesIns_Inst_Sbox_8_L16 ;
    wire SubBytesIns_Inst_Sbox_8_L15 ;
    wire SubBytesIns_Inst_Sbox_8_L14 ;
    wire SubBytesIns_Inst_Sbox_8_L13 ;
    wire SubBytesIns_Inst_Sbox_8_L12 ;
    wire SubBytesIns_Inst_Sbox_8_L11 ;
    wire SubBytesIns_Inst_Sbox_8_L10 ;
    wire SubBytesIns_Inst_Sbox_8_L9 ;
    wire SubBytesIns_Inst_Sbox_8_L8 ;
    wire SubBytesIns_Inst_Sbox_8_L7 ;
    wire SubBytesIns_Inst_Sbox_8_L6 ;
    wire SubBytesIns_Inst_Sbox_8_L5 ;
    wire SubBytesIns_Inst_Sbox_8_L4 ;
    wire SubBytesIns_Inst_Sbox_8_L3 ;
    wire SubBytesIns_Inst_Sbox_8_L2 ;
    wire SubBytesIns_Inst_Sbox_8_L1 ;
    wire SubBytesIns_Inst_Sbox_8_L0 ;
    wire SubBytesIns_Inst_Sbox_8_M63 ;
    wire SubBytesIns_Inst_Sbox_8_M62 ;
    wire SubBytesIns_Inst_Sbox_8_M61 ;
    wire SubBytesIns_Inst_Sbox_8_M60 ;
    wire SubBytesIns_Inst_Sbox_8_M59 ;
    wire SubBytesIns_Inst_Sbox_8_M58 ;
    wire SubBytesIns_Inst_Sbox_8_M57 ;
    wire SubBytesIns_Inst_Sbox_8_M56 ;
    wire SubBytesIns_Inst_Sbox_8_M55 ;
    wire SubBytesIns_Inst_Sbox_8_M54 ;
    wire SubBytesIns_Inst_Sbox_8_M53 ;
    wire SubBytesIns_Inst_Sbox_8_M52 ;
    wire SubBytesIns_Inst_Sbox_8_M51 ;
    wire SubBytesIns_Inst_Sbox_8_M50 ;
    wire SubBytesIns_Inst_Sbox_8_M49 ;
    wire SubBytesIns_Inst_Sbox_8_M48 ;
    wire SubBytesIns_Inst_Sbox_8_M47 ;
    wire SubBytesIns_Inst_Sbox_8_M46 ;
    wire SubBytesIns_Inst_Sbox_8_M45 ;
    wire SubBytesIns_Inst_Sbox_8_M44 ;
    wire SubBytesIns_Inst_Sbox_8_M43 ;
    wire SubBytesIns_Inst_Sbox_8_M42 ;
    wire SubBytesIns_Inst_Sbox_8_M41 ;
    wire SubBytesIns_Inst_Sbox_8_M40 ;
    wire SubBytesIns_Inst_Sbox_8_M39 ;
    wire SubBytesIns_Inst_Sbox_8_M38 ;
    wire SubBytesIns_Inst_Sbox_8_M37 ;
    wire SubBytesIns_Inst_Sbox_8_M36 ;
    wire SubBytesIns_Inst_Sbox_8_M35 ;
    wire SubBytesIns_Inst_Sbox_8_M34 ;
    wire SubBytesIns_Inst_Sbox_8_M33 ;
    wire SubBytesIns_Inst_Sbox_8_M32 ;
    wire SubBytesIns_Inst_Sbox_8_M31 ;
    wire SubBytesIns_Inst_Sbox_8_M30 ;
    wire SubBytesIns_Inst_Sbox_8_M29 ;
    wire SubBytesIns_Inst_Sbox_8_M28 ;
    wire SubBytesIns_Inst_Sbox_8_M27 ;
    wire SubBytesIns_Inst_Sbox_8_M26 ;
    wire SubBytesIns_Inst_Sbox_8_M25 ;
    wire SubBytesIns_Inst_Sbox_8_M24 ;
    wire SubBytesIns_Inst_Sbox_8_M23 ;
    wire SubBytesIns_Inst_Sbox_8_M22 ;
    wire SubBytesIns_Inst_Sbox_8_M21 ;
    wire SubBytesIns_Inst_Sbox_8_M20 ;
    wire SubBytesIns_Inst_Sbox_8_M19 ;
    wire SubBytesIns_Inst_Sbox_8_M18 ;
    wire SubBytesIns_Inst_Sbox_8_M17 ;
    wire SubBytesIns_Inst_Sbox_8_M16 ;
    wire SubBytesIns_Inst_Sbox_8_M15 ;
    wire SubBytesIns_Inst_Sbox_8_M14 ;
    wire SubBytesIns_Inst_Sbox_8_M13 ;
    wire SubBytesIns_Inst_Sbox_8_M12 ;
    wire SubBytesIns_Inst_Sbox_8_M11 ;
    wire SubBytesIns_Inst_Sbox_8_M10 ;
    wire SubBytesIns_Inst_Sbox_8_M9 ;
    wire SubBytesIns_Inst_Sbox_8_M8 ;
    wire SubBytesIns_Inst_Sbox_8_M7 ;
    wire SubBytesIns_Inst_Sbox_8_M6 ;
    wire SubBytesIns_Inst_Sbox_8_M5 ;
    wire SubBytesIns_Inst_Sbox_8_M4 ;
    wire SubBytesIns_Inst_Sbox_8_M3 ;
    wire SubBytesIns_Inst_Sbox_8_M2 ;
    wire SubBytesIns_Inst_Sbox_8_M1 ;
    wire SubBytesIns_Inst_Sbox_8_T27 ;
    wire SubBytesIns_Inst_Sbox_8_T26 ;
    wire SubBytesIns_Inst_Sbox_8_T25 ;
    wire SubBytesIns_Inst_Sbox_8_T24 ;
    wire SubBytesIns_Inst_Sbox_8_T23 ;
    wire SubBytesIns_Inst_Sbox_8_T22 ;
    wire SubBytesIns_Inst_Sbox_8_T21 ;
    wire SubBytesIns_Inst_Sbox_8_T20 ;
    wire SubBytesIns_Inst_Sbox_8_T19 ;
    wire SubBytesIns_Inst_Sbox_8_T18 ;
    wire SubBytesIns_Inst_Sbox_8_T17 ;
    wire SubBytesIns_Inst_Sbox_8_T16 ;
    wire SubBytesIns_Inst_Sbox_8_T15 ;
    wire SubBytesIns_Inst_Sbox_8_T14 ;
    wire SubBytesIns_Inst_Sbox_8_T13 ;
    wire SubBytesIns_Inst_Sbox_8_T12 ;
    wire SubBytesIns_Inst_Sbox_8_T11 ;
    wire SubBytesIns_Inst_Sbox_8_T10 ;
    wire SubBytesIns_Inst_Sbox_8_T9 ;
    wire SubBytesIns_Inst_Sbox_8_T8 ;
    wire SubBytesIns_Inst_Sbox_8_T7 ;
    wire SubBytesIns_Inst_Sbox_8_T6 ;
    wire SubBytesIns_Inst_Sbox_8_T5 ;
    wire SubBytesIns_Inst_Sbox_8_T4 ;
    wire SubBytesIns_Inst_Sbox_8_T3 ;
    wire SubBytesIns_Inst_Sbox_8_T2 ;
    wire SubBytesIns_Inst_Sbox_8_T1 ;
    wire SubBytesIns_Inst_Sbox_9_L29 ;
    wire SubBytesIns_Inst_Sbox_9_L28 ;
    wire SubBytesIns_Inst_Sbox_9_L27 ;
    wire SubBytesIns_Inst_Sbox_9_L26 ;
    wire SubBytesIns_Inst_Sbox_9_L25 ;
    wire SubBytesIns_Inst_Sbox_9_L24 ;
    wire SubBytesIns_Inst_Sbox_9_L23 ;
    wire SubBytesIns_Inst_Sbox_9_L22 ;
    wire SubBytesIns_Inst_Sbox_9_L21 ;
    wire SubBytesIns_Inst_Sbox_9_L20 ;
    wire SubBytesIns_Inst_Sbox_9_L19 ;
    wire SubBytesIns_Inst_Sbox_9_L18 ;
    wire SubBytesIns_Inst_Sbox_9_L17 ;
    wire SubBytesIns_Inst_Sbox_9_L16 ;
    wire SubBytesIns_Inst_Sbox_9_L15 ;
    wire SubBytesIns_Inst_Sbox_9_L14 ;
    wire SubBytesIns_Inst_Sbox_9_L13 ;
    wire SubBytesIns_Inst_Sbox_9_L12 ;
    wire SubBytesIns_Inst_Sbox_9_L11 ;
    wire SubBytesIns_Inst_Sbox_9_L10 ;
    wire SubBytesIns_Inst_Sbox_9_L9 ;
    wire SubBytesIns_Inst_Sbox_9_L8 ;
    wire SubBytesIns_Inst_Sbox_9_L7 ;
    wire SubBytesIns_Inst_Sbox_9_L6 ;
    wire SubBytesIns_Inst_Sbox_9_L5 ;
    wire SubBytesIns_Inst_Sbox_9_L4 ;
    wire SubBytesIns_Inst_Sbox_9_L3 ;
    wire SubBytesIns_Inst_Sbox_9_L2 ;
    wire SubBytesIns_Inst_Sbox_9_L1 ;
    wire SubBytesIns_Inst_Sbox_9_L0 ;
    wire SubBytesIns_Inst_Sbox_9_M63 ;
    wire SubBytesIns_Inst_Sbox_9_M62 ;
    wire SubBytesIns_Inst_Sbox_9_M61 ;
    wire SubBytesIns_Inst_Sbox_9_M60 ;
    wire SubBytesIns_Inst_Sbox_9_M59 ;
    wire SubBytesIns_Inst_Sbox_9_M58 ;
    wire SubBytesIns_Inst_Sbox_9_M57 ;
    wire SubBytesIns_Inst_Sbox_9_M56 ;
    wire SubBytesIns_Inst_Sbox_9_M55 ;
    wire SubBytesIns_Inst_Sbox_9_M54 ;
    wire SubBytesIns_Inst_Sbox_9_M53 ;
    wire SubBytesIns_Inst_Sbox_9_M52 ;
    wire SubBytesIns_Inst_Sbox_9_M51 ;
    wire SubBytesIns_Inst_Sbox_9_M50 ;
    wire SubBytesIns_Inst_Sbox_9_M49 ;
    wire SubBytesIns_Inst_Sbox_9_M48 ;
    wire SubBytesIns_Inst_Sbox_9_M47 ;
    wire SubBytesIns_Inst_Sbox_9_M46 ;
    wire SubBytesIns_Inst_Sbox_9_M45 ;
    wire SubBytesIns_Inst_Sbox_9_M44 ;
    wire SubBytesIns_Inst_Sbox_9_M43 ;
    wire SubBytesIns_Inst_Sbox_9_M42 ;
    wire SubBytesIns_Inst_Sbox_9_M41 ;
    wire SubBytesIns_Inst_Sbox_9_M40 ;
    wire SubBytesIns_Inst_Sbox_9_M39 ;
    wire SubBytesIns_Inst_Sbox_9_M38 ;
    wire SubBytesIns_Inst_Sbox_9_M37 ;
    wire SubBytesIns_Inst_Sbox_9_M36 ;
    wire SubBytesIns_Inst_Sbox_9_M35 ;
    wire SubBytesIns_Inst_Sbox_9_M34 ;
    wire SubBytesIns_Inst_Sbox_9_M33 ;
    wire SubBytesIns_Inst_Sbox_9_M32 ;
    wire SubBytesIns_Inst_Sbox_9_M31 ;
    wire SubBytesIns_Inst_Sbox_9_M30 ;
    wire SubBytesIns_Inst_Sbox_9_M29 ;
    wire SubBytesIns_Inst_Sbox_9_M28 ;
    wire SubBytesIns_Inst_Sbox_9_M27 ;
    wire SubBytesIns_Inst_Sbox_9_M26 ;
    wire SubBytesIns_Inst_Sbox_9_M25 ;
    wire SubBytesIns_Inst_Sbox_9_M24 ;
    wire SubBytesIns_Inst_Sbox_9_M23 ;
    wire SubBytesIns_Inst_Sbox_9_M22 ;
    wire SubBytesIns_Inst_Sbox_9_M21 ;
    wire SubBytesIns_Inst_Sbox_9_M20 ;
    wire SubBytesIns_Inst_Sbox_9_M19 ;
    wire SubBytesIns_Inst_Sbox_9_M18 ;
    wire SubBytesIns_Inst_Sbox_9_M17 ;
    wire SubBytesIns_Inst_Sbox_9_M16 ;
    wire SubBytesIns_Inst_Sbox_9_M15 ;
    wire SubBytesIns_Inst_Sbox_9_M14 ;
    wire SubBytesIns_Inst_Sbox_9_M13 ;
    wire SubBytesIns_Inst_Sbox_9_M12 ;
    wire SubBytesIns_Inst_Sbox_9_M11 ;
    wire SubBytesIns_Inst_Sbox_9_M10 ;
    wire SubBytesIns_Inst_Sbox_9_M9 ;
    wire SubBytesIns_Inst_Sbox_9_M8 ;
    wire SubBytesIns_Inst_Sbox_9_M7 ;
    wire SubBytesIns_Inst_Sbox_9_M6 ;
    wire SubBytesIns_Inst_Sbox_9_M5 ;
    wire SubBytesIns_Inst_Sbox_9_M4 ;
    wire SubBytesIns_Inst_Sbox_9_M3 ;
    wire SubBytesIns_Inst_Sbox_9_M2 ;
    wire SubBytesIns_Inst_Sbox_9_M1 ;
    wire SubBytesIns_Inst_Sbox_9_T27 ;
    wire SubBytesIns_Inst_Sbox_9_T26 ;
    wire SubBytesIns_Inst_Sbox_9_T25 ;
    wire SubBytesIns_Inst_Sbox_9_T24 ;
    wire SubBytesIns_Inst_Sbox_9_T23 ;
    wire SubBytesIns_Inst_Sbox_9_T22 ;
    wire SubBytesIns_Inst_Sbox_9_T21 ;
    wire SubBytesIns_Inst_Sbox_9_T20 ;
    wire SubBytesIns_Inst_Sbox_9_T19 ;
    wire SubBytesIns_Inst_Sbox_9_T18 ;
    wire SubBytesIns_Inst_Sbox_9_T17 ;
    wire SubBytesIns_Inst_Sbox_9_T16 ;
    wire SubBytesIns_Inst_Sbox_9_T15 ;
    wire SubBytesIns_Inst_Sbox_9_T14 ;
    wire SubBytesIns_Inst_Sbox_9_T13 ;
    wire SubBytesIns_Inst_Sbox_9_T12 ;
    wire SubBytesIns_Inst_Sbox_9_T11 ;
    wire SubBytesIns_Inst_Sbox_9_T10 ;
    wire SubBytesIns_Inst_Sbox_9_T9 ;
    wire SubBytesIns_Inst_Sbox_9_T8 ;
    wire SubBytesIns_Inst_Sbox_9_T7 ;
    wire SubBytesIns_Inst_Sbox_9_T6 ;
    wire SubBytesIns_Inst_Sbox_9_T5 ;
    wire SubBytesIns_Inst_Sbox_9_T4 ;
    wire SubBytesIns_Inst_Sbox_9_T3 ;
    wire SubBytesIns_Inst_Sbox_9_T2 ;
    wire SubBytesIns_Inst_Sbox_9_T1 ;
    wire SubBytesIns_Inst_Sbox_10_L29 ;
    wire SubBytesIns_Inst_Sbox_10_L28 ;
    wire SubBytesIns_Inst_Sbox_10_L27 ;
    wire SubBytesIns_Inst_Sbox_10_L26 ;
    wire SubBytesIns_Inst_Sbox_10_L25 ;
    wire SubBytesIns_Inst_Sbox_10_L24 ;
    wire SubBytesIns_Inst_Sbox_10_L23 ;
    wire SubBytesIns_Inst_Sbox_10_L22 ;
    wire SubBytesIns_Inst_Sbox_10_L21 ;
    wire SubBytesIns_Inst_Sbox_10_L20 ;
    wire SubBytesIns_Inst_Sbox_10_L19 ;
    wire SubBytesIns_Inst_Sbox_10_L18 ;
    wire SubBytesIns_Inst_Sbox_10_L17 ;
    wire SubBytesIns_Inst_Sbox_10_L16 ;
    wire SubBytesIns_Inst_Sbox_10_L15 ;
    wire SubBytesIns_Inst_Sbox_10_L14 ;
    wire SubBytesIns_Inst_Sbox_10_L13 ;
    wire SubBytesIns_Inst_Sbox_10_L12 ;
    wire SubBytesIns_Inst_Sbox_10_L11 ;
    wire SubBytesIns_Inst_Sbox_10_L10 ;
    wire SubBytesIns_Inst_Sbox_10_L9 ;
    wire SubBytesIns_Inst_Sbox_10_L8 ;
    wire SubBytesIns_Inst_Sbox_10_L7 ;
    wire SubBytesIns_Inst_Sbox_10_L6 ;
    wire SubBytesIns_Inst_Sbox_10_L5 ;
    wire SubBytesIns_Inst_Sbox_10_L4 ;
    wire SubBytesIns_Inst_Sbox_10_L3 ;
    wire SubBytesIns_Inst_Sbox_10_L2 ;
    wire SubBytesIns_Inst_Sbox_10_L1 ;
    wire SubBytesIns_Inst_Sbox_10_L0 ;
    wire SubBytesIns_Inst_Sbox_10_M63 ;
    wire SubBytesIns_Inst_Sbox_10_M62 ;
    wire SubBytesIns_Inst_Sbox_10_M61 ;
    wire SubBytesIns_Inst_Sbox_10_M60 ;
    wire SubBytesIns_Inst_Sbox_10_M59 ;
    wire SubBytesIns_Inst_Sbox_10_M58 ;
    wire SubBytesIns_Inst_Sbox_10_M57 ;
    wire SubBytesIns_Inst_Sbox_10_M56 ;
    wire SubBytesIns_Inst_Sbox_10_M55 ;
    wire SubBytesIns_Inst_Sbox_10_M54 ;
    wire SubBytesIns_Inst_Sbox_10_M53 ;
    wire SubBytesIns_Inst_Sbox_10_M52 ;
    wire SubBytesIns_Inst_Sbox_10_M51 ;
    wire SubBytesIns_Inst_Sbox_10_M50 ;
    wire SubBytesIns_Inst_Sbox_10_M49 ;
    wire SubBytesIns_Inst_Sbox_10_M48 ;
    wire SubBytesIns_Inst_Sbox_10_M47 ;
    wire SubBytesIns_Inst_Sbox_10_M46 ;
    wire SubBytesIns_Inst_Sbox_10_M45 ;
    wire SubBytesIns_Inst_Sbox_10_M44 ;
    wire SubBytesIns_Inst_Sbox_10_M43 ;
    wire SubBytesIns_Inst_Sbox_10_M42 ;
    wire SubBytesIns_Inst_Sbox_10_M41 ;
    wire SubBytesIns_Inst_Sbox_10_M40 ;
    wire SubBytesIns_Inst_Sbox_10_M39 ;
    wire SubBytesIns_Inst_Sbox_10_M38 ;
    wire SubBytesIns_Inst_Sbox_10_M37 ;
    wire SubBytesIns_Inst_Sbox_10_M36 ;
    wire SubBytesIns_Inst_Sbox_10_M35 ;
    wire SubBytesIns_Inst_Sbox_10_M34 ;
    wire SubBytesIns_Inst_Sbox_10_M33 ;
    wire SubBytesIns_Inst_Sbox_10_M32 ;
    wire SubBytesIns_Inst_Sbox_10_M31 ;
    wire SubBytesIns_Inst_Sbox_10_M30 ;
    wire SubBytesIns_Inst_Sbox_10_M29 ;
    wire SubBytesIns_Inst_Sbox_10_M28 ;
    wire SubBytesIns_Inst_Sbox_10_M27 ;
    wire SubBytesIns_Inst_Sbox_10_M26 ;
    wire SubBytesIns_Inst_Sbox_10_M25 ;
    wire SubBytesIns_Inst_Sbox_10_M24 ;
    wire SubBytesIns_Inst_Sbox_10_M23 ;
    wire SubBytesIns_Inst_Sbox_10_M22 ;
    wire SubBytesIns_Inst_Sbox_10_M21 ;
    wire SubBytesIns_Inst_Sbox_10_M20 ;
    wire SubBytesIns_Inst_Sbox_10_M19 ;
    wire SubBytesIns_Inst_Sbox_10_M18 ;
    wire SubBytesIns_Inst_Sbox_10_M17 ;
    wire SubBytesIns_Inst_Sbox_10_M16 ;
    wire SubBytesIns_Inst_Sbox_10_M15 ;
    wire SubBytesIns_Inst_Sbox_10_M14 ;
    wire SubBytesIns_Inst_Sbox_10_M13 ;
    wire SubBytesIns_Inst_Sbox_10_M12 ;
    wire SubBytesIns_Inst_Sbox_10_M11 ;
    wire SubBytesIns_Inst_Sbox_10_M10 ;
    wire SubBytesIns_Inst_Sbox_10_M9 ;
    wire SubBytesIns_Inst_Sbox_10_M8 ;
    wire SubBytesIns_Inst_Sbox_10_M7 ;
    wire SubBytesIns_Inst_Sbox_10_M6 ;
    wire SubBytesIns_Inst_Sbox_10_M5 ;
    wire SubBytesIns_Inst_Sbox_10_M4 ;
    wire SubBytesIns_Inst_Sbox_10_M3 ;
    wire SubBytesIns_Inst_Sbox_10_M2 ;
    wire SubBytesIns_Inst_Sbox_10_M1 ;
    wire SubBytesIns_Inst_Sbox_10_T27 ;
    wire SubBytesIns_Inst_Sbox_10_T26 ;
    wire SubBytesIns_Inst_Sbox_10_T25 ;
    wire SubBytesIns_Inst_Sbox_10_T24 ;
    wire SubBytesIns_Inst_Sbox_10_T23 ;
    wire SubBytesIns_Inst_Sbox_10_T22 ;
    wire SubBytesIns_Inst_Sbox_10_T21 ;
    wire SubBytesIns_Inst_Sbox_10_T20 ;
    wire SubBytesIns_Inst_Sbox_10_T19 ;
    wire SubBytesIns_Inst_Sbox_10_T18 ;
    wire SubBytesIns_Inst_Sbox_10_T17 ;
    wire SubBytesIns_Inst_Sbox_10_T16 ;
    wire SubBytesIns_Inst_Sbox_10_T15 ;
    wire SubBytesIns_Inst_Sbox_10_T14 ;
    wire SubBytesIns_Inst_Sbox_10_T13 ;
    wire SubBytesIns_Inst_Sbox_10_T12 ;
    wire SubBytesIns_Inst_Sbox_10_T11 ;
    wire SubBytesIns_Inst_Sbox_10_T10 ;
    wire SubBytesIns_Inst_Sbox_10_T9 ;
    wire SubBytesIns_Inst_Sbox_10_T8 ;
    wire SubBytesIns_Inst_Sbox_10_T7 ;
    wire SubBytesIns_Inst_Sbox_10_T6 ;
    wire SubBytesIns_Inst_Sbox_10_T5 ;
    wire SubBytesIns_Inst_Sbox_10_T4 ;
    wire SubBytesIns_Inst_Sbox_10_T3 ;
    wire SubBytesIns_Inst_Sbox_10_T2 ;
    wire SubBytesIns_Inst_Sbox_10_T1 ;
    wire SubBytesIns_Inst_Sbox_11_L29 ;
    wire SubBytesIns_Inst_Sbox_11_L28 ;
    wire SubBytesIns_Inst_Sbox_11_L27 ;
    wire SubBytesIns_Inst_Sbox_11_L26 ;
    wire SubBytesIns_Inst_Sbox_11_L25 ;
    wire SubBytesIns_Inst_Sbox_11_L24 ;
    wire SubBytesIns_Inst_Sbox_11_L23 ;
    wire SubBytesIns_Inst_Sbox_11_L22 ;
    wire SubBytesIns_Inst_Sbox_11_L21 ;
    wire SubBytesIns_Inst_Sbox_11_L20 ;
    wire SubBytesIns_Inst_Sbox_11_L19 ;
    wire SubBytesIns_Inst_Sbox_11_L18 ;
    wire SubBytesIns_Inst_Sbox_11_L17 ;
    wire SubBytesIns_Inst_Sbox_11_L16 ;
    wire SubBytesIns_Inst_Sbox_11_L15 ;
    wire SubBytesIns_Inst_Sbox_11_L14 ;
    wire SubBytesIns_Inst_Sbox_11_L13 ;
    wire SubBytesIns_Inst_Sbox_11_L12 ;
    wire SubBytesIns_Inst_Sbox_11_L11 ;
    wire SubBytesIns_Inst_Sbox_11_L10 ;
    wire SubBytesIns_Inst_Sbox_11_L9 ;
    wire SubBytesIns_Inst_Sbox_11_L8 ;
    wire SubBytesIns_Inst_Sbox_11_L7 ;
    wire SubBytesIns_Inst_Sbox_11_L6 ;
    wire SubBytesIns_Inst_Sbox_11_L5 ;
    wire SubBytesIns_Inst_Sbox_11_L4 ;
    wire SubBytesIns_Inst_Sbox_11_L3 ;
    wire SubBytesIns_Inst_Sbox_11_L2 ;
    wire SubBytesIns_Inst_Sbox_11_L1 ;
    wire SubBytesIns_Inst_Sbox_11_L0 ;
    wire SubBytesIns_Inst_Sbox_11_M63 ;
    wire SubBytesIns_Inst_Sbox_11_M62 ;
    wire SubBytesIns_Inst_Sbox_11_M61 ;
    wire SubBytesIns_Inst_Sbox_11_M60 ;
    wire SubBytesIns_Inst_Sbox_11_M59 ;
    wire SubBytesIns_Inst_Sbox_11_M58 ;
    wire SubBytesIns_Inst_Sbox_11_M57 ;
    wire SubBytesIns_Inst_Sbox_11_M56 ;
    wire SubBytesIns_Inst_Sbox_11_M55 ;
    wire SubBytesIns_Inst_Sbox_11_M54 ;
    wire SubBytesIns_Inst_Sbox_11_M53 ;
    wire SubBytesIns_Inst_Sbox_11_M52 ;
    wire SubBytesIns_Inst_Sbox_11_M51 ;
    wire SubBytesIns_Inst_Sbox_11_M50 ;
    wire SubBytesIns_Inst_Sbox_11_M49 ;
    wire SubBytesIns_Inst_Sbox_11_M48 ;
    wire SubBytesIns_Inst_Sbox_11_M47 ;
    wire SubBytesIns_Inst_Sbox_11_M46 ;
    wire SubBytesIns_Inst_Sbox_11_M45 ;
    wire SubBytesIns_Inst_Sbox_11_M44 ;
    wire SubBytesIns_Inst_Sbox_11_M43 ;
    wire SubBytesIns_Inst_Sbox_11_M42 ;
    wire SubBytesIns_Inst_Sbox_11_M41 ;
    wire SubBytesIns_Inst_Sbox_11_M40 ;
    wire SubBytesIns_Inst_Sbox_11_M39 ;
    wire SubBytesIns_Inst_Sbox_11_M38 ;
    wire SubBytesIns_Inst_Sbox_11_M37 ;
    wire SubBytesIns_Inst_Sbox_11_M36 ;
    wire SubBytesIns_Inst_Sbox_11_M35 ;
    wire SubBytesIns_Inst_Sbox_11_M34 ;
    wire SubBytesIns_Inst_Sbox_11_M33 ;
    wire SubBytesIns_Inst_Sbox_11_M32 ;
    wire SubBytesIns_Inst_Sbox_11_M31 ;
    wire SubBytesIns_Inst_Sbox_11_M30 ;
    wire SubBytesIns_Inst_Sbox_11_M29 ;
    wire SubBytesIns_Inst_Sbox_11_M28 ;
    wire SubBytesIns_Inst_Sbox_11_M27 ;
    wire SubBytesIns_Inst_Sbox_11_M26 ;
    wire SubBytesIns_Inst_Sbox_11_M25 ;
    wire SubBytesIns_Inst_Sbox_11_M24 ;
    wire SubBytesIns_Inst_Sbox_11_M23 ;
    wire SubBytesIns_Inst_Sbox_11_M22 ;
    wire SubBytesIns_Inst_Sbox_11_M21 ;
    wire SubBytesIns_Inst_Sbox_11_M20 ;
    wire SubBytesIns_Inst_Sbox_11_M19 ;
    wire SubBytesIns_Inst_Sbox_11_M18 ;
    wire SubBytesIns_Inst_Sbox_11_M17 ;
    wire SubBytesIns_Inst_Sbox_11_M16 ;
    wire SubBytesIns_Inst_Sbox_11_M15 ;
    wire SubBytesIns_Inst_Sbox_11_M14 ;
    wire SubBytesIns_Inst_Sbox_11_M13 ;
    wire SubBytesIns_Inst_Sbox_11_M12 ;
    wire SubBytesIns_Inst_Sbox_11_M11 ;
    wire SubBytesIns_Inst_Sbox_11_M10 ;
    wire SubBytesIns_Inst_Sbox_11_M9 ;
    wire SubBytesIns_Inst_Sbox_11_M8 ;
    wire SubBytesIns_Inst_Sbox_11_M7 ;
    wire SubBytesIns_Inst_Sbox_11_M6 ;
    wire SubBytesIns_Inst_Sbox_11_M5 ;
    wire SubBytesIns_Inst_Sbox_11_M4 ;
    wire SubBytesIns_Inst_Sbox_11_M3 ;
    wire SubBytesIns_Inst_Sbox_11_M2 ;
    wire SubBytesIns_Inst_Sbox_11_M1 ;
    wire SubBytesIns_Inst_Sbox_11_T27 ;
    wire SubBytesIns_Inst_Sbox_11_T26 ;
    wire SubBytesIns_Inst_Sbox_11_T25 ;
    wire SubBytesIns_Inst_Sbox_11_T24 ;
    wire SubBytesIns_Inst_Sbox_11_T23 ;
    wire SubBytesIns_Inst_Sbox_11_T22 ;
    wire SubBytesIns_Inst_Sbox_11_T21 ;
    wire SubBytesIns_Inst_Sbox_11_T20 ;
    wire SubBytesIns_Inst_Sbox_11_T19 ;
    wire SubBytesIns_Inst_Sbox_11_T18 ;
    wire SubBytesIns_Inst_Sbox_11_T17 ;
    wire SubBytesIns_Inst_Sbox_11_T16 ;
    wire SubBytesIns_Inst_Sbox_11_T15 ;
    wire SubBytesIns_Inst_Sbox_11_T14 ;
    wire SubBytesIns_Inst_Sbox_11_T13 ;
    wire SubBytesIns_Inst_Sbox_11_T12 ;
    wire SubBytesIns_Inst_Sbox_11_T11 ;
    wire SubBytesIns_Inst_Sbox_11_T10 ;
    wire SubBytesIns_Inst_Sbox_11_T9 ;
    wire SubBytesIns_Inst_Sbox_11_T8 ;
    wire SubBytesIns_Inst_Sbox_11_T7 ;
    wire SubBytesIns_Inst_Sbox_11_T6 ;
    wire SubBytesIns_Inst_Sbox_11_T5 ;
    wire SubBytesIns_Inst_Sbox_11_T4 ;
    wire SubBytesIns_Inst_Sbox_11_T3 ;
    wire SubBytesIns_Inst_Sbox_11_T2 ;
    wire SubBytesIns_Inst_Sbox_11_T1 ;
    wire SubBytesIns_Inst_Sbox_12_L29 ;
    wire SubBytesIns_Inst_Sbox_12_L28 ;
    wire SubBytesIns_Inst_Sbox_12_L27 ;
    wire SubBytesIns_Inst_Sbox_12_L26 ;
    wire SubBytesIns_Inst_Sbox_12_L25 ;
    wire SubBytesIns_Inst_Sbox_12_L24 ;
    wire SubBytesIns_Inst_Sbox_12_L23 ;
    wire SubBytesIns_Inst_Sbox_12_L22 ;
    wire SubBytesIns_Inst_Sbox_12_L21 ;
    wire SubBytesIns_Inst_Sbox_12_L20 ;
    wire SubBytesIns_Inst_Sbox_12_L19 ;
    wire SubBytesIns_Inst_Sbox_12_L18 ;
    wire SubBytesIns_Inst_Sbox_12_L17 ;
    wire SubBytesIns_Inst_Sbox_12_L16 ;
    wire SubBytesIns_Inst_Sbox_12_L15 ;
    wire SubBytesIns_Inst_Sbox_12_L14 ;
    wire SubBytesIns_Inst_Sbox_12_L13 ;
    wire SubBytesIns_Inst_Sbox_12_L12 ;
    wire SubBytesIns_Inst_Sbox_12_L11 ;
    wire SubBytesIns_Inst_Sbox_12_L10 ;
    wire SubBytesIns_Inst_Sbox_12_L9 ;
    wire SubBytesIns_Inst_Sbox_12_L8 ;
    wire SubBytesIns_Inst_Sbox_12_L7 ;
    wire SubBytesIns_Inst_Sbox_12_L6 ;
    wire SubBytesIns_Inst_Sbox_12_L5 ;
    wire SubBytesIns_Inst_Sbox_12_L4 ;
    wire SubBytesIns_Inst_Sbox_12_L3 ;
    wire SubBytesIns_Inst_Sbox_12_L2 ;
    wire SubBytesIns_Inst_Sbox_12_L1 ;
    wire SubBytesIns_Inst_Sbox_12_L0 ;
    wire SubBytesIns_Inst_Sbox_12_M63 ;
    wire SubBytesIns_Inst_Sbox_12_M62 ;
    wire SubBytesIns_Inst_Sbox_12_M61 ;
    wire SubBytesIns_Inst_Sbox_12_M60 ;
    wire SubBytesIns_Inst_Sbox_12_M59 ;
    wire SubBytesIns_Inst_Sbox_12_M58 ;
    wire SubBytesIns_Inst_Sbox_12_M57 ;
    wire SubBytesIns_Inst_Sbox_12_M56 ;
    wire SubBytesIns_Inst_Sbox_12_M55 ;
    wire SubBytesIns_Inst_Sbox_12_M54 ;
    wire SubBytesIns_Inst_Sbox_12_M53 ;
    wire SubBytesIns_Inst_Sbox_12_M52 ;
    wire SubBytesIns_Inst_Sbox_12_M51 ;
    wire SubBytesIns_Inst_Sbox_12_M50 ;
    wire SubBytesIns_Inst_Sbox_12_M49 ;
    wire SubBytesIns_Inst_Sbox_12_M48 ;
    wire SubBytesIns_Inst_Sbox_12_M47 ;
    wire SubBytesIns_Inst_Sbox_12_M46 ;
    wire SubBytesIns_Inst_Sbox_12_M45 ;
    wire SubBytesIns_Inst_Sbox_12_M44 ;
    wire SubBytesIns_Inst_Sbox_12_M43 ;
    wire SubBytesIns_Inst_Sbox_12_M42 ;
    wire SubBytesIns_Inst_Sbox_12_M41 ;
    wire SubBytesIns_Inst_Sbox_12_M40 ;
    wire SubBytesIns_Inst_Sbox_12_M39 ;
    wire SubBytesIns_Inst_Sbox_12_M38 ;
    wire SubBytesIns_Inst_Sbox_12_M37 ;
    wire SubBytesIns_Inst_Sbox_12_M36 ;
    wire SubBytesIns_Inst_Sbox_12_M35 ;
    wire SubBytesIns_Inst_Sbox_12_M34 ;
    wire SubBytesIns_Inst_Sbox_12_M33 ;
    wire SubBytesIns_Inst_Sbox_12_M32 ;
    wire SubBytesIns_Inst_Sbox_12_M31 ;
    wire SubBytesIns_Inst_Sbox_12_M30 ;
    wire SubBytesIns_Inst_Sbox_12_M29 ;
    wire SubBytesIns_Inst_Sbox_12_M28 ;
    wire SubBytesIns_Inst_Sbox_12_M27 ;
    wire SubBytesIns_Inst_Sbox_12_M26 ;
    wire SubBytesIns_Inst_Sbox_12_M25 ;
    wire SubBytesIns_Inst_Sbox_12_M24 ;
    wire SubBytesIns_Inst_Sbox_12_M23 ;
    wire SubBytesIns_Inst_Sbox_12_M22 ;
    wire SubBytesIns_Inst_Sbox_12_M21 ;
    wire SubBytesIns_Inst_Sbox_12_M20 ;
    wire SubBytesIns_Inst_Sbox_12_M19 ;
    wire SubBytesIns_Inst_Sbox_12_M18 ;
    wire SubBytesIns_Inst_Sbox_12_M17 ;
    wire SubBytesIns_Inst_Sbox_12_M16 ;
    wire SubBytesIns_Inst_Sbox_12_M15 ;
    wire SubBytesIns_Inst_Sbox_12_M14 ;
    wire SubBytesIns_Inst_Sbox_12_M13 ;
    wire SubBytesIns_Inst_Sbox_12_M12 ;
    wire SubBytesIns_Inst_Sbox_12_M11 ;
    wire SubBytesIns_Inst_Sbox_12_M10 ;
    wire SubBytesIns_Inst_Sbox_12_M9 ;
    wire SubBytesIns_Inst_Sbox_12_M8 ;
    wire SubBytesIns_Inst_Sbox_12_M7 ;
    wire SubBytesIns_Inst_Sbox_12_M6 ;
    wire SubBytesIns_Inst_Sbox_12_M5 ;
    wire SubBytesIns_Inst_Sbox_12_M4 ;
    wire SubBytesIns_Inst_Sbox_12_M3 ;
    wire SubBytesIns_Inst_Sbox_12_M2 ;
    wire SubBytesIns_Inst_Sbox_12_M1 ;
    wire SubBytesIns_Inst_Sbox_12_T27 ;
    wire SubBytesIns_Inst_Sbox_12_T26 ;
    wire SubBytesIns_Inst_Sbox_12_T25 ;
    wire SubBytesIns_Inst_Sbox_12_T24 ;
    wire SubBytesIns_Inst_Sbox_12_T23 ;
    wire SubBytesIns_Inst_Sbox_12_T22 ;
    wire SubBytesIns_Inst_Sbox_12_T21 ;
    wire SubBytesIns_Inst_Sbox_12_T20 ;
    wire SubBytesIns_Inst_Sbox_12_T19 ;
    wire SubBytesIns_Inst_Sbox_12_T18 ;
    wire SubBytesIns_Inst_Sbox_12_T17 ;
    wire SubBytesIns_Inst_Sbox_12_T16 ;
    wire SubBytesIns_Inst_Sbox_12_T15 ;
    wire SubBytesIns_Inst_Sbox_12_T14 ;
    wire SubBytesIns_Inst_Sbox_12_T13 ;
    wire SubBytesIns_Inst_Sbox_12_T12 ;
    wire SubBytesIns_Inst_Sbox_12_T11 ;
    wire SubBytesIns_Inst_Sbox_12_T10 ;
    wire SubBytesIns_Inst_Sbox_12_T9 ;
    wire SubBytesIns_Inst_Sbox_12_T8 ;
    wire SubBytesIns_Inst_Sbox_12_T7 ;
    wire SubBytesIns_Inst_Sbox_12_T6 ;
    wire SubBytesIns_Inst_Sbox_12_T5 ;
    wire SubBytesIns_Inst_Sbox_12_T4 ;
    wire SubBytesIns_Inst_Sbox_12_T3 ;
    wire SubBytesIns_Inst_Sbox_12_T2 ;
    wire SubBytesIns_Inst_Sbox_12_T1 ;
    wire SubBytesIns_Inst_Sbox_13_L29 ;
    wire SubBytesIns_Inst_Sbox_13_L28 ;
    wire SubBytesIns_Inst_Sbox_13_L27 ;
    wire SubBytesIns_Inst_Sbox_13_L26 ;
    wire SubBytesIns_Inst_Sbox_13_L25 ;
    wire SubBytesIns_Inst_Sbox_13_L24 ;
    wire SubBytesIns_Inst_Sbox_13_L23 ;
    wire SubBytesIns_Inst_Sbox_13_L22 ;
    wire SubBytesIns_Inst_Sbox_13_L21 ;
    wire SubBytesIns_Inst_Sbox_13_L20 ;
    wire SubBytesIns_Inst_Sbox_13_L19 ;
    wire SubBytesIns_Inst_Sbox_13_L18 ;
    wire SubBytesIns_Inst_Sbox_13_L17 ;
    wire SubBytesIns_Inst_Sbox_13_L16 ;
    wire SubBytesIns_Inst_Sbox_13_L15 ;
    wire SubBytesIns_Inst_Sbox_13_L14 ;
    wire SubBytesIns_Inst_Sbox_13_L13 ;
    wire SubBytesIns_Inst_Sbox_13_L12 ;
    wire SubBytesIns_Inst_Sbox_13_L11 ;
    wire SubBytesIns_Inst_Sbox_13_L10 ;
    wire SubBytesIns_Inst_Sbox_13_L9 ;
    wire SubBytesIns_Inst_Sbox_13_L8 ;
    wire SubBytesIns_Inst_Sbox_13_L7 ;
    wire SubBytesIns_Inst_Sbox_13_L6 ;
    wire SubBytesIns_Inst_Sbox_13_L5 ;
    wire SubBytesIns_Inst_Sbox_13_L4 ;
    wire SubBytesIns_Inst_Sbox_13_L3 ;
    wire SubBytesIns_Inst_Sbox_13_L2 ;
    wire SubBytesIns_Inst_Sbox_13_L1 ;
    wire SubBytesIns_Inst_Sbox_13_L0 ;
    wire SubBytesIns_Inst_Sbox_13_M63 ;
    wire SubBytesIns_Inst_Sbox_13_M62 ;
    wire SubBytesIns_Inst_Sbox_13_M61 ;
    wire SubBytesIns_Inst_Sbox_13_M60 ;
    wire SubBytesIns_Inst_Sbox_13_M59 ;
    wire SubBytesIns_Inst_Sbox_13_M58 ;
    wire SubBytesIns_Inst_Sbox_13_M57 ;
    wire SubBytesIns_Inst_Sbox_13_M56 ;
    wire SubBytesIns_Inst_Sbox_13_M55 ;
    wire SubBytesIns_Inst_Sbox_13_M54 ;
    wire SubBytesIns_Inst_Sbox_13_M53 ;
    wire SubBytesIns_Inst_Sbox_13_M52 ;
    wire SubBytesIns_Inst_Sbox_13_M51 ;
    wire SubBytesIns_Inst_Sbox_13_M50 ;
    wire SubBytesIns_Inst_Sbox_13_M49 ;
    wire SubBytesIns_Inst_Sbox_13_M48 ;
    wire SubBytesIns_Inst_Sbox_13_M47 ;
    wire SubBytesIns_Inst_Sbox_13_M46 ;
    wire SubBytesIns_Inst_Sbox_13_M45 ;
    wire SubBytesIns_Inst_Sbox_13_M44 ;
    wire SubBytesIns_Inst_Sbox_13_M43 ;
    wire SubBytesIns_Inst_Sbox_13_M42 ;
    wire SubBytesIns_Inst_Sbox_13_M41 ;
    wire SubBytesIns_Inst_Sbox_13_M40 ;
    wire SubBytesIns_Inst_Sbox_13_M39 ;
    wire SubBytesIns_Inst_Sbox_13_M38 ;
    wire SubBytesIns_Inst_Sbox_13_M37 ;
    wire SubBytesIns_Inst_Sbox_13_M36 ;
    wire SubBytesIns_Inst_Sbox_13_M35 ;
    wire SubBytesIns_Inst_Sbox_13_M34 ;
    wire SubBytesIns_Inst_Sbox_13_M33 ;
    wire SubBytesIns_Inst_Sbox_13_M32 ;
    wire SubBytesIns_Inst_Sbox_13_M31 ;
    wire SubBytesIns_Inst_Sbox_13_M30 ;
    wire SubBytesIns_Inst_Sbox_13_M29 ;
    wire SubBytesIns_Inst_Sbox_13_M28 ;
    wire SubBytesIns_Inst_Sbox_13_M27 ;
    wire SubBytesIns_Inst_Sbox_13_M26 ;
    wire SubBytesIns_Inst_Sbox_13_M25 ;
    wire SubBytesIns_Inst_Sbox_13_M24 ;
    wire SubBytesIns_Inst_Sbox_13_M23 ;
    wire SubBytesIns_Inst_Sbox_13_M22 ;
    wire SubBytesIns_Inst_Sbox_13_M21 ;
    wire SubBytesIns_Inst_Sbox_13_M20 ;
    wire SubBytesIns_Inst_Sbox_13_M19 ;
    wire SubBytesIns_Inst_Sbox_13_M18 ;
    wire SubBytesIns_Inst_Sbox_13_M17 ;
    wire SubBytesIns_Inst_Sbox_13_M16 ;
    wire SubBytesIns_Inst_Sbox_13_M15 ;
    wire SubBytesIns_Inst_Sbox_13_M14 ;
    wire SubBytesIns_Inst_Sbox_13_M13 ;
    wire SubBytesIns_Inst_Sbox_13_M12 ;
    wire SubBytesIns_Inst_Sbox_13_M11 ;
    wire SubBytesIns_Inst_Sbox_13_M10 ;
    wire SubBytesIns_Inst_Sbox_13_M9 ;
    wire SubBytesIns_Inst_Sbox_13_M8 ;
    wire SubBytesIns_Inst_Sbox_13_M7 ;
    wire SubBytesIns_Inst_Sbox_13_M6 ;
    wire SubBytesIns_Inst_Sbox_13_M5 ;
    wire SubBytesIns_Inst_Sbox_13_M4 ;
    wire SubBytesIns_Inst_Sbox_13_M3 ;
    wire SubBytesIns_Inst_Sbox_13_M2 ;
    wire SubBytesIns_Inst_Sbox_13_M1 ;
    wire SubBytesIns_Inst_Sbox_13_T27 ;
    wire SubBytesIns_Inst_Sbox_13_T26 ;
    wire SubBytesIns_Inst_Sbox_13_T25 ;
    wire SubBytesIns_Inst_Sbox_13_T24 ;
    wire SubBytesIns_Inst_Sbox_13_T23 ;
    wire SubBytesIns_Inst_Sbox_13_T22 ;
    wire SubBytesIns_Inst_Sbox_13_T21 ;
    wire SubBytesIns_Inst_Sbox_13_T20 ;
    wire SubBytesIns_Inst_Sbox_13_T19 ;
    wire SubBytesIns_Inst_Sbox_13_T18 ;
    wire SubBytesIns_Inst_Sbox_13_T17 ;
    wire SubBytesIns_Inst_Sbox_13_T16 ;
    wire SubBytesIns_Inst_Sbox_13_T15 ;
    wire SubBytesIns_Inst_Sbox_13_T14 ;
    wire SubBytesIns_Inst_Sbox_13_T13 ;
    wire SubBytesIns_Inst_Sbox_13_T12 ;
    wire SubBytesIns_Inst_Sbox_13_T11 ;
    wire SubBytesIns_Inst_Sbox_13_T10 ;
    wire SubBytesIns_Inst_Sbox_13_T9 ;
    wire SubBytesIns_Inst_Sbox_13_T8 ;
    wire SubBytesIns_Inst_Sbox_13_T7 ;
    wire SubBytesIns_Inst_Sbox_13_T6 ;
    wire SubBytesIns_Inst_Sbox_13_T5 ;
    wire SubBytesIns_Inst_Sbox_13_T4 ;
    wire SubBytesIns_Inst_Sbox_13_T3 ;
    wire SubBytesIns_Inst_Sbox_13_T2 ;
    wire SubBytesIns_Inst_Sbox_13_T1 ;
    wire SubBytesIns_Inst_Sbox_14_L29 ;
    wire SubBytesIns_Inst_Sbox_14_L28 ;
    wire SubBytesIns_Inst_Sbox_14_L27 ;
    wire SubBytesIns_Inst_Sbox_14_L26 ;
    wire SubBytesIns_Inst_Sbox_14_L25 ;
    wire SubBytesIns_Inst_Sbox_14_L24 ;
    wire SubBytesIns_Inst_Sbox_14_L23 ;
    wire SubBytesIns_Inst_Sbox_14_L22 ;
    wire SubBytesIns_Inst_Sbox_14_L21 ;
    wire SubBytesIns_Inst_Sbox_14_L20 ;
    wire SubBytesIns_Inst_Sbox_14_L19 ;
    wire SubBytesIns_Inst_Sbox_14_L18 ;
    wire SubBytesIns_Inst_Sbox_14_L17 ;
    wire SubBytesIns_Inst_Sbox_14_L16 ;
    wire SubBytesIns_Inst_Sbox_14_L15 ;
    wire SubBytesIns_Inst_Sbox_14_L14 ;
    wire SubBytesIns_Inst_Sbox_14_L13 ;
    wire SubBytesIns_Inst_Sbox_14_L12 ;
    wire SubBytesIns_Inst_Sbox_14_L11 ;
    wire SubBytesIns_Inst_Sbox_14_L10 ;
    wire SubBytesIns_Inst_Sbox_14_L9 ;
    wire SubBytesIns_Inst_Sbox_14_L8 ;
    wire SubBytesIns_Inst_Sbox_14_L7 ;
    wire SubBytesIns_Inst_Sbox_14_L6 ;
    wire SubBytesIns_Inst_Sbox_14_L5 ;
    wire SubBytesIns_Inst_Sbox_14_L4 ;
    wire SubBytesIns_Inst_Sbox_14_L3 ;
    wire SubBytesIns_Inst_Sbox_14_L2 ;
    wire SubBytesIns_Inst_Sbox_14_L1 ;
    wire SubBytesIns_Inst_Sbox_14_L0 ;
    wire SubBytesIns_Inst_Sbox_14_M63 ;
    wire SubBytesIns_Inst_Sbox_14_M62 ;
    wire SubBytesIns_Inst_Sbox_14_M61 ;
    wire SubBytesIns_Inst_Sbox_14_M60 ;
    wire SubBytesIns_Inst_Sbox_14_M59 ;
    wire SubBytesIns_Inst_Sbox_14_M58 ;
    wire SubBytesIns_Inst_Sbox_14_M57 ;
    wire SubBytesIns_Inst_Sbox_14_M56 ;
    wire SubBytesIns_Inst_Sbox_14_M55 ;
    wire SubBytesIns_Inst_Sbox_14_M54 ;
    wire SubBytesIns_Inst_Sbox_14_M53 ;
    wire SubBytesIns_Inst_Sbox_14_M52 ;
    wire SubBytesIns_Inst_Sbox_14_M51 ;
    wire SubBytesIns_Inst_Sbox_14_M50 ;
    wire SubBytesIns_Inst_Sbox_14_M49 ;
    wire SubBytesIns_Inst_Sbox_14_M48 ;
    wire SubBytesIns_Inst_Sbox_14_M47 ;
    wire SubBytesIns_Inst_Sbox_14_M46 ;
    wire SubBytesIns_Inst_Sbox_14_M45 ;
    wire SubBytesIns_Inst_Sbox_14_M44 ;
    wire SubBytesIns_Inst_Sbox_14_M43 ;
    wire SubBytesIns_Inst_Sbox_14_M42 ;
    wire SubBytesIns_Inst_Sbox_14_M41 ;
    wire SubBytesIns_Inst_Sbox_14_M40 ;
    wire SubBytesIns_Inst_Sbox_14_M39 ;
    wire SubBytesIns_Inst_Sbox_14_M38 ;
    wire SubBytesIns_Inst_Sbox_14_M37 ;
    wire SubBytesIns_Inst_Sbox_14_M36 ;
    wire SubBytesIns_Inst_Sbox_14_M35 ;
    wire SubBytesIns_Inst_Sbox_14_M34 ;
    wire SubBytesIns_Inst_Sbox_14_M33 ;
    wire SubBytesIns_Inst_Sbox_14_M32 ;
    wire SubBytesIns_Inst_Sbox_14_M31 ;
    wire SubBytesIns_Inst_Sbox_14_M30 ;
    wire SubBytesIns_Inst_Sbox_14_M29 ;
    wire SubBytesIns_Inst_Sbox_14_M28 ;
    wire SubBytesIns_Inst_Sbox_14_M27 ;
    wire SubBytesIns_Inst_Sbox_14_M26 ;
    wire SubBytesIns_Inst_Sbox_14_M25 ;
    wire SubBytesIns_Inst_Sbox_14_M24 ;
    wire SubBytesIns_Inst_Sbox_14_M23 ;
    wire SubBytesIns_Inst_Sbox_14_M22 ;
    wire SubBytesIns_Inst_Sbox_14_M21 ;
    wire SubBytesIns_Inst_Sbox_14_M20 ;
    wire SubBytesIns_Inst_Sbox_14_M19 ;
    wire SubBytesIns_Inst_Sbox_14_M18 ;
    wire SubBytesIns_Inst_Sbox_14_M17 ;
    wire SubBytesIns_Inst_Sbox_14_M16 ;
    wire SubBytesIns_Inst_Sbox_14_M15 ;
    wire SubBytesIns_Inst_Sbox_14_M14 ;
    wire SubBytesIns_Inst_Sbox_14_M13 ;
    wire SubBytesIns_Inst_Sbox_14_M12 ;
    wire SubBytesIns_Inst_Sbox_14_M11 ;
    wire SubBytesIns_Inst_Sbox_14_M10 ;
    wire SubBytesIns_Inst_Sbox_14_M9 ;
    wire SubBytesIns_Inst_Sbox_14_M8 ;
    wire SubBytesIns_Inst_Sbox_14_M7 ;
    wire SubBytesIns_Inst_Sbox_14_M6 ;
    wire SubBytesIns_Inst_Sbox_14_M5 ;
    wire SubBytesIns_Inst_Sbox_14_M4 ;
    wire SubBytesIns_Inst_Sbox_14_M3 ;
    wire SubBytesIns_Inst_Sbox_14_M2 ;
    wire SubBytesIns_Inst_Sbox_14_M1 ;
    wire SubBytesIns_Inst_Sbox_14_T27 ;
    wire SubBytesIns_Inst_Sbox_14_T26 ;
    wire SubBytesIns_Inst_Sbox_14_T25 ;
    wire SubBytesIns_Inst_Sbox_14_T24 ;
    wire SubBytesIns_Inst_Sbox_14_T23 ;
    wire SubBytesIns_Inst_Sbox_14_T22 ;
    wire SubBytesIns_Inst_Sbox_14_T21 ;
    wire SubBytesIns_Inst_Sbox_14_T20 ;
    wire SubBytesIns_Inst_Sbox_14_T19 ;
    wire SubBytesIns_Inst_Sbox_14_T18 ;
    wire SubBytesIns_Inst_Sbox_14_T17 ;
    wire SubBytesIns_Inst_Sbox_14_T16 ;
    wire SubBytesIns_Inst_Sbox_14_T15 ;
    wire SubBytesIns_Inst_Sbox_14_T14 ;
    wire SubBytesIns_Inst_Sbox_14_T13 ;
    wire SubBytesIns_Inst_Sbox_14_T12 ;
    wire SubBytesIns_Inst_Sbox_14_T11 ;
    wire SubBytesIns_Inst_Sbox_14_T10 ;
    wire SubBytesIns_Inst_Sbox_14_T9 ;
    wire SubBytesIns_Inst_Sbox_14_T8 ;
    wire SubBytesIns_Inst_Sbox_14_T7 ;
    wire SubBytesIns_Inst_Sbox_14_T6 ;
    wire SubBytesIns_Inst_Sbox_14_T5 ;
    wire SubBytesIns_Inst_Sbox_14_T4 ;
    wire SubBytesIns_Inst_Sbox_14_T3 ;
    wire SubBytesIns_Inst_Sbox_14_T2 ;
    wire SubBytesIns_Inst_Sbox_14_T1 ;
    wire SubBytesIns_Inst_Sbox_15_L29 ;
    wire SubBytesIns_Inst_Sbox_15_L28 ;
    wire SubBytesIns_Inst_Sbox_15_L27 ;
    wire SubBytesIns_Inst_Sbox_15_L26 ;
    wire SubBytesIns_Inst_Sbox_15_L25 ;
    wire SubBytesIns_Inst_Sbox_15_L24 ;
    wire SubBytesIns_Inst_Sbox_15_L23 ;
    wire SubBytesIns_Inst_Sbox_15_L22 ;
    wire SubBytesIns_Inst_Sbox_15_L21 ;
    wire SubBytesIns_Inst_Sbox_15_L20 ;
    wire SubBytesIns_Inst_Sbox_15_L19 ;
    wire SubBytesIns_Inst_Sbox_15_L18 ;
    wire SubBytesIns_Inst_Sbox_15_L17 ;
    wire SubBytesIns_Inst_Sbox_15_L16 ;
    wire SubBytesIns_Inst_Sbox_15_L15 ;
    wire SubBytesIns_Inst_Sbox_15_L14 ;
    wire SubBytesIns_Inst_Sbox_15_L13 ;
    wire SubBytesIns_Inst_Sbox_15_L12 ;
    wire SubBytesIns_Inst_Sbox_15_L11 ;
    wire SubBytesIns_Inst_Sbox_15_L10 ;
    wire SubBytesIns_Inst_Sbox_15_L9 ;
    wire SubBytesIns_Inst_Sbox_15_L8 ;
    wire SubBytesIns_Inst_Sbox_15_L7 ;
    wire SubBytesIns_Inst_Sbox_15_L6 ;
    wire SubBytesIns_Inst_Sbox_15_L5 ;
    wire SubBytesIns_Inst_Sbox_15_L4 ;
    wire SubBytesIns_Inst_Sbox_15_L3 ;
    wire SubBytesIns_Inst_Sbox_15_L2 ;
    wire SubBytesIns_Inst_Sbox_15_L1 ;
    wire SubBytesIns_Inst_Sbox_15_L0 ;
    wire SubBytesIns_Inst_Sbox_15_M63 ;
    wire SubBytesIns_Inst_Sbox_15_M62 ;
    wire SubBytesIns_Inst_Sbox_15_M61 ;
    wire SubBytesIns_Inst_Sbox_15_M60 ;
    wire SubBytesIns_Inst_Sbox_15_M59 ;
    wire SubBytesIns_Inst_Sbox_15_M58 ;
    wire SubBytesIns_Inst_Sbox_15_M57 ;
    wire SubBytesIns_Inst_Sbox_15_M56 ;
    wire SubBytesIns_Inst_Sbox_15_M55 ;
    wire SubBytesIns_Inst_Sbox_15_M54 ;
    wire SubBytesIns_Inst_Sbox_15_M53 ;
    wire SubBytesIns_Inst_Sbox_15_M52 ;
    wire SubBytesIns_Inst_Sbox_15_M51 ;
    wire SubBytesIns_Inst_Sbox_15_M50 ;
    wire SubBytesIns_Inst_Sbox_15_M49 ;
    wire SubBytesIns_Inst_Sbox_15_M48 ;
    wire SubBytesIns_Inst_Sbox_15_M47 ;
    wire SubBytesIns_Inst_Sbox_15_M46 ;
    wire SubBytesIns_Inst_Sbox_15_M45 ;
    wire SubBytesIns_Inst_Sbox_15_M44 ;
    wire SubBytesIns_Inst_Sbox_15_M43 ;
    wire SubBytesIns_Inst_Sbox_15_M42 ;
    wire SubBytesIns_Inst_Sbox_15_M41 ;
    wire SubBytesIns_Inst_Sbox_15_M40 ;
    wire SubBytesIns_Inst_Sbox_15_M39 ;
    wire SubBytesIns_Inst_Sbox_15_M38 ;
    wire SubBytesIns_Inst_Sbox_15_M37 ;
    wire SubBytesIns_Inst_Sbox_15_M36 ;
    wire SubBytesIns_Inst_Sbox_15_M35 ;
    wire SubBytesIns_Inst_Sbox_15_M34 ;
    wire SubBytesIns_Inst_Sbox_15_M33 ;
    wire SubBytesIns_Inst_Sbox_15_M32 ;
    wire SubBytesIns_Inst_Sbox_15_M31 ;
    wire SubBytesIns_Inst_Sbox_15_M30 ;
    wire SubBytesIns_Inst_Sbox_15_M29 ;
    wire SubBytesIns_Inst_Sbox_15_M28 ;
    wire SubBytesIns_Inst_Sbox_15_M27 ;
    wire SubBytesIns_Inst_Sbox_15_M26 ;
    wire SubBytesIns_Inst_Sbox_15_M25 ;
    wire SubBytesIns_Inst_Sbox_15_M24 ;
    wire SubBytesIns_Inst_Sbox_15_M23 ;
    wire SubBytesIns_Inst_Sbox_15_M22 ;
    wire SubBytesIns_Inst_Sbox_15_M21 ;
    wire SubBytesIns_Inst_Sbox_15_M20 ;
    wire SubBytesIns_Inst_Sbox_15_M19 ;
    wire SubBytesIns_Inst_Sbox_15_M18 ;
    wire SubBytesIns_Inst_Sbox_15_M17 ;
    wire SubBytesIns_Inst_Sbox_15_M16 ;
    wire SubBytesIns_Inst_Sbox_15_M15 ;
    wire SubBytesIns_Inst_Sbox_15_M14 ;
    wire SubBytesIns_Inst_Sbox_15_M13 ;
    wire SubBytesIns_Inst_Sbox_15_M12 ;
    wire SubBytesIns_Inst_Sbox_15_M11 ;
    wire SubBytesIns_Inst_Sbox_15_M10 ;
    wire SubBytesIns_Inst_Sbox_15_M9 ;
    wire SubBytesIns_Inst_Sbox_15_M8 ;
    wire SubBytesIns_Inst_Sbox_15_M7 ;
    wire SubBytesIns_Inst_Sbox_15_M6 ;
    wire SubBytesIns_Inst_Sbox_15_M5 ;
    wire SubBytesIns_Inst_Sbox_15_M4 ;
    wire SubBytesIns_Inst_Sbox_15_M3 ;
    wire SubBytesIns_Inst_Sbox_15_M2 ;
    wire SubBytesIns_Inst_Sbox_15_M1 ;
    wire SubBytesIns_Inst_Sbox_15_T27 ;
    wire SubBytesIns_Inst_Sbox_15_T26 ;
    wire SubBytesIns_Inst_Sbox_15_T25 ;
    wire SubBytesIns_Inst_Sbox_15_T24 ;
    wire SubBytesIns_Inst_Sbox_15_T23 ;
    wire SubBytesIns_Inst_Sbox_15_T22 ;
    wire SubBytesIns_Inst_Sbox_15_T21 ;
    wire SubBytesIns_Inst_Sbox_15_T20 ;
    wire SubBytesIns_Inst_Sbox_15_T19 ;
    wire SubBytesIns_Inst_Sbox_15_T18 ;
    wire SubBytesIns_Inst_Sbox_15_T17 ;
    wire SubBytesIns_Inst_Sbox_15_T16 ;
    wire SubBytesIns_Inst_Sbox_15_T15 ;
    wire SubBytesIns_Inst_Sbox_15_T14 ;
    wire SubBytesIns_Inst_Sbox_15_T13 ;
    wire SubBytesIns_Inst_Sbox_15_T12 ;
    wire SubBytesIns_Inst_Sbox_15_T11 ;
    wire SubBytesIns_Inst_Sbox_15_T10 ;
    wire SubBytesIns_Inst_Sbox_15_T9 ;
    wire SubBytesIns_Inst_Sbox_15_T8 ;
    wire SubBytesIns_Inst_Sbox_15_T7 ;
    wire SubBytesIns_Inst_Sbox_15_T6 ;
    wire SubBytesIns_Inst_Sbox_15_T5 ;
    wire SubBytesIns_Inst_Sbox_15_T4 ;
    wire SubBytesIns_Inst_Sbox_15_T3 ;
    wire SubBytesIns_Inst_Sbox_15_T2 ;
    wire SubBytesIns_Inst_Sbox_15_T1 ;
    wire MixColumnsIns_MixOneColumnInst_0_n64 ;
    wire MixColumnsIns_MixOneColumnInst_0_n63 ;
    wire MixColumnsIns_MixOneColumnInst_0_n62 ;
    wire MixColumnsIns_MixOneColumnInst_0_n61 ;
    wire MixColumnsIns_MixOneColumnInst_0_n60 ;
    wire MixColumnsIns_MixOneColumnInst_0_n59 ;
    wire MixColumnsIns_MixOneColumnInst_0_n58 ;
    wire MixColumnsIns_MixOneColumnInst_0_n57 ;
    wire MixColumnsIns_MixOneColumnInst_0_n56 ;
    wire MixColumnsIns_MixOneColumnInst_0_n55 ;
    wire MixColumnsIns_MixOneColumnInst_0_n54 ;
    wire MixColumnsIns_MixOneColumnInst_0_n53 ;
    wire MixColumnsIns_MixOneColumnInst_0_n52 ;
    wire MixColumnsIns_MixOneColumnInst_0_n51 ;
    wire MixColumnsIns_MixOneColumnInst_0_n50 ;
    wire MixColumnsIns_MixOneColumnInst_0_n49 ;
    wire MixColumnsIns_MixOneColumnInst_0_n48 ;
    wire MixColumnsIns_MixOneColumnInst_0_n47 ;
    wire MixColumnsIns_MixOneColumnInst_0_n46 ;
    wire MixColumnsIns_MixOneColumnInst_0_n45 ;
    wire MixColumnsIns_MixOneColumnInst_0_n44 ;
    wire MixColumnsIns_MixOneColumnInst_0_n43 ;
    wire MixColumnsIns_MixOneColumnInst_0_n42 ;
    wire MixColumnsIns_MixOneColumnInst_0_n41 ;
    wire MixColumnsIns_MixOneColumnInst_0_n40 ;
    wire MixColumnsIns_MixOneColumnInst_0_n39 ;
    wire MixColumnsIns_MixOneColumnInst_0_n38 ;
    wire MixColumnsIns_MixOneColumnInst_0_n37 ;
    wire MixColumnsIns_MixOneColumnInst_0_n36 ;
    wire MixColumnsIns_MixOneColumnInst_0_n35 ;
    wire MixColumnsIns_MixOneColumnInst_0_n34 ;
    wire MixColumnsIns_MixOneColumnInst_0_n33 ;
    wire MixColumnsIns_MixOneColumnInst_0_n32 ;
    wire MixColumnsIns_MixOneColumnInst_0_n31 ;
    wire MixColumnsIns_MixOneColumnInst_0_n30 ;
    wire MixColumnsIns_MixOneColumnInst_0_n29 ;
    wire MixColumnsIns_MixOneColumnInst_0_n28 ;
    wire MixColumnsIns_MixOneColumnInst_0_n27 ;
    wire MixColumnsIns_MixOneColumnInst_0_n26 ;
    wire MixColumnsIns_MixOneColumnInst_0_n25 ;
    wire MixColumnsIns_MixOneColumnInst_0_n24 ;
    wire MixColumnsIns_MixOneColumnInst_0_n23 ;
    wire MixColumnsIns_MixOneColumnInst_0_n22 ;
    wire MixColumnsIns_MixOneColumnInst_0_n21 ;
    wire MixColumnsIns_MixOneColumnInst_0_n20 ;
    wire MixColumnsIns_MixOneColumnInst_0_n19 ;
    wire MixColumnsIns_MixOneColumnInst_0_n18 ;
    wire MixColumnsIns_MixOneColumnInst_0_n17 ;
    wire MixColumnsIns_MixOneColumnInst_0_n16 ;
    wire MixColumnsIns_MixOneColumnInst_0_n15 ;
    wire MixColumnsIns_MixOneColumnInst_0_n14 ;
    wire MixColumnsIns_MixOneColumnInst_0_n13 ;
    wire MixColumnsIns_MixOneColumnInst_0_n12 ;
    wire MixColumnsIns_MixOneColumnInst_0_n11 ;
    wire MixColumnsIns_MixOneColumnInst_0_n10 ;
    wire MixColumnsIns_MixOneColumnInst_0_n9 ;
    wire MixColumnsIns_MixOneColumnInst_0_n8 ;
    wire MixColumnsIns_MixOneColumnInst_0_n7 ;
    wire MixColumnsIns_MixOneColumnInst_0_n6 ;
    wire MixColumnsIns_MixOneColumnInst_0_n5 ;
    wire MixColumnsIns_MixOneColumnInst_0_n4 ;
    wire MixColumnsIns_MixOneColumnInst_0_n3 ;
    wire MixColumnsIns_MixOneColumnInst_0_n2 ;
    wire MixColumnsIns_MixOneColumnInst_0_n1 ;
    wire MixColumnsIns_MixOneColumnInst_1_n64 ;
    wire MixColumnsIns_MixOneColumnInst_1_n63 ;
    wire MixColumnsIns_MixOneColumnInst_1_n62 ;
    wire MixColumnsIns_MixOneColumnInst_1_n61 ;
    wire MixColumnsIns_MixOneColumnInst_1_n60 ;
    wire MixColumnsIns_MixOneColumnInst_1_n59 ;
    wire MixColumnsIns_MixOneColumnInst_1_n58 ;
    wire MixColumnsIns_MixOneColumnInst_1_n57 ;
    wire MixColumnsIns_MixOneColumnInst_1_n56 ;
    wire MixColumnsIns_MixOneColumnInst_1_n55 ;
    wire MixColumnsIns_MixOneColumnInst_1_n54 ;
    wire MixColumnsIns_MixOneColumnInst_1_n53 ;
    wire MixColumnsIns_MixOneColumnInst_1_n52 ;
    wire MixColumnsIns_MixOneColumnInst_1_n51 ;
    wire MixColumnsIns_MixOneColumnInst_1_n50 ;
    wire MixColumnsIns_MixOneColumnInst_1_n49 ;
    wire MixColumnsIns_MixOneColumnInst_1_n48 ;
    wire MixColumnsIns_MixOneColumnInst_1_n47 ;
    wire MixColumnsIns_MixOneColumnInst_1_n46 ;
    wire MixColumnsIns_MixOneColumnInst_1_n45 ;
    wire MixColumnsIns_MixOneColumnInst_1_n44 ;
    wire MixColumnsIns_MixOneColumnInst_1_n43 ;
    wire MixColumnsIns_MixOneColumnInst_1_n42 ;
    wire MixColumnsIns_MixOneColumnInst_1_n41 ;
    wire MixColumnsIns_MixOneColumnInst_1_n40 ;
    wire MixColumnsIns_MixOneColumnInst_1_n39 ;
    wire MixColumnsIns_MixOneColumnInst_1_n38 ;
    wire MixColumnsIns_MixOneColumnInst_1_n37 ;
    wire MixColumnsIns_MixOneColumnInst_1_n36 ;
    wire MixColumnsIns_MixOneColumnInst_1_n35 ;
    wire MixColumnsIns_MixOneColumnInst_1_n34 ;
    wire MixColumnsIns_MixOneColumnInst_1_n33 ;
    wire MixColumnsIns_MixOneColumnInst_1_n32 ;
    wire MixColumnsIns_MixOneColumnInst_1_n31 ;
    wire MixColumnsIns_MixOneColumnInst_1_n30 ;
    wire MixColumnsIns_MixOneColumnInst_1_n29 ;
    wire MixColumnsIns_MixOneColumnInst_1_n28 ;
    wire MixColumnsIns_MixOneColumnInst_1_n27 ;
    wire MixColumnsIns_MixOneColumnInst_1_n26 ;
    wire MixColumnsIns_MixOneColumnInst_1_n25 ;
    wire MixColumnsIns_MixOneColumnInst_1_n24 ;
    wire MixColumnsIns_MixOneColumnInst_1_n23 ;
    wire MixColumnsIns_MixOneColumnInst_1_n22 ;
    wire MixColumnsIns_MixOneColumnInst_1_n21 ;
    wire MixColumnsIns_MixOneColumnInst_1_n20 ;
    wire MixColumnsIns_MixOneColumnInst_1_n19 ;
    wire MixColumnsIns_MixOneColumnInst_1_n18 ;
    wire MixColumnsIns_MixOneColumnInst_1_n17 ;
    wire MixColumnsIns_MixOneColumnInst_1_n16 ;
    wire MixColumnsIns_MixOneColumnInst_1_n15 ;
    wire MixColumnsIns_MixOneColumnInst_1_n14 ;
    wire MixColumnsIns_MixOneColumnInst_1_n13 ;
    wire MixColumnsIns_MixOneColumnInst_1_n12 ;
    wire MixColumnsIns_MixOneColumnInst_1_n11 ;
    wire MixColumnsIns_MixOneColumnInst_1_n10 ;
    wire MixColumnsIns_MixOneColumnInst_1_n9 ;
    wire MixColumnsIns_MixOneColumnInst_1_n8 ;
    wire MixColumnsIns_MixOneColumnInst_1_n7 ;
    wire MixColumnsIns_MixOneColumnInst_1_n6 ;
    wire MixColumnsIns_MixOneColumnInst_1_n5 ;
    wire MixColumnsIns_MixOneColumnInst_1_n4 ;
    wire MixColumnsIns_MixOneColumnInst_1_n3 ;
    wire MixColumnsIns_MixOneColumnInst_1_n2 ;
    wire MixColumnsIns_MixOneColumnInst_1_n1 ;
    wire MixColumnsIns_MixOneColumnInst_2_n64 ;
    wire MixColumnsIns_MixOneColumnInst_2_n63 ;
    wire MixColumnsIns_MixOneColumnInst_2_n62 ;
    wire MixColumnsIns_MixOneColumnInst_2_n61 ;
    wire MixColumnsIns_MixOneColumnInst_2_n60 ;
    wire MixColumnsIns_MixOneColumnInst_2_n59 ;
    wire MixColumnsIns_MixOneColumnInst_2_n58 ;
    wire MixColumnsIns_MixOneColumnInst_2_n57 ;
    wire MixColumnsIns_MixOneColumnInst_2_n56 ;
    wire MixColumnsIns_MixOneColumnInst_2_n55 ;
    wire MixColumnsIns_MixOneColumnInst_2_n54 ;
    wire MixColumnsIns_MixOneColumnInst_2_n53 ;
    wire MixColumnsIns_MixOneColumnInst_2_n52 ;
    wire MixColumnsIns_MixOneColumnInst_2_n51 ;
    wire MixColumnsIns_MixOneColumnInst_2_n50 ;
    wire MixColumnsIns_MixOneColumnInst_2_n49 ;
    wire MixColumnsIns_MixOneColumnInst_2_n48 ;
    wire MixColumnsIns_MixOneColumnInst_2_n47 ;
    wire MixColumnsIns_MixOneColumnInst_2_n46 ;
    wire MixColumnsIns_MixOneColumnInst_2_n45 ;
    wire MixColumnsIns_MixOneColumnInst_2_n44 ;
    wire MixColumnsIns_MixOneColumnInst_2_n43 ;
    wire MixColumnsIns_MixOneColumnInst_2_n42 ;
    wire MixColumnsIns_MixOneColumnInst_2_n41 ;
    wire MixColumnsIns_MixOneColumnInst_2_n40 ;
    wire MixColumnsIns_MixOneColumnInst_2_n39 ;
    wire MixColumnsIns_MixOneColumnInst_2_n38 ;
    wire MixColumnsIns_MixOneColumnInst_2_n37 ;
    wire MixColumnsIns_MixOneColumnInst_2_n36 ;
    wire MixColumnsIns_MixOneColumnInst_2_n35 ;
    wire MixColumnsIns_MixOneColumnInst_2_n34 ;
    wire MixColumnsIns_MixOneColumnInst_2_n33 ;
    wire MixColumnsIns_MixOneColumnInst_2_n32 ;
    wire MixColumnsIns_MixOneColumnInst_2_n31 ;
    wire MixColumnsIns_MixOneColumnInst_2_n30 ;
    wire MixColumnsIns_MixOneColumnInst_2_n29 ;
    wire MixColumnsIns_MixOneColumnInst_2_n28 ;
    wire MixColumnsIns_MixOneColumnInst_2_n27 ;
    wire MixColumnsIns_MixOneColumnInst_2_n26 ;
    wire MixColumnsIns_MixOneColumnInst_2_n25 ;
    wire MixColumnsIns_MixOneColumnInst_2_n24 ;
    wire MixColumnsIns_MixOneColumnInst_2_n23 ;
    wire MixColumnsIns_MixOneColumnInst_2_n22 ;
    wire MixColumnsIns_MixOneColumnInst_2_n21 ;
    wire MixColumnsIns_MixOneColumnInst_2_n20 ;
    wire MixColumnsIns_MixOneColumnInst_2_n19 ;
    wire MixColumnsIns_MixOneColumnInst_2_n18 ;
    wire MixColumnsIns_MixOneColumnInst_2_n17 ;
    wire MixColumnsIns_MixOneColumnInst_2_n16 ;
    wire MixColumnsIns_MixOneColumnInst_2_n15 ;
    wire MixColumnsIns_MixOneColumnInst_2_n14 ;
    wire MixColumnsIns_MixOneColumnInst_2_n13 ;
    wire MixColumnsIns_MixOneColumnInst_2_n12 ;
    wire MixColumnsIns_MixOneColumnInst_2_n11 ;
    wire MixColumnsIns_MixOneColumnInst_2_n10 ;
    wire MixColumnsIns_MixOneColumnInst_2_n9 ;
    wire MixColumnsIns_MixOneColumnInst_2_n8 ;
    wire MixColumnsIns_MixOneColumnInst_2_n7 ;
    wire MixColumnsIns_MixOneColumnInst_2_n6 ;
    wire MixColumnsIns_MixOneColumnInst_2_n5 ;
    wire MixColumnsIns_MixOneColumnInst_2_n4 ;
    wire MixColumnsIns_MixOneColumnInst_2_n3 ;
    wire MixColumnsIns_MixOneColumnInst_2_n2 ;
    wire MixColumnsIns_MixOneColumnInst_2_n1 ;
    wire MixColumnsIns_MixOneColumnInst_3_n64 ;
    wire MixColumnsIns_MixOneColumnInst_3_n63 ;
    wire MixColumnsIns_MixOneColumnInst_3_n62 ;
    wire MixColumnsIns_MixOneColumnInst_3_n61 ;
    wire MixColumnsIns_MixOneColumnInst_3_n60 ;
    wire MixColumnsIns_MixOneColumnInst_3_n59 ;
    wire MixColumnsIns_MixOneColumnInst_3_n58 ;
    wire MixColumnsIns_MixOneColumnInst_3_n57 ;
    wire MixColumnsIns_MixOneColumnInst_3_n56 ;
    wire MixColumnsIns_MixOneColumnInst_3_n55 ;
    wire MixColumnsIns_MixOneColumnInst_3_n54 ;
    wire MixColumnsIns_MixOneColumnInst_3_n53 ;
    wire MixColumnsIns_MixOneColumnInst_3_n52 ;
    wire MixColumnsIns_MixOneColumnInst_3_n51 ;
    wire MixColumnsIns_MixOneColumnInst_3_n50 ;
    wire MixColumnsIns_MixOneColumnInst_3_n49 ;
    wire MixColumnsIns_MixOneColumnInst_3_n48 ;
    wire MixColumnsIns_MixOneColumnInst_3_n47 ;
    wire MixColumnsIns_MixOneColumnInst_3_n46 ;
    wire MixColumnsIns_MixOneColumnInst_3_n45 ;
    wire MixColumnsIns_MixOneColumnInst_3_n44 ;
    wire MixColumnsIns_MixOneColumnInst_3_n43 ;
    wire MixColumnsIns_MixOneColumnInst_3_n42 ;
    wire MixColumnsIns_MixOneColumnInst_3_n41 ;
    wire MixColumnsIns_MixOneColumnInst_3_n40 ;
    wire MixColumnsIns_MixOneColumnInst_3_n39 ;
    wire MixColumnsIns_MixOneColumnInst_3_n38 ;
    wire MixColumnsIns_MixOneColumnInst_3_n37 ;
    wire MixColumnsIns_MixOneColumnInst_3_n36 ;
    wire MixColumnsIns_MixOneColumnInst_3_n35 ;
    wire MixColumnsIns_MixOneColumnInst_3_n34 ;
    wire MixColumnsIns_MixOneColumnInst_3_n33 ;
    wire MixColumnsIns_MixOneColumnInst_3_n32 ;
    wire MixColumnsIns_MixOneColumnInst_3_n31 ;
    wire MixColumnsIns_MixOneColumnInst_3_n30 ;
    wire MixColumnsIns_MixOneColumnInst_3_n29 ;
    wire MixColumnsIns_MixOneColumnInst_3_n28 ;
    wire MixColumnsIns_MixOneColumnInst_3_n27 ;
    wire MixColumnsIns_MixOneColumnInst_3_n26 ;
    wire MixColumnsIns_MixOneColumnInst_3_n25 ;
    wire MixColumnsIns_MixOneColumnInst_3_n24 ;
    wire MixColumnsIns_MixOneColumnInst_3_n23 ;
    wire MixColumnsIns_MixOneColumnInst_3_n22 ;
    wire MixColumnsIns_MixOneColumnInst_3_n21 ;
    wire MixColumnsIns_MixOneColumnInst_3_n20 ;
    wire MixColumnsIns_MixOneColumnInst_3_n19 ;
    wire MixColumnsIns_MixOneColumnInst_3_n18 ;
    wire MixColumnsIns_MixOneColumnInst_3_n17 ;
    wire MixColumnsIns_MixOneColumnInst_3_n16 ;
    wire MixColumnsIns_MixOneColumnInst_3_n15 ;
    wire MixColumnsIns_MixOneColumnInst_3_n14 ;
    wire MixColumnsIns_MixOneColumnInst_3_n13 ;
    wire MixColumnsIns_MixOneColumnInst_3_n12 ;
    wire MixColumnsIns_MixOneColumnInst_3_n11 ;
    wire MixColumnsIns_MixOneColumnInst_3_n10 ;
    wire MixColumnsIns_MixOneColumnInst_3_n9 ;
    wire MixColumnsIns_MixOneColumnInst_3_n8 ;
    wire MixColumnsIns_MixOneColumnInst_3_n7 ;
    wire MixColumnsIns_MixOneColumnInst_3_n6 ;
    wire MixColumnsIns_MixOneColumnInst_3_n5 ;
    wire MixColumnsIns_MixOneColumnInst_3_n4 ;
    wire MixColumnsIns_MixOneColumnInst_3_n3 ;
    wire MixColumnsIns_MixOneColumnInst_3_n2 ;
    wire MixColumnsIns_MixOneColumnInst_3_n1 ;
    wire KeyReg_Inst_ff_SDE_0_next_state ;
    wire KeyReg_Inst_ff_SDE_1_next_state ;
    wire KeyReg_Inst_ff_SDE_2_next_state ;
    wire KeyReg_Inst_ff_SDE_3_next_state ;
    wire KeyReg_Inst_ff_SDE_4_next_state ;
    wire KeyReg_Inst_ff_SDE_5_next_state ;
    wire KeyReg_Inst_ff_SDE_6_next_state ;
    wire KeyReg_Inst_ff_SDE_7_next_state ;
    wire KeyReg_Inst_ff_SDE_8_next_state ;
    wire KeyReg_Inst_ff_SDE_9_next_state ;
    wire KeyReg_Inst_ff_SDE_10_next_state ;
    wire KeyReg_Inst_ff_SDE_11_next_state ;
    wire KeyReg_Inst_ff_SDE_12_next_state ;
    wire KeyReg_Inst_ff_SDE_13_next_state ;
    wire KeyReg_Inst_ff_SDE_14_next_state ;
    wire KeyReg_Inst_ff_SDE_15_next_state ;
    wire KeyReg_Inst_ff_SDE_16_next_state ;
    wire KeyReg_Inst_ff_SDE_17_next_state ;
    wire KeyReg_Inst_ff_SDE_18_next_state ;
    wire KeyReg_Inst_ff_SDE_19_next_state ;
    wire KeyReg_Inst_ff_SDE_20_next_state ;
    wire KeyReg_Inst_ff_SDE_21_next_state ;
    wire KeyReg_Inst_ff_SDE_22_next_state ;
    wire KeyReg_Inst_ff_SDE_23_next_state ;
    wire KeyReg_Inst_ff_SDE_24_next_state ;
    wire KeyReg_Inst_ff_SDE_25_next_state ;
    wire KeyReg_Inst_ff_SDE_26_next_state ;
    wire KeyReg_Inst_ff_SDE_27_next_state ;
    wire KeyReg_Inst_ff_SDE_28_next_state ;
    wire KeyReg_Inst_ff_SDE_29_next_state ;
    wire KeyReg_Inst_ff_SDE_30_next_state ;
    wire KeyReg_Inst_ff_SDE_31_next_state ;
    wire KeyReg_Inst_ff_SDE_32_next_state ;
    wire KeyReg_Inst_ff_SDE_33_next_state ;
    wire KeyReg_Inst_ff_SDE_34_next_state ;
    wire KeyReg_Inst_ff_SDE_35_next_state ;
    wire KeyReg_Inst_ff_SDE_36_next_state ;
    wire KeyReg_Inst_ff_SDE_37_next_state ;
    wire KeyReg_Inst_ff_SDE_38_next_state ;
    wire KeyReg_Inst_ff_SDE_39_next_state ;
    wire KeyReg_Inst_ff_SDE_40_next_state ;
    wire KeyReg_Inst_ff_SDE_41_next_state ;
    wire KeyReg_Inst_ff_SDE_42_next_state ;
    wire KeyReg_Inst_ff_SDE_43_next_state ;
    wire KeyReg_Inst_ff_SDE_44_next_state ;
    wire KeyReg_Inst_ff_SDE_45_next_state ;
    wire KeyReg_Inst_ff_SDE_46_next_state ;
    wire KeyReg_Inst_ff_SDE_47_next_state ;
    wire KeyReg_Inst_ff_SDE_48_next_state ;
    wire KeyReg_Inst_ff_SDE_49_next_state ;
    wire KeyReg_Inst_ff_SDE_50_next_state ;
    wire KeyReg_Inst_ff_SDE_51_next_state ;
    wire KeyReg_Inst_ff_SDE_52_next_state ;
    wire KeyReg_Inst_ff_SDE_53_next_state ;
    wire KeyReg_Inst_ff_SDE_54_next_state ;
    wire KeyReg_Inst_ff_SDE_55_next_state ;
    wire KeyReg_Inst_ff_SDE_56_next_state ;
    wire KeyReg_Inst_ff_SDE_57_next_state ;
    wire KeyReg_Inst_ff_SDE_58_next_state ;
    wire KeyReg_Inst_ff_SDE_59_next_state ;
    wire KeyReg_Inst_ff_SDE_60_next_state ;
    wire KeyReg_Inst_ff_SDE_61_next_state ;
    wire KeyReg_Inst_ff_SDE_62_next_state ;
    wire KeyReg_Inst_ff_SDE_63_next_state ;
    wire KeyReg_Inst_ff_SDE_64_next_state ;
    wire KeyReg_Inst_ff_SDE_65_next_state ;
    wire KeyReg_Inst_ff_SDE_66_next_state ;
    wire KeyReg_Inst_ff_SDE_67_next_state ;
    wire KeyReg_Inst_ff_SDE_68_next_state ;
    wire KeyReg_Inst_ff_SDE_69_next_state ;
    wire KeyReg_Inst_ff_SDE_70_next_state ;
    wire KeyReg_Inst_ff_SDE_71_next_state ;
    wire KeyReg_Inst_ff_SDE_72_next_state ;
    wire KeyReg_Inst_ff_SDE_73_next_state ;
    wire KeyReg_Inst_ff_SDE_74_next_state ;
    wire KeyReg_Inst_ff_SDE_75_next_state ;
    wire KeyReg_Inst_ff_SDE_76_next_state ;
    wire KeyReg_Inst_ff_SDE_77_next_state ;
    wire KeyReg_Inst_ff_SDE_78_next_state ;
    wire KeyReg_Inst_ff_SDE_79_next_state ;
    wire KeyReg_Inst_ff_SDE_80_next_state ;
    wire KeyReg_Inst_ff_SDE_81_next_state ;
    wire KeyReg_Inst_ff_SDE_82_next_state ;
    wire KeyReg_Inst_ff_SDE_83_next_state ;
    wire KeyReg_Inst_ff_SDE_84_next_state ;
    wire KeyReg_Inst_ff_SDE_85_next_state ;
    wire KeyReg_Inst_ff_SDE_86_next_state ;
    wire KeyReg_Inst_ff_SDE_87_next_state ;
    wire KeyReg_Inst_ff_SDE_88_next_state ;
    wire KeyReg_Inst_ff_SDE_89_next_state ;
    wire KeyReg_Inst_ff_SDE_90_next_state ;
    wire KeyReg_Inst_ff_SDE_91_next_state ;
    wire KeyReg_Inst_ff_SDE_92_next_state ;
    wire KeyReg_Inst_ff_SDE_93_next_state ;
    wire KeyReg_Inst_ff_SDE_94_next_state ;
    wire KeyReg_Inst_ff_SDE_95_next_state ;
    wire KeyReg_Inst_ff_SDE_96_next_state ;
    wire KeyReg_Inst_ff_SDE_97_next_state ;
    wire KeyReg_Inst_ff_SDE_98_next_state ;
    wire KeyReg_Inst_ff_SDE_99_next_state ;
    wire KeyReg_Inst_ff_SDE_100_next_state ;
    wire KeyReg_Inst_ff_SDE_101_next_state ;
    wire KeyReg_Inst_ff_SDE_102_next_state ;
    wire KeyReg_Inst_ff_SDE_103_next_state ;
    wire KeyReg_Inst_ff_SDE_104_next_state ;
    wire KeyReg_Inst_ff_SDE_105_next_state ;
    wire KeyReg_Inst_ff_SDE_106_next_state ;
    wire KeyReg_Inst_ff_SDE_107_next_state ;
    wire KeyReg_Inst_ff_SDE_108_next_state ;
    wire KeyReg_Inst_ff_SDE_109_next_state ;
    wire KeyReg_Inst_ff_SDE_110_next_state ;
    wire KeyReg_Inst_ff_SDE_111_next_state ;
    wire KeyReg_Inst_ff_SDE_112_next_state ;
    wire KeyReg_Inst_ff_SDE_113_next_state ;
    wire KeyReg_Inst_ff_SDE_114_next_state ;
    wire KeyReg_Inst_ff_SDE_115_next_state ;
    wire KeyReg_Inst_ff_SDE_116_next_state ;
    wire KeyReg_Inst_ff_SDE_117_next_state ;
    wire KeyReg_Inst_ff_SDE_118_next_state ;
    wire KeyReg_Inst_ff_SDE_119_next_state ;
    wire KeyReg_Inst_ff_SDE_120_next_state ;
    wire KeyReg_Inst_ff_SDE_121_next_state ;
    wire KeyReg_Inst_ff_SDE_122_next_state ;
    wire KeyReg_Inst_ff_SDE_123_next_state ;
    wire KeyReg_Inst_ff_SDE_124_next_state ;
    wire KeyReg_Inst_ff_SDE_125_next_state ;
    wire KeyReg_Inst_ff_SDE_126_next_state ;
    wire KeyReg_Inst_ff_SDE_127_next_state ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_ ;
    wire KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_ ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2 ;
    wire KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1 ;
    wire RoundCounterIns_n13 ;
    wire RoundCounterIns_n12 ;
    wire RoundCounterIns_n11 ;
    wire RoundCounterIns_n10 ;
    wire RoundCounterIns_n9 ;
    wire RoundCounterIns_n8 ;
    wire RoundCounterIns_n7 ;
    wire RoundCounterIns_n4 ;
    wire RoundCounterIns_n3 ;
    wire RoundCounterIns_n2 ;
    wire RoundCounterIns_n1 ;
    wire RoundCounterIns_N10 ;
    wire RoundCounterIns_n5 ;
    wire RoundCounterIns_N8 ;
    wire RoundCounterIns_n6 ;
    wire RoundCounterIns_N7 ;
    wire [127:0] RoundOutput ;
    wire [127:0] RoundInput ;
    wire [123:0] MixColumnsInput ;
    wire [127:0] MixColumnsOutput ;
    wire [127:0] KeyExpansionOutput ;
    wire [127:0] RoundKey ;
    wire [5:0] Rcon ;
    wire [3:0] RoundCounter ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_0_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_1_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_2_DoubleBytes ;
    wire [31:0] MixColumnsIns_MixOneColumnInst_3_DoubleBytes ;
    wire [31:0] KeyExpansionIns_tmp ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;
    wire new_AGEMA_signal_5184 ;
    wire new_AGEMA_signal_5188 ;
    wire new_AGEMA_signal_5189 ;
    wire new_AGEMA_signal_5190 ;
    wire new_AGEMA_signal_5191 ;
    wire new_AGEMA_signal_5192 ;
    wire new_AGEMA_signal_5193 ;
    wire new_AGEMA_signal_5197 ;
    wire new_AGEMA_signal_5198 ;
    wire new_AGEMA_signal_5199 ;
    wire new_AGEMA_signal_5200 ;
    wire new_AGEMA_signal_5201 ;
    wire new_AGEMA_signal_5202 ;
    wire new_AGEMA_signal_5206 ;
    wire new_AGEMA_signal_5207 ;
    wire new_AGEMA_signal_5208 ;
    wire new_AGEMA_signal_5209 ;
    wire new_AGEMA_signal_5210 ;
    wire new_AGEMA_signal_5211 ;
    wire new_AGEMA_signal_5215 ;
    wire new_AGEMA_signal_5216 ;
    wire new_AGEMA_signal_5217 ;
    wire new_AGEMA_signal_5218 ;
    wire new_AGEMA_signal_5219 ;
    wire new_AGEMA_signal_5220 ;
    wire new_AGEMA_signal_5224 ;
    wire new_AGEMA_signal_5225 ;
    wire new_AGEMA_signal_5226 ;
    wire new_AGEMA_signal_5227 ;
    wire new_AGEMA_signal_5228 ;
    wire new_AGEMA_signal_5229 ;
    wire new_AGEMA_signal_5233 ;
    wire new_AGEMA_signal_5234 ;
    wire new_AGEMA_signal_5235 ;
    wire new_AGEMA_signal_5236 ;
    wire new_AGEMA_signal_5237 ;
    wire new_AGEMA_signal_5238 ;
    wire new_AGEMA_signal_5242 ;
    wire new_AGEMA_signal_5243 ;
    wire new_AGEMA_signal_5244 ;
    wire new_AGEMA_signal_5245 ;
    wire new_AGEMA_signal_5246 ;
    wire new_AGEMA_signal_5247 ;
    wire new_AGEMA_signal_5251 ;
    wire new_AGEMA_signal_5252 ;
    wire new_AGEMA_signal_5253 ;
    wire new_AGEMA_signal_5254 ;
    wire new_AGEMA_signal_5255 ;
    wire new_AGEMA_signal_5256 ;
    wire new_AGEMA_signal_5260 ;
    wire new_AGEMA_signal_5261 ;
    wire new_AGEMA_signal_5262 ;
    wire new_AGEMA_signal_5263 ;
    wire new_AGEMA_signal_5264 ;
    wire new_AGEMA_signal_5265 ;
    wire new_AGEMA_signal_5269 ;
    wire new_AGEMA_signal_5270 ;
    wire new_AGEMA_signal_5271 ;
    wire new_AGEMA_signal_5272 ;
    wire new_AGEMA_signal_5273 ;
    wire new_AGEMA_signal_5274 ;
    wire new_AGEMA_signal_5278 ;
    wire new_AGEMA_signal_5279 ;
    wire new_AGEMA_signal_5280 ;
    wire new_AGEMA_signal_5281 ;
    wire new_AGEMA_signal_5282 ;
    wire new_AGEMA_signal_5283 ;
    wire new_AGEMA_signal_5287 ;
    wire new_AGEMA_signal_5288 ;
    wire new_AGEMA_signal_5289 ;
    wire new_AGEMA_signal_5290 ;
    wire new_AGEMA_signal_5291 ;
    wire new_AGEMA_signal_5292 ;
    wire new_AGEMA_signal_5296 ;
    wire new_AGEMA_signal_5297 ;
    wire new_AGEMA_signal_5298 ;
    wire new_AGEMA_signal_5299 ;
    wire new_AGEMA_signal_5300 ;
    wire new_AGEMA_signal_5301 ;
    wire new_AGEMA_signal_5305 ;
    wire new_AGEMA_signal_5306 ;
    wire new_AGEMA_signal_5307 ;
    wire new_AGEMA_signal_5308 ;
    wire new_AGEMA_signal_5309 ;
    wire new_AGEMA_signal_5310 ;
    wire new_AGEMA_signal_5314 ;
    wire new_AGEMA_signal_5315 ;
    wire new_AGEMA_signal_5316 ;
    wire new_AGEMA_signal_5317 ;
    wire new_AGEMA_signal_5318 ;
    wire new_AGEMA_signal_5319 ;
    wire new_AGEMA_signal_5323 ;
    wire new_AGEMA_signal_5324 ;
    wire new_AGEMA_signal_5325 ;
    wire new_AGEMA_signal_5326 ;
    wire new_AGEMA_signal_5327 ;
    wire new_AGEMA_signal_5328 ;
    wire new_AGEMA_signal_5332 ;
    wire new_AGEMA_signal_5333 ;
    wire new_AGEMA_signal_5334 ;
    wire new_AGEMA_signal_5335 ;
    wire new_AGEMA_signal_5336 ;
    wire new_AGEMA_signal_5337 ;
    wire new_AGEMA_signal_5341 ;
    wire new_AGEMA_signal_5342 ;
    wire new_AGEMA_signal_5343 ;
    wire new_AGEMA_signal_5344 ;
    wire new_AGEMA_signal_5345 ;
    wire new_AGEMA_signal_5346 ;
    wire new_AGEMA_signal_5350 ;
    wire new_AGEMA_signal_5351 ;
    wire new_AGEMA_signal_5352 ;
    wire new_AGEMA_signal_5353 ;
    wire new_AGEMA_signal_5354 ;
    wire new_AGEMA_signal_5355 ;
    wire new_AGEMA_signal_5359 ;
    wire new_AGEMA_signal_5360 ;
    wire new_AGEMA_signal_5361 ;
    wire new_AGEMA_signal_5362 ;
    wire new_AGEMA_signal_5363 ;
    wire new_AGEMA_signal_5364 ;
    wire new_AGEMA_signal_5368 ;
    wire new_AGEMA_signal_5369 ;
    wire new_AGEMA_signal_5370 ;
    wire new_AGEMA_signal_5371 ;
    wire new_AGEMA_signal_5372 ;
    wire new_AGEMA_signal_5373 ;
    wire new_AGEMA_signal_5377 ;
    wire new_AGEMA_signal_5378 ;
    wire new_AGEMA_signal_5379 ;
    wire new_AGEMA_signal_5380 ;
    wire new_AGEMA_signal_5381 ;
    wire new_AGEMA_signal_5382 ;
    wire new_AGEMA_signal_5386 ;
    wire new_AGEMA_signal_5387 ;
    wire new_AGEMA_signal_5388 ;
    wire new_AGEMA_signal_5389 ;
    wire new_AGEMA_signal_5390 ;
    wire new_AGEMA_signal_5391 ;
    wire new_AGEMA_signal_5395 ;
    wire new_AGEMA_signal_5396 ;
    wire new_AGEMA_signal_5397 ;
    wire new_AGEMA_signal_5398 ;
    wire new_AGEMA_signal_5399 ;
    wire new_AGEMA_signal_5400 ;
    wire new_AGEMA_signal_5404 ;
    wire new_AGEMA_signal_5405 ;
    wire new_AGEMA_signal_5406 ;
    wire new_AGEMA_signal_5407 ;
    wire new_AGEMA_signal_5408 ;
    wire new_AGEMA_signal_5409 ;
    wire new_AGEMA_signal_5413 ;
    wire new_AGEMA_signal_5414 ;
    wire new_AGEMA_signal_5415 ;
    wire new_AGEMA_signal_5416 ;
    wire new_AGEMA_signal_5417 ;
    wire new_AGEMA_signal_5418 ;
    wire new_AGEMA_signal_5422 ;
    wire new_AGEMA_signal_5423 ;
    wire new_AGEMA_signal_5424 ;
    wire new_AGEMA_signal_5425 ;
    wire new_AGEMA_signal_5426 ;
    wire new_AGEMA_signal_5427 ;
    wire new_AGEMA_signal_5431 ;
    wire new_AGEMA_signal_5432 ;
    wire new_AGEMA_signal_5433 ;
    wire new_AGEMA_signal_5434 ;
    wire new_AGEMA_signal_5435 ;
    wire new_AGEMA_signal_5436 ;
    wire new_AGEMA_signal_5440 ;
    wire new_AGEMA_signal_5441 ;
    wire new_AGEMA_signal_5442 ;
    wire new_AGEMA_signal_5443 ;
    wire new_AGEMA_signal_5444 ;
    wire new_AGEMA_signal_5445 ;
    wire new_AGEMA_signal_5449 ;
    wire new_AGEMA_signal_5450 ;
    wire new_AGEMA_signal_5451 ;
    wire new_AGEMA_signal_5452 ;
    wire new_AGEMA_signal_5453 ;
    wire new_AGEMA_signal_5454 ;
    wire new_AGEMA_signal_5458 ;
    wire new_AGEMA_signal_5459 ;
    wire new_AGEMA_signal_5460 ;
    wire new_AGEMA_signal_5461 ;
    wire new_AGEMA_signal_5462 ;
    wire new_AGEMA_signal_5463 ;
    wire new_AGEMA_signal_5467 ;
    wire new_AGEMA_signal_5468 ;
    wire new_AGEMA_signal_5469 ;
    wire new_AGEMA_signal_5470 ;
    wire new_AGEMA_signal_5471 ;
    wire new_AGEMA_signal_5472 ;
    wire new_AGEMA_signal_5476 ;
    wire new_AGEMA_signal_5477 ;
    wire new_AGEMA_signal_5478 ;
    wire new_AGEMA_signal_5479 ;
    wire new_AGEMA_signal_5480 ;
    wire new_AGEMA_signal_5481 ;
    wire new_AGEMA_signal_5485 ;
    wire new_AGEMA_signal_5486 ;
    wire new_AGEMA_signal_5487 ;
    wire new_AGEMA_signal_5488 ;
    wire new_AGEMA_signal_5489 ;
    wire new_AGEMA_signal_5490 ;
    wire new_AGEMA_signal_5494 ;
    wire new_AGEMA_signal_5495 ;
    wire new_AGEMA_signal_5496 ;
    wire new_AGEMA_signal_5497 ;
    wire new_AGEMA_signal_5498 ;
    wire new_AGEMA_signal_5499 ;
    wire new_AGEMA_signal_5503 ;
    wire new_AGEMA_signal_5504 ;
    wire new_AGEMA_signal_5505 ;
    wire new_AGEMA_signal_5506 ;
    wire new_AGEMA_signal_5507 ;
    wire new_AGEMA_signal_5508 ;
    wire new_AGEMA_signal_5512 ;
    wire new_AGEMA_signal_5513 ;
    wire new_AGEMA_signal_5514 ;
    wire new_AGEMA_signal_5515 ;
    wire new_AGEMA_signal_5516 ;
    wire new_AGEMA_signal_5517 ;
    wire new_AGEMA_signal_5521 ;
    wire new_AGEMA_signal_5522 ;
    wire new_AGEMA_signal_5523 ;
    wire new_AGEMA_signal_5524 ;
    wire new_AGEMA_signal_5525 ;
    wire new_AGEMA_signal_5526 ;
    wire new_AGEMA_signal_5530 ;
    wire new_AGEMA_signal_5531 ;
    wire new_AGEMA_signal_5532 ;
    wire new_AGEMA_signal_5533 ;
    wire new_AGEMA_signal_5534 ;
    wire new_AGEMA_signal_5535 ;
    wire new_AGEMA_signal_5539 ;
    wire new_AGEMA_signal_5540 ;
    wire new_AGEMA_signal_5541 ;
    wire new_AGEMA_signal_5542 ;
    wire new_AGEMA_signal_5543 ;
    wire new_AGEMA_signal_5544 ;
    wire new_AGEMA_signal_5548 ;
    wire new_AGEMA_signal_5549 ;
    wire new_AGEMA_signal_5550 ;
    wire new_AGEMA_signal_5551 ;
    wire new_AGEMA_signal_5552 ;
    wire new_AGEMA_signal_5553 ;
    wire new_AGEMA_signal_5557 ;
    wire new_AGEMA_signal_5558 ;
    wire new_AGEMA_signal_5559 ;
    wire new_AGEMA_signal_5560 ;
    wire new_AGEMA_signal_5561 ;
    wire new_AGEMA_signal_5562 ;
    wire new_AGEMA_signal_5566 ;
    wire new_AGEMA_signal_5567 ;
    wire new_AGEMA_signal_5568 ;
    wire new_AGEMA_signal_5569 ;
    wire new_AGEMA_signal_5570 ;
    wire new_AGEMA_signal_5571 ;
    wire new_AGEMA_signal_5575 ;
    wire new_AGEMA_signal_5576 ;
    wire new_AGEMA_signal_5577 ;
    wire new_AGEMA_signal_5578 ;
    wire new_AGEMA_signal_5579 ;
    wire new_AGEMA_signal_5580 ;
    wire new_AGEMA_signal_5584 ;
    wire new_AGEMA_signal_5585 ;
    wire new_AGEMA_signal_5586 ;
    wire new_AGEMA_signal_5587 ;
    wire new_AGEMA_signal_5588 ;
    wire new_AGEMA_signal_5589 ;
    wire new_AGEMA_signal_5593 ;
    wire new_AGEMA_signal_5594 ;
    wire new_AGEMA_signal_5595 ;
    wire new_AGEMA_signal_5596 ;
    wire new_AGEMA_signal_5597 ;
    wire new_AGEMA_signal_5598 ;
    wire new_AGEMA_signal_5602 ;
    wire new_AGEMA_signal_5603 ;
    wire new_AGEMA_signal_5604 ;
    wire new_AGEMA_signal_5605 ;
    wire new_AGEMA_signal_5606 ;
    wire new_AGEMA_signal_5607 ;
    wire new_AGEMA_signal_5611 ;
    wire new_AGEMA_signal_5612 ;
    wire new_AGEMA_signal_5613 ;
    wire new_AGEMA_signal_5614 ;
    wire new_AGEMA_signal_5615 ;
    wire new_AGEMA_signal_5616 ;
    wire new_AGEMA_signal_5620 ;
    wire new_AGEMA_signal_5621 ;
    wire new_AGEMA_signal_5622 ;
    wire new_AGEMA_signal_5623 ;
    wire new_AGEMA_signal_5624 ;
    wire new_AGEMA_signal_5625 ;
    wire new_AGEMA_signal_5629 ;
    wire new_AGEMA_signal_5630 ;
    wire new_AGEMA_signal_5631 ;
    wire new_AGEMA_signal_5632 ;
    wire new_AGEMA_signal_5633 ;
    wire new_AGEMA_signal_5634 ;
    wire new_AGEMA_signal_5638 ;
    wire new_AGEMA_signal_5639 ;
    wire new_AGEMA_signal_5640 ;
    wire new_AGEMA_signal_5641 ;
    wire new_AGEMA_signal_5642 ;
    wire new_AGEMA_signal_5643 ;
    wire new_AGEMA_signal_5647 ;
    wire new_AGEMA_signal_5648 ;
    wire new_AGEMA_signal_5649 ;
    wire new_AGEMA_signal_5650 ;
    wire new_AGEMA_signal_5651 ;
    wire new_AGEMA_signal_5652 ;
    wire new_AGEMA_signal_5656 ;
    wire new_AGEMA_signal_5657 ;
    wire new_AGEMA_signal_5658 ;
    wire new_AGEMA_signal_5659 ;
    wire new_AGEMA_signal_5660 ;
    wire new_AGEMA_signal_5661 ;
    wire new_AGEMA_signal_5665 ;
    wire new_AGEMA_signal_5666 ;
    wire new_AGEMA_signal_5667 ;
    wire new_AGEMA_signal_5668 ;
    wire new_AGEMA_signal_5669 ;
    wire new_AGEMA_signal_5670 ;
    wire new_AGEMA_signal_5674 ;
    wire new_AGEMA_signal_5675 ;
    wire new_AGEMA_signal_5676 ;
    wire new_AGEMA_signal_5677 ;
    wire new_AGEMA_signal_5678 ;
    wire new_AGEMA_signal_5679 ;
    wire new_AGEMA_signal_5683 ;
    wire new_AGEMA_signal_5684 ;
    wire new_AGEMA_signal_5685 ;
    wire new_AGEMA_signal_5686 ;
    wire new_AGEMA_signal_5687 ;
    wire new_AGEMA_signal_5688 ;
    wire new_AGEMA_signal_5692 ;
    wire new_AGEMA_signal_5693 ;
    wire new_AGEMA_signal_5694 ;
    wire new_AGEMA_signal_5695 ;
    wire new_AGEMA_signal_5696 ;
    wire new_AGEMA_signal_5697 ;
    wire new_AGEMA_signal_5701 ;
    wire new_AGEMA_signal_5702 ;
    wire new_AGEMA_signal_5703 ;
    wire new_AGEMA_signal_5704 ;
    wire new_AGEMA_signal_5705 ;
    wire new_AGEMA_signal_5706 ;
    wire new_AGEMA_signal_5707 ;
    wire new_AGEMA_signal_5708 ;
    wire new_AGEMA_signal_5709 ;
    wire new_AGEMA_signal_5710 ;
    wire new_AGEMA_signal_5711 ;
    wire new_AGEMA_signal_5712 ;
    wire new_AGEMA_signal_5713 ;
    wire new_AGEMA_signal_5714 ;
    wire new_AGEMA_signal_5715 ;
    wire new_AGEMA_signal_5716 ;
    wire new_AGEMA_signal_5717 ;
    wire new_AGEMA_signal_5718 ;
    wire new_AGEMA_signal_5719 ;
    wire new_AGEMA_signal_5720 ;
    wire new_AGEMA_signal_5721 ;
    wire new_AGEMA_signal_5722 ;
    wire new_AGEMA_signal_5723 ;
    wire new_AGEMA_signal_5724 ;
    wire new_AGEMA_signal_5725 ;
    wire new_AGEMA_signal_5726 ;
    wire new_AGEMA_signal_5727 ;
    wire new_AGEMA_signal_5728 ;
    wire new_AGEMA_signal_5729 ;
    wire new_AGEMA_signal_5730 ;
    wire new_AGEMA_signal_5731 ;
    wire new_AGEMA_signal_5732 ;
    wire new_AGEMA_signal_5733 ;
    wire new_AGEMA_signal_5734 ;
    wire new_AGEMA_signal_5735 ;
    wire new_AGEMA_signal_5736 ;
    wire new_AGEMA_signal_5737 ;
    wire new_AGEMA_signal_5738 ;
    wire new_AGEMA_signal_5739 ;
    wire new_AGEMA_signal_5740 ;
    wire new_AGEMA_signal_5741 ;
    wire new_AGEMA_signal_5742 ;
    wire new_AGEMA_signal_5743 ;
    wire new_AGEMA_signal_5744 ;
    wire new_AGEMA_signal_5745 ;
    wire new_AGEMA_signal_5746 ;
    wire new_AGEMA_signal_5747 ;
    wire new_AGEMA_signal_5748 ;
    wire new_AGEMA_signal_5749 ;
    wire new_AGEMA_signal_5750 ;
    wire new_AGEMA_signal_5751 ;
    wire new_AGEMA_signal_5752 ;
    wire new_AGEMA_signal_5753 ;
    wire new_AGEMA_signal_5754 ;
    wire new_AGEMA_signal_5755 ;
    wire new_AGEMA_signal_5756 ;
    wire new_AGEMA_signal_5757 ;
    wire new_AGEMA_signal_5758 ;
    wire new_AGEMA_signal_5759 ;
    wire new_AGEMA_signal_5760 ;
    wire new_AGEMA_signal_5761 ;
    wire new_AGEMA_signal_5762 ;
    wire new_AGEMA_signal_5763 ;
    wire new_AGEMA_signal_5764 ;
    wire new_AGEMA_signal_5765 ;
    wire new_AGEMA_signal_5766 ;
    wire new_AGEMA_signal_5767 ;
    wire new_AGEMA_signal_5768 ;
    wire new_AGEMA_signal_5769 ;
    wire new_AGEMA_signal_5770 ;
    wire new_AGEMA_signal_5771 ;
    wire new_AGEMA_signal_5772 ;
    wire new_AGEMA_signal_5773 ;
    wire new_AGEMA_signal_5774 ;
    wire new_AGEMA_signal_5775 ;
    wire new_AGEMA_signal_5776 ;
    wire new_AGEMA_signal_5777 ;
    wire new_AGEMA_signal_5778 ;
    wire new_AGEMA_signal_5779 ;
    wire new_AGEMA_signal_5780 ;
    wire new_AGEMA_signal_5781 ;
    wire new_AGEMA_signal_5782 ;
    wire new_AGEMA_signal_5783 ;
    wire new_AGEMA_signal_5784 ;
    wire new_AGEMA_signal_5785 ;
    wire new_AGEMA_signal_5786 ;
    wire new_AGEMA_signal_5787 ;
    wire new_AGEMA_signal_5788 ;
    wire new_AGEMA_signal_5789 ;
    wire new_AGEMA_signal_5790 ;
    wire new_AGEMA_signal_5791 ;
    wire new_AGEMA_signal_5792 ;
    wire new_AGEMA_signal_5793 ;
    wire new_AGEMA_signal_5794 ;
    wire new_AGEMA_signal_5795 ;
    wire new_AGEMA_signal_5796 ;
    wire new_AGEMA_signal_5797 ;
    wire new_AGEMA_signal_5798 ;
    wire new_AGEMA_signal_5799 ;
    wire new_AGEMA_signal_5800 ;
    wire new_AGEMA_signal_5801 ;
    wire new_AGEMA_signal_5802 ;
    wire new_AGEMA_signal_5803 ;
    wire new_AGEMA_signal_5804 ;
    wire new_AGEMA_signal_5805 ;
    wire new_AGEMA_signal_5806 ;
    wire new_AGEMA_signal_5807 ;
    wire new_AGEMA_signal_5808 ;
    wire new_AGEMA_signal_5809 ;
    wire new_AGEMA_signal_5810 ;
    wire new_AGEMA_signal_5811 ;
    wire new_AGEMA_signal_5812 ;
    wire new_AGEMA_signal_5813 ;
    wire new_AGEMA_signal_5814 ;
    wire new_AGEMA_signal_5815 ;
    wire new_AGEMA_signal_5816 ;
    wire new_AGEMA_signal_5817 ;
    wire new_AGEMA_signal_5818 ;
    wire new_AGEMA_signal_5819 ;
    wire new_AGEMA_signal_5820 ;
    wire new_AGEMA_signal_5821 ;
    wire new_AGEMA_signal_5822 ;
    wire new_AGEMA_signal_5823 ;
    wire new_AGEMA_signal_5824 ;
    wire new_AGEMA_signal_5825 ;
    wire new_AGEMA_signal_5826 ;
    wire new_AGEMA_signal_5827 ;
    wire new_AGEMA_signal_5828 ;
    wire new_AGEMA_signal_5829 ;
    wire new_AGEMA_signal_5830 ;
    wire new_AGEMA_signal_5831 ;
    wire new_AGEMA_signal_5832 ;
    wire new_AGEMA_signal_5833 ;
    wire new_AGEMA_signal_5834 ;
    wire new_AGEMA_signal_5835 ;
    wire new_AGEMA_signal_5836 ;
    wire new_AGEMA_signal_5837 ;
    wire new_AGEMA_signal_5838 ;
    wire new_AGEMA_signal_5839 ;
    wire new_AGEMA_signal_5840 ;
    wire new_AGEMA_signal_5841 ;
    wire new_AGEMA_signal_5842 ;
    wire new_AGEMA_signal_5843 ;
    wire new_AGEMA_signal_5844 ;
    wire new_AGEMA_signal_5845 ;
    wire new_AGEMA_signal_5846 ;
    wire new_AGEMA_signal_5847 ;
    wire new_AGEMA_signal_5848 ;
    wire new_AGEMA_signal_5849 ;
    wire new_AGEMA_signal_5850 ;
    wire new_AGEMA_signal_5851 ;
    wire new_AGEMA_signal_5852 ;
    wire new_AGEMA_signal_5853 ;
    wire new_AGEMA_signal_5854 ;
    wire new_AGEMA_signal_5855 ;
    wire new_AGEMA_signal_5856 ;
    wire new_AGEMA_signal_5857 ;
    wire new_AGEMA_signal_5858 ;
    wire new_AGEMA_signal_5859 ;
    wire new_AGEMA_signal_5860 ;
    wire new_AGEMA_signal_5861 ;
    wire new_AGEMA_signal_5862 ;
    wire new_AGEMA_signal_5863 ;
    wire new_AGEMA_signal_5864 ;
    wire new_AGEMA_signal_5865 ;
    wire new_AGEMA_signal_5866 ;
    wire new_AGEMA_signal_5867 ;
    wire new_AGEMA_signal_5868 ;
    wire new_AGEMA_signal_5869 ;
    wire new_AGEMA_signal_5870 ;
    wire new_AGEMA_signal_5871 ;
    wire new_AGEMA_signal_5872 ;
    wire new_AGEMA_signal_5873 ;
    wire new_AGEMA_signal_5874 ;
    wire new_AGEMA_signal_5875 ;
    wire new_AGEMA_signal_5876 ;
    wire new_AGEMA_signal_5877 ;
    wire new_AGEMA_signal_5878 ;
    wire new_AGEMA_signal_5879 ;
    wire new_AGEMA_signal_5880 ;
    wire new_AGEMA_signal_5881 ;
    wire new_AGEMA_signal_5882 ;
    wire new_AGEMA_signal_5883 ;
    wire new_AGEMA_signal_5884 ;
    wire new_AGEMA_signal_5885 ;
    wire new_AGEMA_signal_5886 ;
    wire new_AGEMA_signal_5887 ;
    wire new_AGEMA_signal_5888 ;
    wire new_AGEMA_signal_5889 ;
    wire new_AGEMA_signal_5890 ;
    wire new_AGEMA_signal_5891 ;
    wire new_AGEMA_signal_5892 ;
    wire new_AGEMA_signal_5893 ;
    wire new_AGEMA_signal_5894 ;
    wire new_AGEMA_signal_5895 ;
    wire new_AGEMA_signal_5896 ;
    wire new_AGEMA_signal_5897 ;
    wire new_AGEMA_signal_5898 ;
    wire new_AGEMA_signal_5899 ;
    wire new_AGEMA_signal_5900 ;
    wire new_AGEMA_signal_5901 ;
    wire new_AGEMA_signal_5902 ;
    wire new_AGEMA_signal_5903 ;
    wire new_AGEMA_signal_5904 ;
    wire new_AGEMA_signal_5905 ;
    wire new_AGEMA_signal_5906 ;
    wire new_AGEMA_signal_5907 ;
    wire new_AGEMA_signal_5908 ;
    wire new_AGEMA_signal_5909 ;
    wire new_AGEMA_signal_5910 ;
    wire new_AGEMA_signal_5911 ;
    wire new_AGEMA_signal_5912 ;
    wire new_AGEMA_signal_5913 ;
    wire new_AGEMA_signal_5914 ;
    wire new_AGEMA_signal_5915 ;
    wire new_AGEMA_signal_5916 ;
    wire new_AGEMA_signal_5917 ;
    wire new_AGEMA_signal_5918 ;
    wire new_AGEMA_signal_5919 ;
    wire new_AGEMA_signal_5920 ;
    wire new_AGEMA_signal_5921 ;
    wire new_AGEMA_signal_5922 ;
    wire new_AGEMA_signal_5923 ;
    wire new_AGEMA_signal_5924 ;
    wire new_AGEMA_signal_5925 ;
    wire new_AGEMA_signal_5926 ;
    wire new_AGEMA_signal_5927 ;
    wire new_AGEMA_signal_5928 ;
    wire new_AGEMA_signal_5929 ;
    wire new_AGEMA_signal_5930 ;
    wire new_AGEMA_signal_5931 ;
    wire new_AGEMA_signal_5932 ;
    wire new_AGEMA_signal_5933 ;
    wire new_AGEMA_signal_5934 ;
    wire new_AGEMA_signal_5935 ;
    wire new_AGEMA_signal_5936 ;
    wire new_AGEMA_signal_5937 ;
    wire new_AGEMA_signal_5938 ;
    wire new_AGEMA_signal_5939 ;
    wire new_AGEMA_signal_5940 ;
    wire new_AGEMA_signal_5941 ;
    wire new_AGEMA_signal_5942 ;
    wire new_AGEMA_signal_5943 ;
    wire new_AGEMA_signal_5944 ;
    wire new_AGEMA_signal_5945 ;
    wire new_AGEMA_signal_5946 ;
    wire new_AGEMA_signal_5947 ;
    wire new_AGEMA_signal_5948 ;
    wire new_AGEMA_signal_5949 ;
    wire new_AGEMA_signal_5950 ;
    wire new_AGEMA_signal_5951 ;
    wire new_AGEMA_signal_5952 ;
    wire new_AGEMA_signal_5953 ;
    wire new_AGEMA_signal_5954 ;
    wire new_AGEMA_signal_5955 ;
    wire new_AGEMA_signal_5956 ;
    wire new_AGEMA_signal_5957 ;
    wire new_AGEMA_signal_5958 ;
    wire new_AGEMA_signal_5959 ;
    wire new_AGEMA_signal_5960 ;
    wire new_AGEMA_signal_5961 ;
    wire new_AGEMA_signal_5962 ;
    wire new_AGEMA_signal_5963 ;
    wire new_AGEMA_signal_5964 ;
    wire new_AGEMA_signal_5965 ;
    wire new_AGEMA_signal_5966 ;
    wire new_AGEMA_signal_5967 ;
    wire new_AGEMA_signal_5968 ;
    wire new_AGEMA_signal_5969 ;
    wire new_AGEMA_signal_5970 ;
    wire new_AGEMA_signal_5971 ;
    wire new_AGEMA_signal_5972 ;
    wire new_AGEMA_signal_5973 ;
    wire new_AGEMA_signal_5974 ;
    wire new_AGEMA_signal_5975 ;
    wire new_AGEMA_signal_5976 ;
    wire new_AGEMA_signal_5977 ;
    wire new_AGEMA_signal_5978 ;
    wire new_AGEMA_signal_5979 ;
    wire new_AGEMA_signal_5980 ;
    wire new_AGEMA_signal_5981 ;
    wire new_AGEMA_signal_5982 ;
    wire new_AGEMA_signal_5983 ;
    wire new_AGEMA_signal_5984 ;
    wire new_AGEMA_signal_5985 ;
    wire new_AGEMA_signal_5986 ;
    wire new_AGEMA_signal_5987 ;
    wire new_AGEMA_signal_5988 ;
    wire new_AGEMA_signal_5989 ;
    wire new_AGEMA_signal_5990 ;
    wire new_AGEMA_signal_5991 ;
    wire new_AGEMA_signal_5992 ;
    wire new_AGEMA_signal_5993 ;
    wire new_AGEMA_signal_5994 ;
    wire new_AGEMA_signal_5995 ;
    wire new_AGEMA_signal_5996 ;
    wire new_AGEMA_signal_5997 ;
    wire new_AGEMA_signal_5998 ;
    wire new_AGEMA_signal_5999 ;
    wire new_AGEMA_signal_6000 ;
    wire new_AGEMA_signal_6001 ;
    wire new_AGEMA_signal_6002 ;
    wire new_AGEMA_signal_6003 ;
    wire new_AGEMA_signal_6004 ;
    wire new_AGEMA_signal_6005 ;
    wire new_AGEMA_signal_6006 ;
    wire new_AGEMA_signal_6007 ;
    wire new_AGEMA_signal_6008 ;
    wire new_AGEMA_signal_6009 ;
    wire new_AGEMA_signal_6010 ;
    wire new_AGEMA_signal_6011 ;
    wire new_AGEMA_signal_6012 ;
    wire new_AGEMA_signal_6013 ;
    wire new_AGEMA_signal_6014 ;
    wire new_AGEMA_signal_6015 ;
    wire new_AGEMA_signal_6016 ;
    wire new_AGEMA_signal_6017 ;
    wire new_AGEMA_signal_6018 ;
    wire new_AGEMA_signal_6019 ;
    wire new_AGEMA_signal_6020 ;
    wire new_AGEMA_signal_6021 ;
    wire new_AGEMA_signal_6022 ;
    wire new_AGEMA_signal_6023 ;
    wire new_AGEMA_signal_6024 ;
    wire new_AGEMA_signal_6025 ;
    wire new_AGEMA_signal_6026 ;
    wire new_AGEMA_signal_6027 ;
    wire new_AGEMA_signal_6028 ;
    wire new_AGEMA_signal_6029 ;
    wire new_AGEMA_signal_6030 ;
    wire new_AGEMA_signal_6031 ;
    wire new_AGEMA_signal_6032 ;
    wire new_AGEMA_signal_6033 ;
    wire new_AGEMA_signal_6034 ;
    wire new_AGEMA_signal_6035 ;
    wire new_AGEMA_signal_6036 ;
    wire new_AGEMA_signal_6037 ;
    wire new_AGEMA_signal_6038 ;
    wire new_AGEMA_signal_6039 ;
    wire new_AGEMA_signal_6040 ;
    wire new_AGEMA_signal_6041 ;
    wire new_AGEMA_signal_6042 ;
    wire new_AGEMA_signal_6043 ;
    wire new_AGEMA_signal_6044 ;
    wire new_AGEMA_signal_6045 ;
    wire new_AGEMA_signal_6046 ;
    wire new_AGEMA_signal_6047 ;
    wire new_AGEMA_signal_6048 ;
    wire new_AGEMA_signal_6049 ;
    wire new_AGEMA_signal_6050 ;
    wire new_AGEMA_signal_6051 ;
    wire new_AGEMA_signal_6052 ;
    wire new_AGEMA_signal_6053 ;
    wire new_AGEMA_signal_6054 ;
    wire new_AGEMA_signal_6055 ;
    wire new_AGEMA_signal_6056 ;
    wire new_AGEMA_signal_6057 ;
    wire new_AGEMA_signal_6058 ;
    wire new_AGEMA_signal_6059 ;
    wire new_AGEMA_signal_6060 ;
    wire new_AGEMA_signal_6061 ;
    wire new_AGEMA_signal_6062 ;
    wire new_AGEMA_signal_6063 ;
    wire new_AGEMA_signal_6064 ;
    wire new_AGEMA_signal_6065 ;
    wire new_AGEMA_signal_6066 ;
    wire new_AGEMA_signal_6067 ;
    wire new_AGEMA_signal_6068 ;
    wire new_AGEMA_signal_6069 ;
    wire new_AGEMA_signal_6070 ;
    wire new_AGEMA_signal_6071 ;
    wire new_AGEMA_signal_6072 ;
    wire new_AGEMA_signal_6073 ;
    wire new_AGEMA_signal_6074 ;
    wire new_AGEMA_signal_6075 ;
    wire new_AGEMA_signal_6076 ;
    wire new_AGEMA_signal_6077 ;
    wire new_AGEMA_signal_6078 ;
    wire new_AGEMA_signal_6079 ;
    wire new_AGEMA_signal_6080 ;
    wire new_AGEMA_signal_6081 ;
    wire new_AGEMA_signal_6082 ;
    wire new_AGEMA_signal_6083 ;
    wire new_AGEMA_signal_6084 ;
    wire new_AGEMA_signal_6085 ;
    wire new_AGEMA_signal_6086 ;
    wire new_AGEMA_signal_6087 ;
    wire new_AGEMA_signal_6088 ;
    wire new_AGEMA_signal_6089 ;
    wire new_AGEMA_signal_6090 ;
    wire new_AGEMA_signal_6091 ;
    wire new_AGEMA_signal_6092 ;
    wire new_AGEMA_signal_6093 ;
    wire new_AGEMA_signal_6094 ;
    wire new_AGEMA_signal_6095 ;
    wire new_AGEMA_signal_6096 ;
    wire new_AGEMA_signal_6097 ;
    wire new_AGEMA_signal_6098 ;
    wire new_AGEMA_signal_6099 ;
    wire new_AGEMA_signal_6100 ;
    wire new_AGEMA_signal_6101 ;
    wire new_AGEMA_signal_6102 ;
    wire new_AGEMA_signal_6103 ;
    wire new_AGEMA_signal_6104 ;
    wire new_AGEMA_signal_6105 ;
    wire new_AGEMA_signal_6106 ;
    wire new_AGEMA_signal_6107 ;
    wire new_AGEMA_signal_6108 ;
    wire new_AGEMA_signal_6109 ;
    wire new_AGEMA_signal_6110 ;
    wire new_AGEMA_signal_6111 ;
    wire new_AGEMA_signal_6112 ;
    wire new_AGEMA_signal_6113 ;
    wire new_AGEMA_signal_6114 ;
    wire new_AGEMA_signal_6115 ;
    wire new_AGEMA_signal_6116 ;
    wire new_AGEMA_signal_6117 ;
    wire new_AGEMA_signal_6118 ;
    wire new_AGEMA_signal_6119 ;
    wire new_AGEMA_signal_6120 ;
    wire new_AGEMA_signal_6121 ;
    wire new_AGEMA_signal_6122 ;
    wire new_AGEMA_signal_6123 ;
    wire new_AGEMA_signal_6124 ;
    wire new_AGEMA_signal_6125 ;
    wire new_AGEMA_signal_6126 ;
    wire new_AGEMA_signal_6127 ;
    wire new_AGEMA_signal_6128 ;
    wire new_AGEMA_signal_6129 ;
    wire new_AGEMA_signal_6130 ;
    wire new_AGEMA_signal_6131 ;
    wire new_AGEMA_signal_6132 ;
    wire new_AGEMA_signal_6133 ;
    wire new_AGEMA_signal_6134 ;
    wire new_AGEMA_signal_6135 ;
    wire new_AGEMA_signal_6136 ;
    wire new_AGEMA_signal_6137 ;
    wire new_AGEMA_signal_6138 ;
    wire new_AGEMA_signal_6139 ;
    wire new_AGEMA_signal_6140 ;
    wire new_AGEMA_signal_6141 ;
    wire new_AGEMA_signal_6142 ;
    wire new_AGEMA_signal_6143 ;
    wire new_AGEMA_signal_6144 ;
    wire new_AGEMA_signal_6145 ;
    wire new_AGEMA_signal_6146 ;
    wire new_AGEMA_signal_6147 ;
    wire new_AGEMA_signal_6148 ;
    wire new_AGEMA_signal_6149 ;
    wire new_AGEMA_signal_6150 ;
    wire new_AGEMA_signal_6151 ;
    wire new_AGEMA_signal_6152 ;
    wire new_AGEMA_signal_6153 ;
    wire new_AGEMA_signal_6154 ;
    wire new_AGEMA_signal_6155 ;
    wire new_AGEMA_signal_6156 ;
    wire new_AGEMA_signal_6157 ;
    wire new_AGEMA_signal_6158 ;
    wire new_AGEMA_signal_6159 ;
    wire new_AGEMA_signal_6160 ;
    wire new_AGEMA_signal_6161 ;
    wire new_AGEMA_signal_6162 ;
    wire new_AGEMA_signal_6163 ;
    wire new_AGEMA_signal_6164 ;
    wire new_AGEMA_signal_6165 ;
    wire new_AGEMA_signal_6166 ;
    wire new_AGEMA_signal_6167 ;
    wire new_AGEMA_signal_6168 ;
    wire new_AGEMA_signal_6169 ;
    wire new_AGEMA_signal_6170 ;
    wire new_AGEMA_signal_6171 ;
    wire new_AGEMA_signal_6172 ;
    wire new_AGEMA_signal_6173 ;
    wire new_AGEMA_signal_6174 ;
    wire new_AGEMA_signal_6175 ;
    wire new_AGEMA_signal_6176 ;
    wire new_AGEMA_signal_6177 ;
    wire new_AGEMA_signal_6178 ;
    wire new_AGEMA_signal_6179 ;
    wire new_AGEMA_signal_6180 ;
    wire new_AGEMA_signal_6181 ;
    wire new_AGEMA_signal_6182 ;
    wire new_AGEMA_signal_6183 ;
    wire new_AGEMA_signal_6184 ;
    wire new_AGEMA_signal_6185 ;
    wire new_AGEMA_signal_6186 ;
    wire new_AGEMA_signal_6187 ;
    wire new_AGEMA_signal_6188 ;
    wire new_AGEMA_signal_6189 ;
    wire new_AGEMA_signal_6190 ;
    wire new_AGEMA_signal_6191 ;
    wire new_AGEMA_signal_6192 ;
    wire new_AGEMA_signal_6193 ;
    wire new_AGEMA_signal_6194 ;
    wire new_AGEMA_signal_6195 ;
    wire new_AGEMA_signal_6196 ;
    wire new_AGEMA_signal_6197 ;
    wire new_AGEMA_signal_6198 ;
    wire new_AGEMA_signal_6199 ;
    wire new_AGEMA_signal_6200 ;
    wire new_AGEMA_signal_6201 ;
    wire new_AGEMA_signal_6202 ;
    wire new_AGEMA_signal_6203 ;
    wire new_AGEMA_signal_6204 ;
    wire new_AGEMA_signal_6205 ;
    wire new_AGEMA_signal_6206 ;
    wire new_AGEMA_signal_6207 ;
    wire new_AGEMA_signal_6208 ;
    wire new_AGEMA_signal_6209 ;
    wire new_AGEMA_signal_6210 ;
    wire new_AGEMA_signal_6211 ;
    wire new_AGEMA_signal_6212 ;
    wire new_AGEMA_signal_6213 ;
    wire new_AGEMA_signal_6214 ;
    wire new_AGEMA_signal_6215 ;
    wire new_AGEMA_signal_6216 ;
    wire new_AGEMA_signal_6217 ;
    wire new_AGEMA_signal_6218 ;
    wire new_AGEMA_signal_6219 ;
    wire new_AGEMA_signal_6220 ;
    wire new_AGEMA_signal_6221 ;
    wire new_AGEMA_signal_6222 ;
    wire new_AGEMA_signal_6223 ;
    wire new_AGEMA_signal_6224 ;
    wire new_AGEMA_signal_6225 ;
    wire new_AGEMA_signal_6226 ;
    wire new_AGEMA_signal_6227 ;
    wire new_AGEMA_signal_6228 ;
    wire new_AGEMA_signal_6229 ;
    wire new_AGEMA_signal_6230 ;
    wire new_AGEMA_signal_6231 ;
    wire new_AGEMA_signal_6232 ;
    wire new_AGEMA_signal_6233 ;
    wire new_AGEMA_signal_6234 ;
    wire new_AGEMA_signal_6235 ;
    wire new_AGEMA_signal_6236 ;
    wire new_AGEMA_signal_6237 ;
    wire new_AGEMA_signal_6238 ;
    wire new_AGEMA_signal_6239 ;
    wire new_AGEMA_signal_6240 ;
    wire new_AGEMA_signal_6241 ;
    wire new_AGEMA_signal_6242 ;
    wire new_AGEMA_signal_6243 ;
    wire new_AGEMA_signal_6244 ;
    wire new_AGEMA_signal_6245 ;
    wire new_AGEMA_signal_6246 ;
    wire new_AGEMA_signal_6247 ;
    wire new_AGEMA_signal_6248 ;
    wire new_AGEMA_signal_6249 ;
    wire new_AGEMA_signal_6250 ;
    wire new_AGEMA_signal_6251 ;
    wire new_AGEMA_signal_6252 ;
    wire new_AGEMA_signal_6253 ;
    wire new_AGEMA_signal_6254 ;
    wire new_AGEMA_signal_6255 ;
    wire new_AGEMA_signal_6256 ;
    wire new_AGEMA_signal_6257 ;
    wire new_AGEMA_signal_6258 ;
    wire new_AGEMA_signal_6259 ;
    wire new_AGEMA_signal_6260 ;
    wire new_AGEMA_signal_6261 ;
    wire new_AGEMA_signal_6262 ;
    wire new_AGEMA_signal_6263 ;
    wire new_AGEMA_signal_6264 ;
    wire new_AGEMA_signal_6265 ;
    wire new_AGEMA_signal_6266 ;
    wire new_AGEMA_signal_6267 ;
    wire new_AGEMA_signal_6268 ;
    wire new_AGEMA_signal_6269 ;
    wire new_AGEMA_signal_6270 ;
    wire new_AGEMA_signal_6271 ;
    wire new_AGEMA_signal_6272 ;
    wire new_AGEMA_signal_6273 ;
    wire new_AGEMA_signal_6274 ;
    wire new_AGEMA_signal_6275 ;
    wire new_AGEMA_signal_6276 ;
    wire new_AGEMA_signal_6277 ;
    wire new_AGEMA_signal_6278 ;
    wire new_AGEMA_signal_6279 ;
    wire new_AGEMA_signal_6280 ;
    wire new_AGEMA_signal_6281 ;
    wire new_AGEMA_signal_6282 ;
    wire new_AGEMA_signal_6283 ;
    wire new_AGEMA_signal_6284 ;
    wire new_AGEMA_signal_6285 ;
    wire new_AGEMA_signal_6286 ;
    wire new_AGEMA_signal_6287 ;
    wire new_AGEMA_signal_6288 ;
    wire new_AGEMA_signal_6289 ;
    wire new_AGEMA_signal_6290 ;
    wire new_AGEMA_signal_6291 ;
    wire new_AGEMA_signal_6292 ;
    wire new_AGEMA_signal_6293 ;
    wire new_AGEMA_signal_6294 ;
    wire new_AGEMA_signal_6295 ;
    wire new_AGEMA_signal_6296 ;
    wire new_AGEMA_signal_6297 ;
    wire new_AGEMA_signal_6298 ;
    wire new_AGEMA_signal_6299 ;
    wire new_AGEMA_signal_6300 ;
    wire new_AGEMA_signal_6301 ;
    wire new_AGEMA_signal_6302 ;
    wire new_AGEMA_signal_6303 ;
    wire new_AGEMA_signal_6304 ;
    wire new_AGEMA_signal_6305 ;
    wire new_AGEMA_signal_6306 ;
    wire new_AGEMA_signal_6307 ;
    wire new_AGEMA_signal_6308 ;
    wire new_AGEMA_signal_6309 ;
    wire new_AGEMA_signal_6310 ;
    wire new_AGEMA_signal_6311 ;
    wire new_AGEMA_signal_6312 ;
    wire new_AGEMA_signal_6313 ;
    wire new_AGEMA_signal_6314 ;
    wire new_AGEMA_signal_6315 ;
    wire new_AGEMA_signal_6316 ;
    wire new_AGEMA_signal_6317 ;
    wire new_AGEMA_signal_6318 ;
    wire new_AGEMA_signal_6319 ;
    wire new_AGEMA_signal_6320 ;
    wire new_AGEMA_signal_6321 ;
    wire new_AGEMA_signal_6322 ;
    wire new_AGEMA_signal_6323 ;
    wire new_AGEMA_signal_6324 ;
    wire new_AGEMA_signal_6325 ;
    wire new_AGEMA_signal_6326 ;
    wire new_AGEMA_signal_6327 ;
    wire new_AGEMA_signal_6328 ;
    wire new_AGEMA_signal_6329 ;
    wire new_AGEMA_signal_6330 ;
    wire new_AGEMA_signal_6331 ;
    wire new_AGEMA_signal_6332 ;
    wire new_AGEMA_signal_6333 ;
    wire new_AGEMA_signal_6334 ;
    wire new_AGEMA_signal_6335 ;
    wire new_AGEMA_signal_6336 ;
    wire new_AGEMA_signal_6337 ;
    wire new_AGEMA_signal_6338 ;
    wire new_AGEMA_signal_6339 ;
    wire new_AGEMA_signal_6340 ;
    wire new_AGEMA_signal_6341 ;
    wire new_AGEMA_signal_6342 ;
    wire new_AGEMA_signal_6343 ;
    wire new_AGEMA_signal_6344 ;
    wire new_AGEMA_signal_6345 ;
    wire new_AGEMA_signal_6346 ;
    wire new_AGEMA_signal_6347 ;
    wire new_AGEMA_signal_6348 ;
    wire new_AGEMA_signal_6349 ;
    wire new_AGEMA_signal_6350 ;
    wire new_AGEMA_signal_6351 ;
    wire new_AGEMA_signal_6352 ;
    wire new_AGEMA_signal_6353 ;
    wire new_AGEMA_signal_6354 ;
    wire new_AGEMA_signal_6355 ;
    wire new_AGEMA_signal_6356 ;
    wire new_AGEMA_signal_6357 ;
    wire new_AGEMA_signal_6358 ;
    wire new_AGEMA_signal_6359 ;
    wire new_AGEMA_signal_6360 ;
    wire new_AGEMA_signal_6361 ;
    wire new_AGEMA_signal_6362 ;
    wire new_AGEMA_signal_6363 ;
    wire new_AGEMA_signal_6364 ;
    wire new_AGEMA_signal_6365 ;
    wire new_AGEMA_signal_6366 ;
    wire new_AGEMA_signal_6367 ;
    wire new_AGEMA_signal_6368 ;
    wire new_AGEMA_signal_6369 ;
    wire new_AGEMA_signal_6370 ;
    wire new_AGEMA_signal_6371 ;
    wire new_AGEMA_signal_6372 ;
    wire new_AGEMA_signal_6373 ;
    wire new_AGEMA_signal_6374 ;
    wire new_AGEMA_signal_6375 ;
    wire new_AGEMA_signal_6376 ;
    wire new_AGEMA_signal_6377 ;
    wire new_AGEMA_signal_6378 ;
    wire new_AGEMA_signal_6379 ;
    wire new_AGEMA_signal_6380 ;
    wire new_AGEMA_signal_6381 ;
    wire new_AGEMA_signal_6382 ;
    wire new_AGEMA_signal_6383 ;
    wire new_AGEMA_signal_6384 ;
    wire new_AGEMA_signal_6385 ;
    wire new_AGEMA_signal_6386 ;
    wire new_AGEMA_signal_6387 ;
    wire new_AGEMA_signal_6388 ;
    wire new_AGEMA_signal_6389 ;
    wire new_AGEMA_signal_6390 ;
    wire new_AGEMA_signal_6391 ;
    wire new_AGEMA_signal_6392 ;
    wire new_AGEMA_signal_6393 ;
    wire new_AGEMA_signal_6394 ;
    wire new_AGEMA_signal_6395 ;
    wire new_AGEMA_signal_6396 ;
    wire new_AGEMA_signal_6397 ;
    wire new_AGEMA_signal_6398 ;
    wire new_AGEMA_signal_6399 ;
    wire new_AGEMA_signal_6400 ;
    wire new_AGEMA_signal_6401 ;
    wire new_AGEMA_signal_6402 ;
    wire new_AGEMA_signal_6403 ;
    wire new_AGEMA_signal_6404 ;
    wire new_AGEMA_signal_6405 ;
    wire new_AGEMA_signal_6406 ;
    wire new_AGEMA_signal_6407 ;
    wire new_AGEMA_signal_6408 ;
    wire new_AGEMA_signal_6409 ;
    wire new_AGEMA_signal_6410 ;
    wire new_AGEMA_signal_6411 ;
    wire new_AGEMA_signal_6412 ;
    wire new_AGEMA_signal_6413 ;
    wire new_AGEMA_signal_6414 ;
    wire new_AGEMA_signal_6415 ;
    wire new_AGEMA_signal_6416 ;
    wire new_AGEMA_signal_6417 ;
    wire new_AGEMA_signal_6418 ;
    wire new_AGEMA_signal_6419 ;
    wire new_AGEMA_signal_6420 ;
    wire new_AGEMA_signal_6421 ;
    wire new_AGEMA_signal_6422 ;
    wire new_AGEMA_signal_6423 ;
    wire new_AGEMA_signal_6424 ;
    wire new_AGEMA_signal_6425 ;
    wire new_AGEMA_signal_6426 ;
    wire new_AGEMA_signal_6427 ;
    wire new_AGEMA_signal_6428 ;
    wire new_AGEMA_signal_6429 ;
    wire new_AGEMA_signal_6430 ;
    wire new_AGEMA_signal_6431 ;
    wire new_AGEMA_signal_6432 ;
    wire new_AGEMA_signal_6433 ;
    wire new_AGEMA_signal_6434 ;
    wire new_AGEMA_signal_6435 ;
    wire new_AGEMA_signal_6436 ;
    wire new_AGEMA_signal_6437 ;
    wire new_AGEMA_signal_6438 ;
    wire new_AGEMA_signal_6439 ;
    wire new_AGEMA_signal_6440 ;
    wire new_AGEMA_signal_6441 ;
    wire new_AGEMA_signal_6442 ;
    wire new_AGEMA_signal_6443 ;
    wire new_AGEMA_signal_6444 ;
    wire new_AGEMA_signal_6445 ;
    wire new_AGEMA_signal_6446 ;
    wire new_AGEMA_signal_6447 ;
    wire new_AGEMA_signal_6448 ;
    wire new_AGEMA_signal_6449 ;
    wire new_AGEMA_signal_6450 ;
    wire new_AGEMA_signal_6451 ;
    wire new_AGEMA_signal_6452 ;
    wire new_AGEMA_signal_6453 ;
    wire new_AGEMA_signal_6454 ;
    wire new_AGEMA_signal_6455 ;
    wire new_AGEMA_signal_6456 ;
    wire new_AGEMA_signal_6457 ;
    wire new_AGEMA_signal_6458 ;
    wire new_AGEMA_signal_6459 ;
    wire new_AGEMA_signal_6460 ;
    wire new_AGEMA_signal_6461 ;
    wire new_AGEMA_signal_6462 ;
    wire new_AGEMA_signal_6463 ;
    wire new_AGEMA_signal_6464 ;
    wire new_AGEMA_signal_6465 ;
    wire new_AGEMA_signal_6466 ;
    wire new_AGEMA_signal_6467 ;
    wire new_AGEMA_signal_6468 ;
    wire new_AGEMA_signal_6469 ;
    wire new_AGEMA_signal_6470 ;
    wire new_AGEMA_signal_6471 ;
    wire new_AGEMA_signal_6472 ;
    wire new_AGEMA_signal_6473 ;
    wire new_AGEMA_signal_6474 ;
    wire new_AGEMA_signal_6475 ;
    wire new_AGEMA_signal_6476 ;
    wire new_AGEMA_signal_6477 ;
    wire new_AGEMA_signal_6478 ;
    wire new_AGEMA_signal_6479 ;
    wire new_AGEMA_signal_6480 ;
    wire new_AGEMA_signal_6481 ;
    wire new_AGEMA_signal_6482 ;
    wire new_AGEMA_signal_6483 ;
    wire new_AGEMA_signal_6484 ;
    wire new_AGEMA_signal_6485 ;
    wire new_AGEMA_signal_6486 ;
    wire new_AGEMA_signal_6487 ;
    wire new_AGEMA_signal_6488 ;
    wire new_AGEMA_signal_6489 ;
    wire new_AGEMA_signal_6490 ;
    wire new_AGEMA_signal_6491 ;
    wire new_AGEMA_signal_6492 ;
    wire new_AGEMA_signal_6493 ;
    wire new_AGEMA_signal_6494 ;
    wire new_AGEMA_signal_6495 ;
    wire new_AGEMA_signal_6496 ;
    wire new_AGEMA_signal_6497 ;
    wire new_AGEMA_signal_6498 ;
    wire new_AGEMA_signal_6499 ;
    wire new_AGEMA_signal_6500 ;
    wire new_AGEMA_signal_6501 ;
    wire new_AGEMA_signal_6502 ;
    wire new_AGEMA_signal_6503 ;
    wire new_AGEMA_signal_6504 ;
    wire new_AGEMA_signal_6505 ;
    wire new_AGEMA_signal_6506 ;
    wire new_AGEMA_signal_6507 ;
    wire new_AGEMA_signal_6508 ;
    wire new_AGEMA_signal_6509 ;
    wire new_AGEMA_signal_6510 ;
    wire new_AGEMA_signal_6511 ;
    wire new_AGEMA_signal_6512 ;
    wire new_AGEMA_signal_6513 ;
    wire new_AGEMA_signal_6514 ;
    wire new_AGEMA_signal_6515 ;
    wire new_AGEMA_signal_6516 ;
    wire new_AGEMA_signal_6517 ;
    wire new_AGEMA_signal_6518 ;
    wire new_AGEMA_signal_6519 ;
    wire new_AGEMA_signal_6520 ;
    wire new_AGEMA_signal_6521 ;
    wire new_AGEMA_signal_6522 ;
    wire new_AGEMA_signal_6523 ;
    wire new_AGEMA_signal_6524 ;
    wire new_AGEMA_signal_6525 ;
    wire new_AGEMA_signal_6526 ;
    wire new_AGEMA_signal_6527 ;
    wire new_AGEMA_signal_6528 ;
    wire new_AGEMA_signal_6529 ;
    wire new_AGEMA_signal_6530 ;
    wire new_AGEMA_signal_6531 ;
    wire new_AGEMA_signal_6532 ;
    wire new_AGEMA_signal_6533 ;
    wire new_AGEMA_signal_6534 ;
    wire new_AGEMA_signal_6535 ;
    wire new_AGEMA_signal_6536 ;
    wire new_AGEMA_signal_6537 ;
    wire new_AGEMA_signal_6538 ;
    wire new_AGEMA_signal_6539 ;
    wire new_AGEMA_signal_6540 ;
    wire new_AGEMA_signal_6541 ;
    wire new_AGEMA_signal_6542 ;
    wire new_AGEMA_signal_6543 ;
    wire new_AGEMA_signal_6544 ;
    wire new_AGEMA_signal_6545 ;
    wire new_AGEMA_signal_6546 ;
    wire new_AGEMA_signal_6547 ;
    wire new_AGEMA_signal_6548 ;
    wire new_AGEMA_signal_6549 ;
    wire new_AGEMA_signal_6550 ;
    wire new_AGEMA_signal_6551 ;
    wire new_AGEMA_signal_6552 ;
    wire new_AGEMA_signal_6553 ;
    wire new_AGEMA_signal_6554 ;
    wire new_AGEMA_signal_6555 ;
    wire new_AGEMA_signal_6556 ;
    wire new_AGEMA_signal_6557 ;
    wire new_AGEMA_signal_6558 ;
    wire new_AGEMA_signal_6559 ;
    wire new_AGEMA_signal_6560 ;
    wire new_AGEMA_signal_6561 ;
    wire new_AGEMA_signal_6562 ;
    wire new_AGEMA_signal_6563 ;
    wire new_AGEMA_signal_6564 ;
    wire new_AGEMA_signal_6565 ;
    wire new_AGEMA_signal_6566 ;
    wire new_AGEMA_signal_6567 ;
    wire new_AGEMA_signal_6568 ;
    wire new_AGEMA_signal_6569 ;
    wire new_AGEMA_signal_6570 ;
    wire new_AGEMA_signal_6571 ;
    wire new_AGEMA_signal_6572 ;
    wire new_AGEMA_signal_6573 ;
    wire new_AGEMA_signal_6574 ;
    wire new_AGEMA_signal_6575 ;
    wire new_AGEMA_signal_6576 ;
    wire new_AGEMA_signal_6577 ;
    wire new_AGEMA_signal_6578 ;
    wire new_AGEMA_signal_6579 ;
    wire new_AGEMA_signal_6580 ;
    wire new_AGEMA_signal_6581 ;
    wire new_AGEMA_signal_6582 ;
    wire new_AGEMA_signal_6583 ;
    wire new_AGEMA_signal_6584 ;
    wire new_AGEMA_signal_6585 ;
    wire new_AGEMA_signal_6586 ;
    wire new_AGEMA_signal_6587 ;
    wire new_AGEMA_signal_6588 ;
    wire new_AGEMA_signal_6589 ;
    wire new_AGEMA_signal_6590 ;
    wire new_AGEMA_signal_6591 ;
    wire new_AGEMA_signal_6592 ;
    wire new_AGEMA_signal_6593 ;
    wire new_AGEMA_signal_6594 ;
    wire new_AGEMA_signal_6595 ;
    wire new_AGEMA_signal_6596 ;
    wire new_AGEMA_signal_6597 ;
    wire new_AGEMA_signal_6598 ;
    wire new_AGEMA_signal_6599 ;
    wire new_AGEMA_signal_6600 ;
    wire new_AGEMA_signal_6601 ;
    wire new_AGEMA_signal_6602 ;
    wire new_AGEMA_signal_6603 ;
    wire new_AGEMA_signal_6604 ;
    wire new_AGEMA_signal_6605 ;
    wire new_AGEMA_signal_6606 ;
    wire new_AGEMA_signal_6607 ;
    wire new_AGEMA_signal_6608 ;
    wire new_AGEMA_signal_6609 ;
    wire new_AGEMA_signal_6610 ;
    wire new_AGEMA_signal_6611 ;
    wire new_AGEMA_signal_6612 ;
    wire new_AGEMA_signal_6613 ;
    wire new_AGEMA_signal_6614 ;
    wire new_AGEMA_signal_6615 ;
    wire new_AGEMA_signal_6616 ;
    wire new_AGEMA_signal_6617 ;
    wire new_AGEMA_signal_6618 ;
    wire new_AGEMA_signal_6619 ;
    wire new_AGEMA_signal_6620 ;
    wire new_AGEMA_signal_6621 ;
    wire new_AGEMA_signal_6622 ;
    wire new_AGEMA_signal_6623 ;
    wire new_AGEMA_signal_6624 ;
    wire new_AGEMA_signal_6625 ;
    wire new_AGEMA_signal_6626 ;
    wire new_AGEMA_signal_6627 ;
    wire new_AGEMA_signal_6628 ;
    wire new_AGEMA_signal_6629 ;
    wire new_AGEMA_signal_6630 ;
    wire new_AGEMA_signal_6631 ;
    wire new_AGEMA_signal_6632 ;
    wire new_AGEMA_signal_6633 ;
    wire new_AGEMA_signal_6634 ;
    wire new_AGEMA_signal_6635 ;
    wire new_AGEMA_signal_6636 ;
    wire new_AGEMA_signal_6637 ;
    wire new_AGEMA_signal_6638 ;
    wire new_AGEMA_signal_6639 ;
    wire new_AGEMA_signal_6640 ;
    wire new_AGEMA_signal_6641 ;
    wire new_AGEMA_signal_6642 ;
    wire new_AGEMA_signal_6643 ;
    wire new_AGEMA_signal_6644 ;
    wire new_AGEMA_signal_6645 ;
    wire new_AGEMA_signal_6646 ;
    wire new_AGEMA_signal_6647 ;
    wire new_AGEMA_signal_6648 ;
    wire new_AGEMA_signal_6649 ;
    wire new_AGEMA_signal_6650 ;
    wire new_AGEMA_signal_6651 ;
    wire new_AGEMA_signal_6652 ;
    wire new_AGEMA_signal_6653 ;
    wire new_AGEMA_signal_6654 ;
    wire new_AGEMA_signal_6655 ;
    wire new_AGEMA_signal_6656 ;
    wire new_AGEMA_signal_6657 ;
    wire new_AGEMA_signal_6658 ;
    wire new_AGEMA_signal_6659 ;
    wire new_AGEMA_signal_6660 ;
    wire new_AGEMA_signal_6661 ;
    wire new_AGEMA_signal_6662 ;
    wire new_AGEMA_signal_6663 ;
    wire new_AGEMA_signal_6664 ;
    wire new_AGEMA_signal_6665 ;
    wire new_AGEMA_signal_6666 ;
    wire new_AGEMA_signal_6667 ;
    wire new_AGEMA_signal_6668 ;
    wire new_AGEMA_signal_6669 ;
    wire new_AGEMA_signal_6670 ;
    wire new_AGEMA_signal_6671 ;
    wire new_AGEMA_signal_6672 ;
    wire new_AGEMA_signal_6673 ;
    wire new_AGEMA_signal_6674 ;
    wire new_AGEMA_signal_6675 ;
    wire new_AGEMA_signal_6676 ;
    wire new_AGEMA_signal_6677 ;
    wire new_AGEMA_signal_6678 ;
    wire new_AGEMA_signal_6679 ;
    wire new_AGEMA_signal_6680 ;
    wire new_AGEMA_signal_6681 ;
    wire new_AGEMA_signal_6682 ;
    wire new_AGEMA_signal_6683 ;
    wire new_AGEMA_signal_6684 ;
    wire new_AGEMA_signal_6685 ;
    wire new_AGEMA_signal_6686 ;
    wire new_AGEMA_signal_6687 ;
    wire new_AGEMA_signal_6688 ;
    wire new_AGEMA_signal_6689 ;
    wire new_AGEMA_signal_6690 ;
    wire new_AGEMA_signal_6691 ;
    wire new_AGEMA_signal_6692 ;
    wire new_AGEMA_signal_6693 ;
    wire new_AGEMA_signal_6694 ;
    wire new_AGEMA_signal_6695 ;
    wire new_AGEMA_signal_6696 ;
    wire new_AGEMA_signal_6697 ;
    wire new_AGEMA_signal_6698 ;
    wire new_AGEMA_signal_6699 ;
    wire new_AGEMA_signal_6700 ;
    wire new_AGEMA_signal_6701 ;
    wire new_AGEMA_signal_6702 ;
    wire new_AGEMA_signal_6703 ;
    wire new_AGEMA_signal_6704 ;
    wire new_AGEMA_signal_6705 ;
    wire new_AGEMA_signal_6706 ;
    wire new_AGEMA_signal_6707 ;
    wire new_AGEMA_signal_6708 ;
    wire new_AGEMA_signal_6709 ;
    wire new_AGEMA_signal_6710 ;
    wire new_AGEMA_signal_6711 ;
    wire new_AGEMA_signal_6712 ;
    wire new_AGEMA_signal_6713 ;
    wire new_AGEMA_signal_6714 ;
    wire new_AGEMA_signal_6715 ;
    wire new_AGEMA_signal_6716 ;
    wire new_AGEMA_signal_6717 ;
    wire new_AGEMA_signal_6718 ;
    wire new_AGEMA_signal_6719 ;
    wire new_AGEMA_signal_6720 ;
    wire new_AGEMA_signal_6721 ;
    wire new_AGEMA_signal_6722 ;
    wire new_AGEMA_signal_6723 ;
    wire new_AGEMA_signal_6724 ;
    wire new_AGEMA_signal_6725 ;
    wire new_AGEMA_signal_6726 ;
    wire new_AGEMA_signal_6727 ;
    wire new_AGEMA_signal_6728 ;
    wire new_AGEMA_signal_6729 ;
    wire new_AGEMA_signal_6730 ;
    wire new_AGEMA_signal_6731 ;
    wire new_AGEMA_signal_6732 ;
    wire new_AGEMA_signal_6733 ;
    wire new_AGEMA_signal_6734 ;
    wire new_AGEMA_signal_6735 ;
    wire new_AGEMA_signal_6736 ;
    wire new_AGEMA_signal_6737 ;
    wire new_AGEMA_signal_6738 ;
    wire new_AGEMA_signal_6739 ;
    wire new_AGEMA_signal_6740 ;
    wire new_AGEMA_signal_6741 ;
    wire new_AGEMA_signal_6742 ;
    wire new_AGEMA_signal_6743 ;
    wire new_AGEMA_signal_6744 ;
    wire new_AGEMA_signal_6745 ;
    wire new_AGEMA_signal_6746 ;
    wire new_AGEMA_signal_6747 ;
    wire new_AGEMA_signal_6748 ;
    wire new_AGEMA_signal_6749 ;
    wire new_AGEMA_signal_6750 ;
    wire new_AGEMA_signal_6751 ;
    wire new_AGEMA_signal_6752 ;
    wire new_AGEMA_signal_6753 ;
    wire new_AGEMA_signal_6754 ;
    wire new_AGEMA_signal_6755 ;
    wire new_AGEMA_signal_6756 ;
    wire new_AGEMA_signal_6757 ;
    wire new_AGEMA_signal_6758 ;
    wire new_AGEMA_signal_6759 ;
    wire new_AGEMA_signal_6760 ;
    wire new_AGEMA_signal_6761 ;
    wire new_AGEMA_signal_6762 ;
    wire new_AGEMA_signal_6763 ;
    wire new_AGEMA_signal_6764 ;
    wire new_AGEMA_signal_6765 ;
    wire new_AGEMA_signal_6766 ;
    wire new_AGEMA_signal_6767 ;
    wire new_AGEMA_signal_6768 ;
    wire new_AGEMA_signal_6769 ;
    wire new_AGEMA_signal_6770 ;
    wire new_AGEMA_signal_6771 ;
    wire new_AGEMA_signal_6772 ;
    wire new_AGEMA_signal_6773 ;
    wire new_AGEMA_signal_6774 ;
    wire new_AGEMA_signal_6775 ;
    wire new_AGEMA_signal_6776 ;
    wire new_AGEMA_signal_6777 ;
    wire new_AGEMA_signal_6778 ;
    wire new_AGEMA_signal_6779 ;
    wire new_AGEMA_signal_6780 ;
    wire new_AGEMA_signal_6781 ;
    wire new_AGEMA_signal_6782 ;
    wire new_AGEMA_signal_6783 ;
    wire new_AGEMA_signal_6784 ;
    wire new_AGEMA_signal_6785 ;
    wire new_AGEMA_signal_6786 ;
    wire new_AGEMA_signal_6787 ;
    wire new_AGEMA_signal_6788 ;
    wire new_AGEMA_signal_6789 ;
    wire new_AGEMA_signal_6790 ;
    wire new_AGEMA_signal_6791 ;
    wire new_AGEMA_signal_6792 ;
    wire new_AGEMA_signal_6793 ;
    wire new_AGEMA_signal_6794 ;
    wire new_AGEMA_signal_6795 ;
    wire new_AGEMA_signal_6796 ;
    wire new_AGEMA_signal_6797 ;
    wire new_AGEMA_signal_6798 ;
    wire new_AGEMA_signal_6799 ;
    wire new_AGEMA_signal_6800 ;
    wire new_AGEMA_signal_6801 ;
    wire new_AGEMA_signal_6802 ;
    wire new_AGEMA_signal_6803 ;
    wire new_AGEMA_signal_6804 ;
    wire new_AGEMA_signal_6805 ;
    wire new_AGEMA_signal_6806 ;
    wire new_AGEMA_signal_6807 ;
    wire new_AGEMA_signal_6808 ;
    wire new_AGEMA_signal_6809 ;
    wire new_AGEMA_signal_6810 ;
    wire new_AGEMA_signal_6811 ;
    wire new_AGEMA_signal_6812 ;
    wire new_AGEMA_signal_6813 ;
    wire new_AGEMA_signal_6814 ;
    wire new_AGEMA_signal_6815 ;
    wire new_AGEMA_signal_6816 ;
    wire new_AGEMA_signal_6817 ;
    wire new_AGEMA_signal_6818 ;
    wire new_AGEMA_signal_6819 ;
    wire new_AGEMA_signal_6820 ;
    wire new_AGEMA_signal_6821 ;
    wire new_AGEMA_signal_6822 ;
    wire new_AGEMA_signal_6823 ;
    wire new_AGEMA_signal_6824 ;
    wire new_AGEMA_signal_6825 ;
    wire new_AGEMA_signal_6826 ;
    wire new_AGEMA_signal_6827 ;
    wire new_AGEMA_signal_6828 ;
    wire new_AGEMA_signal_6829 ;
    wire new_AGEMA_signal_6830 ;
    wire new_AGEMA_signal_6831 ;
    wire new_AGEMA_signal_6832 ;
    wire new_AGEMA_signal_6833 ;
    wire new_AGEMA_signal_6834 ;
    wire new_AGEMA_signal_6835 ;
    wire new_AGEMA_signal_6836 ;
    wire new_AGEMA_signal_6837 ;
    wire new_AGEMA_signal_6838 ;
    wire new_AGEMA_signal_6839 ;
    wire new_AGEMA_signal_6840 ;
    wire new_AGEMA_signal_6841 ;
    wire new_AGEMA_signal_6842 ;
    wire new_AGEMA_signal_6843 ;
    wire new_AGEMA_signal_6844 ;
    wire new_AGEMA_signal_6845 ;
    wire new_AGEMA_signal_6846 ;
    wire new_AGEMA_signal_6847 ;
    wire new_AGEMA_signal_6848 ;
    wire new_AGEMA_signal_6849 ;
    wire new_AGEMA_signal_6850 ;
    wire new_AGEMA_signal_6851 ;
    wire new_AGEMA_signal_6852 ;
    wire new_AGEMA_signal_6853 ;
    wire new_AGEMA_signal_6854 ;
    wire new_AGEMA_signal_6855 ;
    wire new_AGEMA_signal_6856 ;
    wire new_AGEMA_signal_6857 ;
    wire new_AGEMA_signal_6858 ;
    wire new_AGEMA_signal_6859 ;
    wire new_AGEMA_signal_6860 ;
    wire new_AGEMA_signal_6861 ;
    wire new_AGEMA_signal_6862 ;
    wire new_AGEMA_signal_6863 ;
    wire new_AGEMA_signal_6864 ;
    wire new_AGEMA_signal_6865 ;
    wire new_AGEMA_signal_6866 ;
    wire new_AGEMA_signal_6867 ;
    wire new_AGEMA_signal_6868 ;
    wire new_AGEMA_signal_6869 ;
    wire new_AGEMA_signal_6870 ;
    wire new_AGEMA_signal_6871 ;
    wire new_AGEMA_signal_6872 ;
    wire new_AGEMA_signal_6873 ;
    wire new_AGEMA_signal_6874 ;
    wire new_AGEMA_signal_6875 ;
    wire new_AGEMA_signal_6876 ;
    wire new_AGEMA_signal_6877 ;
    wire new_AGEMA_signal_6878 ;
    wire new_AGEMA_signal_6879 ;
    wire new_AGEMA_signal_6880 ;
    wire new_AGEMA_signal_6881 ;
    wire new_AGEMA_signal_6882 ;
    wire new_AGEMA_signal_6883 ;
    wire new_AGEMA_signal_6884 ;
    wire new_AGEMA_signal_6885 ;
    wire new_AGEMA_signal_6886 ;
    wire new_AGEMA_signal_6887 ;
    wire new_AGEMA_signal_6888 ;
    wire new_AGEMA_signal_6889 ;
    wire new_AGEMA_signal_6890 ;
    wire new_AGEMA_signal_6891 ;
    wire new_AGEMA_signal_6892 ;
    wire new_AGEMA_signal_6893 ;
    wire new_AGEMA_signal_6894 ;
    wire new_AGEMA_signal_6895 ;
    wire new_AGEMA_signal_6896 ;
    wire new_AGEMA_signal_6897 ;
    wire new_AGEMA_signal_6898 ;
    wire new_AGEMA_signal_6899 ;
    wire new_AGEMA_signal_6900 ;
    wire new_AGEMA_signal_6901 ;
    wire new_AGEMA_signal_6902 ;
    wire new_AGEMA_signal_6903 ;
    wire new_AGEMA_signal_6904 ;
    wire new_AGEMA_signal_6905 ;
    wire new_AGEMA_signal_6906 ;
    wire new_AGEMA_signal_6907 ;
    wire new_AGEMA_signal_6908 ;
    wire new_AGEMA_signal_6909 ;
    wire new_AGEMA_signal_6910 ;
    wire new_AGEMA_signal_6911 ;
    wire new_AGEMA_signal_6912 ;
    wire new_AGEMA_signal_6913 ;
    wire new_AGEMA_signal_6914 ;
    wire new_AGEMA_signal_6915 ;
    wire new_AGEMA_signal_6916 ;
    wire new_AGEMA_signal_6917 ;
    wire new_AGEMA_signal_6918 ;
    wire new_AGEMA_signal_6919 ;
    wire new_AGEMA_signal_6920 ;
    wire new_AGEMA_signal_6921 ;
    wire new_AGEMA_signal_6922 ;
    wire new_AGEMA_signal_6923 ;
    wire new_AGEMA_signal_6924 ;
    wire new_AGEMA_signal_6925 ;
    wire new_AGEMA_signal_6926 ;
    wire new_AGEMA_signal_6927 ;
    wire new_AGEMA_signal_6928 ;
    wire new_AGEMA_signal_6929 ;
    wire new_AGEMA_signal_6930 ;
    wire new_AGEMA_signal_6931 ;
    wire new_AGEMA_signal_6932 ;
    wire new_AGEMA_signal_6933 ;
    wire new_AGEMA_signal_6934 ;
    wire new_AGEMA_signal_6935 ;
    wire new_AGEMA_signal_6936 ;
    wire new_AGEMA_signal_6937 ;
    wire new_AGEMA_signal_6938 ;
    wire new_AGEMA_signal_6939 ;
    wire new_AGEMA_signal_6940 ;
    wire new_AGEMA_signal_6941 ;
    wire new_AGEMA_signal_6942 ;
    wire new_AGEMA_signal_6943 ;
    wire new_AGEMA_signal_6944 ;
    wire new_AGEMA_signal_6945 ;
    wire new_AGEMA_signal_6946 ;
    wire new_AGEMA_signal_6947 ;
    wire new_AGEMA_signal_6948 ;
    wire new_AGEMA_signal_6949 ;
    wire new_AGEMA_signal_6950 ;
    wire new_AGEMA_signal_6951 ;
    wire new_AGEMA_signal_6952 ;
    wire new_AGEMA_signal_6953 ;
    wire new_AGEMA_signal_6954 ;
    wire new_AGEMA_signal_6955 ;
    wire new_AGEMA_signal_6956 ;
    wire new_AGEMA_signal_6957 ;
    wire new_AGEMA_signal_6958 ;
    wire new_AGEMA_signal_6959 ;
    wire new_AGEMA_signal_6960 ;
    wire new_AGEMA_signal_6961 ;
    wire new_AGEMA_signal_6962 ;
    wire new_AGEMA_signal_6963 ;
    wire new_AGEMA_signal_6964 ;
    wire new_AGEMA_signal_6965 ;
    wire new_AGEMA_signal_6966 ;
    wire new_AGEMA_signal_6967 ;
    wire new_AGEMA_signal_6968 ;
    wire new_AGEMA_signal_6969 ;
    wire new_AGEMA_signal_6970 ;
    wire new_AGEMA_signal_6971 ;
    wire new_AGEMA_signal_6972 ;
    wire new_AGEMA_signal_6973 ;
    wire new_AGEMA_signal_6974 ;
    wire new_AGEMA_signal_6975 ;
    wire new_AGEMA_signal_6976 ;
    wire new_AGEMA_signal_6977 ;
    wire new_AGEMA_signal_6978 ;
    wire new_AGEMA_signal_6979 ;
    wire new_AGEMA_signal_6980 ;
    wire new_AGEMA_signal_6981 ;
    wire new_AGEMA_signal_6982 ;
    wire new_AGEMA_signal_6983 ;
    wire new_AGEMA_signal_6984 ;
    wire new_AGEMA_signal_6985 ;
    wire new_AGEMA_signal_6986 ;
    wire new_AGEMA_signal_6987 ;
    wire new_AGEMA_signal_6988 ;
    wire new_AGEMA_signal_6989 ;
    wire new_AGEMA_signal_6990 ;
    wire new_AGEMA_signal_6991 ;
    wire new_AGEMA_signal_6992 ;
    wire new_AGEMA_signal_6993 ;
    wire new_AGEMA_signal_6994 ;
    wire new_AGEMA_signal_6995 ;
    wire new_AGEMA_signal_6996 ;
    wire new_AGEMA_signal_6997 ;
    wire new_AGEMA_signal_6998 ;
    wire new_AGEMA_signal_6999 ;
    wire new_AGEMA_signal_7000 ;
    wire new_AGEMA_signal_7001 ;
    wire new_AGEMA_signal_7002 ;
    wire new_AGEMA_signal_7003 ;
    wire new_AGEMA_signal_7004 ;
    wire new_AGEMA_signal_7005 ;
    wire new_AGEMA_signal_7006 ;
    wire new_AGEMA_signal_7007 ;
    wire new_AGEMA_signal_7008 ;
    wire new_AGEMA_signal_7009 ;
    wire new_AGEMA_signal_7010 ;
    wire new_AGEMA_signal_7011 ;
    wire new_AGEMA_signal_7012 ;
    wire new_AGEMA_signal_7013 ;
    wire new_AGEMA_signal_7014 ;
    wire new_AGEMA_signal_7015 ;
    wire new_AGEMA_signal_7016 ;
    wire new_AGEMA_signal_7017 ;
    wire new_AGEMA_signal_7018 ;
    wire new_AGEMA_signal_7019 ;
    wire new_AGEMA_signal_7020 ;
    wire new_AGEMA_signal_7021 ;
    wire new_AGEMA_signal_7022 ;
    wire new_AGEMA_signal_7023 ;
    wire new_AGEMA_signal_7024 ;
    wire new_AGEMA_signal_7025 ;
    wire new_AGEMA_signal_7026 ;
    wire new_AGEMA_signal_7027 ;
    wire new_AGEMA_signal_7028 ;
    wire new_AGEMA_signal_7029 ;
    wire new_AGEMA_signal_7030 ;
    wire new_AGEMA_signal_7031 ;
    wire new_AGEMA_signal_7032 ;
    wire new_AGEMA_signal_7033 ;
    wire new_AGEMA_signal_7034 ;
    wire new_AGEMA_signal_7035 ;
    wire new_AGEMA_signal_7036 ;
    wire new_AGEMA_signal_7037 ;
    wire new_AGEMA_signal_7038 ;
    wire new_AGEMA_signal_7039 ;
    wire new_AGEMA_signal_7040 ;
    wire new_AGEMA_signal_7041 ;
    wire new_AGEMA_signal_7042 ;
    wire new_AGEMA_signal_7043 ;
    wire new_AGEMA_signal_7044 ;
    wire new_AGEMA_signal_7045 ;
    wire new_AGEMA_signal_7046 ;
    wire new_AGEMA_signal_7047 ;
    wire new_AGEMA_signal_7048 ;
    wire new_AGEMA_signal_7049 ;
    wire new_AGEMA_signal_7050 ;
    wire new_AGEMA_signal_7051 ;
    wire new_AGEMA_signal_7052 ;
    wire new_AGEMA_signal_7053 ;
    wire new_AGEMA_signal_7054 ;
    wire new_AGEMA_signal_7055 ;
    wire new_AGEMA_signal_7056 ;
    wire new_AGEMA_signal_7057 ;
    wire new_AGEMA_signal_7058 ;
    wire new_AGEMA_signal_7059 ;
    wire new_AGEMA_signal_7060 ;
    wire new_AGEMA_signal_7061 ;
    wire new_AGEMA_signal_7062 ;
    wire new_AGEMA_signal_7063 ;
    wire new_AGEMA_signal_7064 ;
    wire new_AGEMA_signal_7065 ;
    wire new_AGEMA_signal_7066 ;
    wire new_AGEMA_signal_7067 ;
    wire new_AGEMA_signal_7068 ;
    wire new_AGEMA_signal_7069 ;
    wire new_AGEMA_signal_7070 ;
    wire new_AGEMA_signal_7071 ;
    wire new_AGEMA_signal_7072 ;
    wire new_AGEMA_signal_7073 ;
    wire new_AGEMA_signal_7074 ;
    wire new_AGEMA_signal_7075 ;
    wire new_AGEMA_signal_7076 ;
    wire new_AGEMA_signal_7077 ;
    wire new_AGEMA_signal_7078 ;
    wire new_AGEMA_signal_7079 ;
    wire new_AGEMA_signal_7080 ;
    wire new_AGEMA_signal_7081 ;
    wire new_AGEMA_signal_7082 ;
    wire new_AGEMA_signal_7083 ;
    wire new_AGEMA_signal_7084 ;
    wire new_AGEMA_signal_7085 ;
    wire new_AGEMA_signal_7086 ;
    wire new_AGEMA_signal_7087 ;
    wire new_AGEMA_signal_7088 ;
    wire new_AGEMA_signal_7089 ;
    wire new_AGEMA_signal_7090 ;
    wire new_AGEMA_signal_7091 ;
    wire new_AGEMA_signal_7092 ;
    wire new_AGEMA_signal_7093 ;
    wire new_AGEMA_signal_7094 ;
    wire new_AGEMA_signal_7095 ;
    wire new_AGEMA_signal_7096 ;
    wire new_AGEMA_signal_7097 ;
    wire new_AGEMA_signal_7098 ;
    wire new_AGEMA_signal_7099 ;
    wire new_AGEMA_signal_7100 ;
    wire new_AGEMA_signal_7101 ;
    wire new_AGEMA_signal_7102 ;
    wire new_AGEMA_signal_7103 ;
    wire new_AGEMA_signal_7104 ;
    wire new_AGEMA_signal_7105 ;
    wire new_AGEMA_signal_7106 ;
    wire new_AGEMA_signal_7107 ;
    wire new_AGEMA_signal_7108 ;
    wire new_AGEMA_signal_7109 ;
    wire new_AGEMA_signal_7110 ;
    wire new_AGEMA_signal_7111 ;
    wire new_AGEMA_signal_7112 ;
    wire new_AGEMA_signal_7113 ;
    wire new_AGEMA_signal_7114 ;
    wire new_AGEMA_signal_7115 ;
    wire new_AGEMA_signal_7116 ;
    wire new_AGEMA_signal_7117 ;
    wire new_AGEMA_signal_7118 ;
    wire new_AGEMA_signal_7119 ;
    wire new_AGEMA_signal_7120 ;
    wire new_AGEMA_signal_7121 ;
    wire new_AGEMA_signal_7122 ;
    wire new_AGEMA_signal_7123 ;
    wire new_AGEMA_signal_7124 ;
    wire new_AGEMA_signal_7125 ;
    wire new_AGEMA_signal_7126 ;
    wire new_AGEMA_signal_7127 ;
    wire new_AGEMA_signal_7128 ;
    wire new_AGEMA_signal_7129 ;
    wire new_AGEMA_signal_7130 ;
    wire new_AGEMA_signal_7131 ;
    wire new_AGEMA_signal_7132 ;
    wire new_AGEMA_signal_7133 ;
    wire new_AGEMA_signal_7134 ;
    wire new_AGEMA_signal_7135 ;
    wire new_AGEMA_signal_7136 ;
    wire new_AGEMA_signal_7137 ;
    wire new_AGEMA_signal_7138 ;
    wire new_AGEMA_signal_7139 ;
    wire new_AGEMA_signal_7140 ;
    wire new_AGEMA_signal_7141 ;
    wire new_AGEMA_signal_7142 ;
    wire new_AGEMA_signal_7143 ;
    wire new_AGEMA_signal_7144 ;
    wire new_AGEMA_signal_7145 ;
    wire new_AGEMA_signal_7146 ;
    wire new_AGEMA_signal_7147 ;
    wire new_AGEMA_signal_7148 ;
    wire new_AGEMA_signal_7149 ;
    wire new_AGEMA_signal_7150 ;
    wire new_AGEMA_signal_7151 ;
    wire new_AGEMA_signal_7152 ;
    wire new_AGEMA_signal_7153 ;
    wire new_AGEMA_signal_7154 ;
    wire new_AGEMA_signal_7155 ;
    wire new_AGEMA_signal_7156 ;
    wire new_AGEMA_signal_7157 ;
    wire new_AGEMA_signal_7158 ;
    wire new_AGEMA_signal_7159 ;
    wire new_AGEMA_signal_7160 ;
    wire new_AGEMA_signal_7161 ;
    wire new_AGEMA_signal_7162 ;
    wire new_AGEMA_signal_7163 ;
    wire new_AGEMA_signal_7164 ;
    wire new_AGEMA_signal_7165 ;
    wire new_AGEMA_signal_7166 ;
    wire new_AGEMA_signal_7167 ;
    wire new_AGEMA_signal_7168 ;
    wire new_AGEMA_signal_7169 ;
    wire new_AGEMA_signal_7170 ;
    wire new_AGEMA_signal_7171 ;
    wire new_AGEMA_signal_7172 ;
    wire new_AGEMA_signal_7173 ;
    wire new_AGEMA_signal_7174 ;
    wire new_AGEMA_signal_7175 ;
    wire new_AGEMA_signal_7176 ;
    wire new_AGEMA_signal_7177 ;
    wire new_AGEMA_signal_7178 ;
    wire new_AGEMA_signal_7179 ;
    wire new_AGEMA_signal_7180 ;
    wire new_AGEMA_signal_7181 ;
    wire new_AGEMA_signal_7182 ;
    wire new_AGEMA_signal_7183 ;
    wire new_AGEMA_signal_7184 ;
    wire new_AGEMA_signal_7185 ;
    wire new_AGEMA_signal_7186 ;
    wire new_AGEMA_signal_7187 ;
    wire new_AGEMA_signal_7188 ;
    wire new_AGEMA_signal_7189 ;
    wire new_AGEMA_signal_7190 ;
    wire new_AGEMA_signal_7191 ;
    wire new_AGEMA_signal_7192 ;
    wire new_AGEMA_signal_7193 ;
    wire new_AGEMA_signal_7194 ;
    wire new_AGEMA_signal_7195 ;
    wire new_AGEMA_signal_7196 ;
    wire new_AGEMA_signal_7197 ;
    wire new_AGEMA_signal_7198 ;
    wire new_AGEMA_signal_7199 ;
    wire new_AGEMA_signal_7200 ;
    wire new_AGEMA_signal_7201 ;
    wire new_AGEMA_signal_7202 ;
    wire new_AGEMA_signal_7203 ;
    wire new_AGEMA_signal_7204 ;
    wire new_AGEMA_signal_7205 ;
    wire new_AGEMA_signal_7206 ;
    wire new_AGEMA_signal_7207 ;
    wire new_AGEMA_signal_7208 ;
    wire new_AGEMA_signal_7209 ;
    wire new_AGEMA_signal_7210 ;
    wire new_AGEMA_signal_7211 ;
    wire new_AGEMA_signal_7212 ;
    wire new_AGEMA_signal_7213 ;
    wire new_AGEMA_signal_7214 ;
    wire new_AGEMA_signal_7215 ;
    wire new_AGEMA_signal_7216 ;
    wire new_AGEMA_signal_7217 ;
    wire new_AGEMA_signal_7218 ;
    wire new_AGEMA_signal_7219 ;
    wire new_AGEMA_signal_7220 ;
    wire new_AGEMA_signal_7221 ;
    wire new_AGEMA_signal_7222 ;
    wire new_AGEMA_signal_7223 ;
    wire new_AGEMA_signal_7224 ;
    wire new_AGEMA_signal_7225 ;
    wire new_AGEMA_signal_7226 ;
    wire new_AGEMA_signal_7227 ;
    wire new_AGEMA_signal_7228 ;
    wire new_AGEMA_signal_7229 ;
    wire new_AGEMA_signal_7230 ;
    wire new_AGEMA_signal_7231 ;
    wire new_AGEMA_signal_7232 ;
    wire new_AGEMA_signal_7233 ;
    wire new_AGEMA_signal_7234 ;
    wire new_AGEMA_signal_7235 ;
    wire new_AGEMA_signal_7236 ;
    wire new_AGEMA_signal_7237 ;
    wire new_AGEMA_signal_7238 ;
    wire new_AGEMA_signal_7239 ;
    wire new_AGEMA_signal_7240 ;
    wire new_AGEMA_signal_7241 ;
    wire new_AGEMA_signal_7242 ;
    wire new_AGEMA_signal_7243 ;
    wire new_AGEMA_signal_7244 ;
    wire new_AGEMA_signal_7245 ;
    wire new_AGEMA_signal_7246 ;
    wire new_AGEMA_signal_7247 ;
    wire new_AGEMA_signal_7248 ;
    wire new_AGEMA_signal_7249 ;
    wire new_AGEMA_signal_7250 ;
    wire new_AGEMA_signal_7251 ;
    wire new_AGEMA_signal_7252 ;
    wire new_AGEMA_signal_7253 ;
    wire new_AGEMA_signal_7254 ;
    wire new_AGEMA_signal_7255 ;
    wire new_AGEMA_signal_7256 ;
    wire new_AGEMA_signal_7257 ;
    wire new_AGEMA_signal_7258 ;
    wire new_AGEMA_signal_7259 ;
    wire new_AGEMA_signal_7260 ;
    wire new_AGEMA_signal_7261 ;
    wire new_AGEMA_signal_7262 ;
    wire new_AGEMA_signal_7263 ;
    wire new_AGEMA_signal_7264 ;
    wire new_AGEMA_signal_7265 ;
    wire new_AGEMA_signal_7266 ;
    wire new_AGEMA_signal_7267 ;
    wire new_AGEMA_signal_7268 ;
    wire new_AGEMA_signal_7269 ;
    wire new_AGEMA_signal_7270 ;
    wire new_AGEMA_signal_7271 ;
    wire new_AGEMA_signal_7272 ;
    wire new_AGEMA_signal_7273 ;
    wire new_AGEMA_signal_7274 ;
    wire new_AGEMA_signal_7275 ;
    wire new_AGEMA_signal_7276 ;
    wire new_AGEMA_signal_7277 ;
    wire new_AGEMA_signal_7278 ;
    wire new_AGEMA_signal_7279 ;
    wire new_AGEMA_signal_7280 ;
    wire new_AGEMA_signal_7281 ;
    wire new_AGEMA_signal_7282 ;
    wire new_AGEMA_signal_7283 ;
    wire new_AGEMA_signal_7284 ;
    wire new_AGEMA_signal_7285 ;
    wire new_AGEMA_signal_7286 ;
    wire new_AGEMA_signal_7287 ;
    wire new_AGEMA_signal_7288 ;
    wire new_AGEMA_signal_7289 ;
    wire new_AGEMA_signal_7290 ;
    wire new_AGEMA_signal_7291 ;
    wire new_AGEMA_signal_7292 ;
    wire new_AGEMA_signal_7293 ;
    wire new_AGEMA_signal_7294 ;
    wire new_AGEMA_signal_7295 ;
    wire new_AGEMA_signal_7296 ;
    wire new_AGEMA_signal_7297 ;
    wire new_AGEMA_signal_7298 ;
    wire new_AGEMA_signal_7299 ;
    wire new_AGEMA_signal_7300 ;
    wire new_AGEMA_signal_7301 ;
    wire new_AGEMA_signal_7302 ;
    wire new_AGEMA_signal_7303 ;
    wire new_AGEMA_signal_7304 ;
    wire new_AGEMA_signal_7305 ;
    wire new_AGEMA_signal_7306 ;
    wire new_AGEMA_signal_7307 ;
    wire new_AGEMA_signal_7308 ;
    wire new_AGEMA_signal_7309 ;
    wire new_AGEMA_signal_7310 ;
    wire new_AGEMA_signal_7311 ;
    wire new_AGEMA_signal_7312 ;
    wire new_AGEMA_signal_7313 ;
    wire new_AGEMA_signal_7314 ;
    wire new_AGEMA_signal_7315 ;
    wire new_AGEMA_signal_7316 ;
    wire new_AGEMA_signal_7317 ;
    wire new_AGEMA_signal_7318 ;
    wire new_AGEMA_signal_7319 ;
    wire new_AGEMA_signal_7320 ;
    wire new_AGEMA_signal_7321 ;
    wire new_AGEMA_signal_7322 ;
    wire new_AGEMA_signal_7323 ;
    wire new_AGEMA_signal_7324 ;
    wire new_AGEMA_signal_7325 ;
    wire new_AGEMA_signal_7326 ;
    wire new_AGEMA_signal_7327 ;
    wire new_AGEMA_signal_7328 ;
    wire new_AGEMA_signal_7329 ;
    wire new_AGEMA_signal_7330 ;
    wire new_AGEMA_signal_7331 ;
    wire new_AGEMA_signal_7332 ;
    wire new_AGEMA_signal_7333 ;
    wire new_AGEMA_signal_7334 ;
    wire new_AGEMA_signal_7335 ;
    wire new_AGEMA_signal_7336 ;
    wire new_AGEMA_signal_7337 ;
    wire new_AGEMA_signal_7338 ;
    wire new_AGEMA_signal_7339 ;
    wire new_AGEMA_signal_7340 ;
    wire new_AGEMA_signal_7341 ;
    wire new_AGEMA_signal_7342 ;
    wire new_AGEMA_signal_7343 ;
    wire new_AGEMA_signal_7344 ;
    wire new_AGEMA_signal_7345 ;
    wire new_AGEMA_signal_7346 ;
    wire new_AGEMA_signal_7347 ;
    wire new_AGEMA_signal_7348 ;
    wire new_AGEMA_signal_7349 ;
    wire new_AGEMA_signal_7350 ;
    wire new_AGEMA_signal_7351 ;
    wire new_AGEMA_signal_7352 ;
    wire new_AGEMA_signal_7353 ;
    wire new_AGEMA_signal_7354 ;
    wire new_AGEMA_signal_7355 ;
    wire new_AGEMA_signal_7356 ;
    wire new_AGEMA_signal_7357 ;
    wire new_AGEMA_signal_7358 ;
    wire new_AGEMA_signal_7359 ;
    wire new_AGEMA_signal_7360 ;
    wire new_AGEMA_signal_7361 ;
    wire new_AGEMA_signal_7362 ;
    wire new_AGEMA_signal_7363 ;
    wire new_AGEMA_signal_7364 ;
    wire new_AGEMA_signal_7365 ;
    wire new_AGEMA_signal_7366 ;
    wire new_AGEMA_signal_7367 ;
    wire new_AGEMA_signal_7368 ;
    wire new_AGEMA_signal_7369 ;
    wire new_AGEMA_signal_7370 ;
    wire new_AGEMA_signal_7371 ;
    wire new_AGEMA_signal_7372 ;
    wire new_AGEMA_signal_7373 ;
    wire new_AGEMA_signal_7374 ;
    wire new_AGEMA_signal_7375 ;
    wire new_AGEMA_signal_7376 ;
    wire new_AGEMA_signal_7377 ;
    wire new_AGEMA_signal_7378 ;
    wire new_AGEMA_signal_7379 ;
    wire new_AGEMA_signal_7380 ;
    wire new_AGEMA_signal_7381 ;
    wire new_AGEMA_signal_7382 ;
    wire new_AGEMA_signal_7383 ;
    wire new_AGEMA_signal_7384 ;
    wire new_AGEMA_signal_7385 ;
    wire new_AGEMA_signal_7386 ;
    wire new_AGEMA_signal_7387 ;
    wire new_AGEMA_signal_7388 ;
    wire new_AGEMA_signal_7389 ;
    wire new_AGEMA_signal_7390 ;
    wire new_AGEMA_signal_7391 ;
    wire new_AGEMA_signal_7392 ;
    wire new_AGEMA_signal_7393 ;
    wire new_AGEMA_signal_7394 ;
    wire new_AGEMA_signal_7395 ;
    wire new_AGEMA_signal_7396 ;
    wire new_AGEMA_signal_7397 ;
    wire new_AGEMA_signal_7398 ;
    wire new_AGEMA_signal_7399 ;
    wire new_AGEMA_signal_7400 ;
    wire new_AGEMA_signal_7401 ;
    wire new_AGEMA_signal_7402 ;
    wire new_AGEMA_signal_7403 ;
    wire new_AGEMA_signal_7404 ;
    wire new_AGEMA_signal_7405 ;
    wire new_AGEMA_signal_7406 ;
    wire new_AGEMA_signal_7407 ;
    wire new_AGEMA_signal_7408 ;
    wire new_AGEMA_signal_7409 ;
    wire new_AGEMA_signal_7410 ;
    wire new_AGEMA_signal_7411 ;
    wire new_AGEMA_signal_7412 ;
    wire new_AGEMA_signal_7413 ;
    wire new_AGEMA_signal_7414 ;
    wire new_AGEMA_signal_7415 ;
    wire new_AGEMA_signal_7416 ;
    wire new_AGEMA_signal_7417 ;
    wire new_AGEMA_signal_7418 ;
    wire new_AGEMA_signal_7419 ;
    wire new_AGEMA_signal_7420 ;
    wire new_AGEMA_signal_7421 ;
    wire new_AGEMA_signal_7422 ;
    wire new_AGEMA_signal_7423 ;
    wire new_AGEMA_signal_7424 ;
    wire new_AGEMA_signal_7425 ;
    wire new_AGEMA_signal_7426 ;
    wire new_AGEMA_signal_7427 ;
    wire new_AGEMA_signal_7428 ;
    wire new_AGEMA_signal_7429 ;
    wire new_AGEMA_signal_7430 ;
    wire new_AGEMA_signal_7431 ;
    wire new_AGEMA_signal_7432 ;
    wire new_AGEMA_signal_7433 ;
    wire new_AGEMA_signal_7434 ;
    wire new_AGEMA_signal_7435 ;
    wire new_AGEMA_signal_7436 ;
    wire new_AGEMA_signal_7437 ;
    wire new_AGEMA_signal_7438 ;
    wire new_AGEMA_signal_7439 ;
    wire new_AGEMA_signal_7440 ;
    wire new_AGEMA_signal_7441 ;
    wire new_AGEMA_signal_7442 ;
    wire new_AGEMA_signal_7443 ;
    wire new_AGEMA_signal_7444 ;
    wire new_AGEMA_signal_7445 ;
    wire new_AGEMA_signal_7446 ;
    wire new_AGEMA_signal_7447 ;
    wire new_AGEMA_signal_7448 ;
    wire new_AGEMA_signal_7449 ;
    wire new_AGEMA_signal_7450 ;
    wire new_AGEMA_signal_7451 ;
    wire new_AGEMA_signal_7452 ;
    wire new_AGEMA_signal_7453 ;
    wire new_AGEMA_signal_7454 ;
    wire new_AGEMA_signal_7455 ;
    wire new_AGEMA_signal_7456 ;
    wire new_AGEMA_signal_7457 ;
    wire new_AGEMA_signal_7458 ;
    wire new_AGEMA_signal_7459 ;
    wire new_AGEMA_signal_7460 ;
    wire new_AGEMA_signal_7461 ;
    wire new_AGEMA_signal_7462 ;
    wire new_AGEMA_signal_7463 ;
    wire new_AGEMA_signal_7464 ;
    wire new_AGEMA_signal_7465 ;
    wire new_AGEMA_signal_7466 ;
    wire new_AGEMA_signal_7467 ;
    wire new_AGEMA_signal_7468 ;
    wire new_AGEMA_signal_7469 ;
    wire new_AGEMA_signal_7470 ;
    wire new_AGEMA_signal_7471 ;
    wire new_AGEMA_signal_7472 ;
    wire new_AGEMA_signal_7473 ;
    wire new_AGEMA_signal_7474 ;
    wire new_AGEMA_signal_7475 ;
    wire new_AGEMA_signal_7476 ;
    wire new_AGEMA_signal_7477 ;
    wire new_AGEMA_signal_7478 ;
    wire new_AGEMA_signal_7479 ;
    wire new_AGEMA_signal_7480 ;
    wire new_AGEMA_signal_7481 ;
    wire new_AGEMA_signal_7482 ;
    wire new_AGEMA_signal_7483 ;
    wire new_AGEMA_signal_7484 ;
    wire new_AGEMA_signal_7485 ;
    wire new_AGEMA_signal_7486 ;
    wire new_AGEMA_signal_7487 ;
    wire new_AGEMA_signal_7488 ;
    wire new_AGEMA_signal_7489 ;
    wire new_AGEMA_signal_7490 ;
    wire new_AGEMA_signal_7491 ;
    wire new_AGEMA_signal_7492 ;
    wire new_AGEMA_signal_7493 ;
    wire new_AGEMA_signal_7494 ;
    wire new_AGEMA_signal_7495 ;
    wire new_AGEMA_signal_7496 ;
    wire new_AGEMA_signal_7497 ;
    wire new_AGEMA_signal_7498 ;
    wire new_AGEMA_signal_7499 ;
    wire new_AGEMA_signal_7500 ;
    wire new_AGEMA_signal_7501 ;
    wire new_AGEMA_signal_7502 ;
    wire new_AGEMA_signal_7503 ;
    wire new_AGEMA_signal_7504 ;
    wire new_AGEMA_signal_7505 ;
    wire new_AGEMA_signal_7506 ;
    wire new_AGEMA_signal_7507 ;
    wire new_AGEMA_signal_7508 ;
    wire new_AGEMA_signal_7509 ;
    wire new_AGEMA_signal_7510 ;
    wire new_AGEMA_signal_7511 ;
    wire new_AGEMA_signal_7512 ;
    wire new_AGEMA_signal_7513 ;
    wire new_AGEMA_signal_7514 ;
    wire new_AGEMA_signal_7515 ;
    wire new_AGEMA_signal_7516 ;
    wire new_AGEMA_signal_7517 ;
    wire new_AGEMA_signal_7518 ;
    wire new_AGEMA_signal_7519 ;
    wire new_AGEMA_signal_7520 ;
    wire new_AGEMA_signal_7521 ;
    wire new_AGEMA_signal_7522 ;
    wire new_AGEMA_signal_7523 ;
    wire new_AGEMA_signal_7524 ;
    wire new_AGEMA_signal_7525 ;
    wire new_AGEMA_signal_7526 ;
    wire new_AGEMA_signal_7527 ;
    wire new_AGEMA_signal_7528 ;
    wire new_AGEMA_signal_7529 ;
    wire new_AGEMA_signal_7530 ;
    wire new_AGEMA_signal_7531 ;
    wire new_AGEMA_signal_7532 ;
    wire new_AGEMA_signal_7533 ;
    wire new_AGEMA_signal_7534 ;
    wire new_AGEMA_signal_7535 ;
    wire new_AGEMA_signal_7536 ;
    wire new_AGEMA_signal_7537 ;
    wire new_AGEMA_signal_7538 ;
    wire new_AGEMA_signal_7539 ;
    wire new_AGEMA_signal_7540 ;
    wire new_AGEMA_signal_7541 ;
    wire new_AGEMA_signal_7542 ;
    wire new_AGEMA_signal_7543 ;
    wire new_AGEMA_signal_7544 ;
    wire new_AGEMA_signal_7545 ;
    wire new_AGEMA_signal_7546 ;
    wire new_AGEMA_signal_7547 ;
    wire new_AGEMA_signal_7548 ;
    wire new_AGEMA_signal_7549 ;
    wire new_AGEMA_signal_7550 ;
    wire new_AGEMA_signal_7551 ;
    wire new_AGEMA_signal_7552 ;
    wire new_AGEMA_signal_7553 ;
    wire new_AGEMA_signal_7554 ;
    wire new_AGEMA_signal_7555 ;
    wire new_AGEMA_signal_7556 ;
    wire new_AGEMA_signal_7557 ;
    wire new_AGEMA_signal_7558 ;
    wire new_AGEMA_signal_7559 ;
    wire new_AGEMA_signal_7560 ;
    wire new_AGEMA_signal_7561 ;
    wire new_AGEMA_signal_7562 ;
    wire new_AGEMA_signal_7563 ;
    wire new_AGEMA_signal_7564 ;
    wire new_AGEMA_signal_7565 ;
    wire new_AGEMA_signal_7566 ;
    wire new_AGEMA_signal_7567 ;
    wire new_AGEMA_signal_7568 ;
    wire new_AGEMA_signal_7569 ;
    wire new_AGEMA_signal_7570 ;
    wire new_AGEMA_signal_7571 ;
    wire new_AGEMA_signal_7572 ;
    wire new_AGEMA_signal_7573 ;
    wire new_AGEMA_signal_7574 ;
    wire new_AGEMA_signal_7575 ;
    wire new_AGEMA_signal_7576 ;
    wire new_AGEMA_signal_7577 ;
    wire new_AGEMA_signal_7578 ;
    wire new_AGEMA_signal_7579 ;
    wire new_AGEMA_signal_7580 ;
    wire new_AGEMA_signal_7581 ;
    wire new_AGEMA_signal_7582 ;
    wire new_AGEMA_signal_7583 ;
    wire new_AGEMA_signal_7584 ;
    wire new_AGEMA_signal_7585 ;
    wire new_AGEMA_signal_7586 ;
    wire new_AGEMA_signal_7587 ;
    wire new_AGEMA_signal_7588 ;
    wire new_AGEMA_signal_7589 ;
    wire new_AGEMA_signal_7590 ;
    wire new_AGEMA_signal_7591 ;
    wire new_AGEMA_signal_7592 ;
    wire new_AGEMA_signal_7593 ;
    wire new_AGEMA_signal_7594 ;
    wire new_AGEMA_signal_7595 ;
    wire new_AGEMA_signal_7596 ;
    wire new_AGEMA_signal_7597 ;
    wire new_AGEMA_signal_7598 ;
    wire new_AGEMA_signal_7599 ;
    wire new_AGEMA_signal_7600 ;
    wire new_AGEMA_signal_7601 ;
    wire new_AGEMA_signal_7602 ;
    wire new_AGEMA_signal_7603 ;
    wire new_AGEMA_signal_7604 ;
    wire new_AGEMA_signal_7605 ;
    wire new_AGEMA_signal_7606 ;
    wire new_AGEMA_signal_7607 ;
    wire new_AGEMA_signal_7608 ;
    wire new_AGEMA_signal_7609 ;
    wire new_AGEMA_signal_7610 ;
    wire new_AGEMA_signal_7611 ;
    wire new_AGEMA_signal_7612 ;
    wire new_AGEMA_signal_7613 ;
    wire new_AGEMA_signal_7614 ;
    wire new_AGEMA_signal_7615 ;
    wire new_AGEMA_signal_7616 ;
    wire new_AGEMA_signal_7617 ;
    wire new_AGEMA_signal_7618 ;
    wire new_AGEMA_signal_7619 ;
    wire new_AGEMA_signal_7620 ;
    wire new_AGEMA_signal_7621 ;
    wire new_AGEMA_signal_7622 ;
    wire new_AGEMA_signal_7623 ;
    wire new_AGEMA_signal_7624 ;
    wire new_AGEMA_signal_7625 ;
    wire new_AGEMA_signal_7626 ;
    wire new_AGEMA_signal_7627 ;
    wire new_AGEMA_signal_7628 ;
    wire new_AGEMA_signal_7629 ;
    wire new_AGEMA_signal_7630 ;
    wire new_AGEMA_signal_7631 ;
    wire new_AGEMA_signal_7632 ;
    wire new_AGEMA_signal_7633 ;
    wire new_AGEMA_signal_7634 ;
    wire new_AGEMA_signal_7635 ;
    wire new_AGEMA_signal_7636 ;
    wire new_AGEMA_signal_7637 ;
    wire new_AGEMA_signal_7638 ;
    wire new_AGEMA_signal_7639 ;
    wire new_AGEMA_signal_7640 ;
    wire new_AGEMA_signal_7641 ;
    wire new_AGEMA_signal_7642 ;
    wire new_AGEMA_signal_7643 ;
    wire new_AGEMA_signal_7644 ;
    wire new_AGEMA_signal_7645 ;
    wire new_AGEMA_signal_7646 ;
    wire new_AGEMA_signal_7647 ;
    wire new_AGEMA_signal_7648 ;
    wire new_AGEMA_signal_7649 ;
    wire new_AGEMA_signal_7650 ;
    wire new_AGEMA_signal_7651 ;
    wire new_AGEMA_signal_7652 ;
    wire new_AGEMA_signal_7653 ;
    wire new_AGEMA_signal_7654 ;
    wire new_AGEMA_signal_7655 ;
    wire new_AGEMA_signal_7656 ;
    wire new_AGEMA_signal_7657 ;
    wire new_AGEMA_signal_7658 ;
    wire new_AGEMA_signal_7659 ;
    wire new_AGEMA_signal_7660 ;
    wire new_AGEMA_signal_7661 ;
    wire new_AGEMA_signal_7662 ;
    wire new_AGEMA_signal_7663 ;
    wire new_AGEMA_signal_7664 ;
    wire new_AGEMA_signal_7665 ;
    wire new_AGEMA_signal_7666 ;
    wire new_AGEMA_signal_7667 ;
    wire new_AGEMA_signal_7668 ;
    wire new_AGEMA_signal_7669 ;
    wire new_AGEMA_signal_7670 ;
    wire new_AGEMA_signal_7671 ;
    wire new_AGEMA_signal_7672 ;
    wire new_AGEMA_signal_7673 ;
    wire new_AGEMA_signal_7674 ;
    wire new_AGEMA_signal_7675 ;
    wire new_AGEMA_signal_7676 ;
    wire new_AGEMA_signal_7677 ;
    wire new_AGEMA_signal_7678 ;
    wire new_AGEMA_signal_7679 ;
    wire new_AGEMA_signal_7680 ;
    wire new_AGEMA_signal_7681 ;
    wire new_AGEMA_signal_7682 ;
    wire new_AGEMA_signal_7683 ;
    wire new_AGEMA_signal_7684 ;
    wire new_AGEMA_signal_7685 ;
    wire new_AGEMA_signal_7686 ;
    wire new_AGEMA_signal_7687 ;
    wire new_AGEMA_signal_7688 ;
    wire new_AGEMA_signal_7689 ;
    wire new_AGEMA_signal_7690 ;
    wire new_AGEMA_signal_7691 ;
    wire new_AGEMA_signal_7692 ;
    wire new_AGEMA_signal_7693 ;
    wire new_AGEMA_signal_7694 ;
    wire new_AGEMA_signal_7695 ;
    wire new_AGEMA_signal_7696 ;
    wire new_AGEMA_signal_7697 ;
    wire new_AGEMA_signal_7698 ;
    wire new_AGEMA_signal_7699 ;
    wire new_AGEMA_signal_7700 ;
    wire new_AGEMA_signal_7701 ;
    wire new_AGEMA_signal_7702 ;
    wire new_AGEMA_signal_7703 ;
    wire new_AGEMA_signal_7704 ;
    wire new_AGEMA_signal_7705 ;
    wire new_AGEMA_signal_7706 ;
    wire new_AGEMA_signal_7707 ;
    wire new_AGEMA_signal_7708 ;
    wire new_AGEMA_signal_7709 ;
    wire new_AGEMA_signal_7710 ;
    wire new_AGEMA_signal_7711 ;
    wire new_AGEMA_signal_7712 ;
    wire new_AGEMA_signal_7713 ;
    wire new_AGEMA_signal_7714 ;
    wire new_AGEMA_signal_7715 ;
    wire new_AGEMA_signal_7716 ;
    wire new_AGEMA_signal_7717 ;
    wire new_AGEMA_signal_7718 ;
    wire new_AGEMA_signal_7719 ;
    wire new_AGEMA_signal_7720 ;
    wire new_AGEMA_signal_7721 ;
    wire new_AGEMA_signal_7722 ;
    wire new_AGEMA_signal_7723 ;
    wire new_AGEMA_signal_7724 ;
    wire new_AGEMA_signal_7725 ;
    wire new_AGEMA_signal_7726 ;
    wire new_AGEMA_signal_7727 ;
    wire new_AGEMA_signal_7728 ;
    wire new_AGEMA_signal_7729 ;
    wire new_AGEMA_signal_7730 ;
    wire new_AGEMA_signal_7731 ;
    wire new_AGEMA_signal_7732 ;
    wire new_AGEMA_signal_7733 ;
    wire new_AGEMA_signal_7734 ;
    wire new_AGEMA_signal_7735 ;
    wire new_AGEMA_signal_7736 ;
    wire new_AGEMA_signal_7737 ;
    wire new_AGEMA_signal_7738 ;
    wire new_AGEMA_signal_7739 ;
    wire new_AGEMA_signal_7740 ;
    wire new_AGEMA_signal_7741 ;
    wire new_AGEMA_signal_7742 ;
    wire new_AGEMA_signal_7743 ;
    wire new_AGEMA_signal_7744 ;
    wire new_AGEMA_signal_7745 ;
    wire new_AGEMA_signal_7746 ;
    wire new_AGEMA_signal_7747 ;
    wire new_AGEMA_signal_7748 ;
    wire new_AGEMA_signal_7749 ;
    wire new_AGEMA_signal_7750 ;
    wire new_AGEMA_signal_7751 ;
    wire new_AGEMA_signal_7752 ;
    wire new_AGEMA_signal_7753 ;
    wire new_AGEMA_signal_7754 ;
    wire new_AGEMA_signal_7755 ;
    wire new_AGEMA_signal_7756 ;
    wire new_AGEMA_signal_7757 ;
    wire new_AGEMA_signal_7758 ;
    wire new_AGEMA_signal_7759 ;
    wire new_AGEMA_signal_7760 ;
    wire new_AGEMA_signal_7761 ;
    wire new_AGEMA_signal_7762 ;
    wire new_AGEMA_signal_7763 ;
    wire new_AGEMA_signal_7764 ;
    wire new_AGEMA_signal_7765 ;
    wire new_AGEMA_signal_7766 ;
    wire new_AGEMA_signal_7767 ;
    wire new_AGEMA_signal_7768 ;
    wire new_AGEMA_signal_7769 ;
    wire new_AGEMA_signal_7770 ;
    wire new_AGEMA_signal_7771 ;
    wire new_AGEMA_signal_7772 ;
    wire new_AGEMA_signal_7773 ;
    wire new_AGEMA_signal_7774 ;
    wire new_AGEMA_signal_7775 ;
    wire new_AGEMA_signal_7776 ;
    wire new_AGEMA_signal_7777 ;
    wire new_AGEMA_signal_7778 ;
    wire new_AGEMA_signal_7779 ;
    wire new_AGEMA_signal_7780 ;
    wire new_AGEMA_signal_7781 ;
    wire new_AGEMA_signal_7782 ;
    wire new_AGEMA_signal_7783 ;
    wire new_AGEMA_signal_7784 ;
    wire new_AGEMA_signal_7785 ;
    wire new_AGEMA_signal_7786 ;
    wire new_AGEMA_signal_7787 ;
    wire new_AGEMA_signal_7788 ;
    wire new_AGEMA_signal_7789 ;
    wire new_AGEMA_signal_7790 ;
    wire new_AGEMA_signal_7791 ;
    wire new_AGEMA_signal_7792 ;
    wire new_AGEMA_signal_7793 ;
    wire new_AGEMA_signal_7794 ;
    wire new_AGEMA_signal_7795 ;
    wire new_AGEMA_signal_7796 ;
    wire new_AGEMA_signal_7797 ;
    wire new_AGEMA_signal_7798 ;
    wire new_AGEMA_signal_7799 ;
    wire new_AGEMA_signal_7800 ;
    wire new_AGEMA_signal_7801 ;
    wire new_AGEMA_signal_7802 ;
    wire new_AGEMA_signal_7803 ;
    wire new_AGEMA_signal_7804 ;
    wire new_AGEMA_signal_7805 ;
    wire new_AGEMA_signal_7806 ;
    wire new_AGEMA_signal_7807 ;
    wire new_AGEMA_signal_7808 ;
    wire new_AGEMA_signal_7809 ;
    wire new_AGEMA_signal_7810 ;
    wire new_AGEMA_signal_7811 ;
    wire new_AGEMA_signal_7812 ;
    wire new_AGEMA_signal_7813 ;
    wire new_AGEMA_signal_7814 ;
    wire new_AGEMA_signal_7815 ;
    wire new_AGEMA_signal_7816 ;
    wire new_AGEMA_signal_7817 ;
    wire new_AGEMA_signal_7818 ;
    wire new_AGEMA_signal_7819 ;
    wire new_AGEMA_signal_7820 ;
    wire new_AGEMA_signal_7821 ;
    wire new_AGEMA_signal_7822 ;
    wire new_AGEMA_signal_7823 ;
    wire new_AGEMA_signal_7824 ;
    wire new_AGEMA_signal_7825 ;
    wire new_AGEMA_signal_7826 ;
    wire new_AGEMA_signal_7827 ;
    wire new_AGEMA_signal_7828 ;
    wire new_AGEMA_signal_7829 ;
    wire new_AGEMA_signal_7830 ;
    wire new_AGEMA_signal_7831 ;
    wire new_AGEMA_signal_7832 ;
    wire new_AGEMA_signal_7833 ;
    wire new_AGEMA_signal_7834 ;
    wire new_AGEMA_signal_7835 ;
    wire new_AGEMA_signal_7836 ;
    wire new_AGEMA_signal_7837 ;
    wire new_AGEMA_signal_7838 ;
    wire new_AGEMA_signal_7839 ;
    wire new_AGEMA_signal_7840 ;
    wire new_AGEMA_signal_7841 ;
    wire new_AGEMA_signal_7842 ;
    wire new_AGEMA_signal_7843 ;
    wire new_AGEMA_signal_7844 ;
    wire new_AGEMA_signal_7845 ;
    wire new_AGEMA_signal_7846 ;
    wire new_AGEMA_signal_7847 ;
    wire new_AGEMA_signal_7848 ;
    wire new_AGEMA_signal_7849 ;
    wire new_AGEMA_signal_7850 ;
    wire new_AGEMA_signal_7851 ;
    wire new_AGEMA_signal_7852 ;
    wire new_AGEMA_signal_7853 ;
    wire new_AGEMA_signal_7854 ;
    wire new_AGEMA_signal_7855 ;
    wire new_AGEMA_signal_7856 ;
    wire new_AGEMA_signal_7857 ;
    wire new_AGEMA_signal_7858 ;
    wire new_AGEMA_signal_7859 ;
    wire new_AGEMA_signal_7860 ;
    wire new_AGEMA_signal_7861 ;
    wire new_AGEMA_signal_7862 ;
    wire new_AGEMA_signal_7863 ;
    wire new_AGEMA_signal_7864 ;
    wire new_AGEMA_signal_7865 ;
    wire new_AGEMA_signal_7866 ;
    wire new_AGEMA_signal_7867 ;
    wire new_AGEMA_signal_7868 ;
    wire new_AGEMA_signal_7869 ;
    wire new_AGEMA_signal_7870 ;
    wire new_AGEMA_signal_7871 ;
    wire new_AGEMA_signal_7872 ;
    wire new_AGEMA_signal_7873 ;
    wire new_AGEMA_signal_7874 ;
    wire new_AGEMA_signal_7875 ;
    wire new_AGEMA_signal_7876 ;
    wire new_AGEMA_signal_7877 ;
    wire new_AGEMA_signal_7878 ;
    wire new_AGEMA_signal_7879 ;
    wire new_AGEMA_signal_7880 ;
    wire new_AGEMA_signal_7881 ;
    wire new_AGEMA_signal_7882 ;
    wire new_AGEMA_signal_7883 ;
    wire new_AGEMA_signal_7884 ;
    wire new_AGEMA_signal_7885 ;
    wire new_AGEMA_signal_7886 ;
    wire new_AGEMA_signal_7887 ;
    wire new_AGEMA_signal_7888 ;
    wire new_AGEMA_signal_7889 ;
    wire new_AGEMA_signal_7890 ;
    wire new_AGEMA_signal_7891 ;
    wire new_AGEMA_signal_7892 ;
    wire new_AGEMA_signal_7893 ;
    wire new_AGEMA_signal_7894 ;
    wire new_AGEMA_signal_7895 ;
    wire new_AGEMA_signal_7896 ;
    wire new_AGEMA_signal_7897 ;
    wire new_AGEMA_signal_7898 ;
    wire new_AGEMA_signal_7899 ;
    wire new_AGEMA_signal_7900 ;
    wire new_AGEMA_signal_7901 ;
    wire new_AGEMA_signal_7902 ;
    wire new_AGEMA_signal_7903 ;
    wire new_AGEMA_signal_7904 ;
    wire new_AGEMA_signal_7905 ;
    wire new_AGEMA_signal_7906 ;
    wire new_AGEMA_signal_7907 ;
    wire new_AGEMA_signal_7908 ;
    wire new_AGEMA_signal_7909 ;
    wire new_AGEMA_signal_7910 ;
    wire new_AGEMA_signal_7911 ;
    wire new_AGEMA_signal_7912 ;
    wire new_AGEMA_signal_7913 ;
    wire new_AGEMA_signal_7914 ;
    wire new_AGEMA_signal_7915 ;
    wire new_AGEMA_signal_7916 ;
    wire new_AGEMA_signal_7917 ;
    wire new_AGEMA_signal_7918 ;
    wire new_AGEMA_signal_7919 ;
    wire new_AGEMA_signal_7920 ;
    wire new_AGEMA_signal_7921 ;
    wire new_AGEMA_signal_7922 ;
    wire new_AGEMA_signal_7923 ;
    wire new_AGEMA_signal_7924 ;
    wire new_AGEMA_signal_7925 ;
    wire new_AGEMA_signal_7926 ;
    wire new_AGEMA_signal_7927 ;
    wire new_AGEMA_signal_7928 ;
    wire new_AGEMA_signal_7929 ;
    wire new_AGEMA_signal_7930 ;
    wire new_AGEMA_signal_7931 ;
    wire new_AGEMA_signal_7932 ;
    wire new_AGEMA_signal_7933 ;
    wire new_AGEMA_signal_7934 ;
    wire new_AGEMA_signal_7935 ;
    wire new_AGEMA_signal_7936 ;
    wire new_AGEMA_signal_7937 ;
    wire new_AGEMA_signal_7938 ;
    wire new_AGEMA_signal_7939 ;
    wire new_AGEMA_signal_7940 ;
    wire new_AGEMA_signal_7941 ;
    wire new_AGEMA_signal_7942 ;
    wire new_AGEMA_signal_7943 ;
    wire new_AGEMA_signal_7944 ;
    wire new_AGEMA_signal_7945 ;
    wire new_AGEMA_signal_7946 ;
    wire new_AGEMA_signal_7947 ;
    wire new_AGEMA_signal_7948 ;
    wire new_AGEMA_signal_7949 ;
    wire new_AGEMA_signal_7950 ;
    wire new_AGEMA_signal_7951 ;
    wire new_AGEMA_signal_7952 ;
    wire new_AGEMA_signal_7953 ;
    wire new_AGEMA_signal_7954 ;
    wire new_AGEMA_signal_7955 ;
    wire new_AGEMA_signal_7956 ;
    wire new_AGEMA_signal_7957 ;
    wire new_AGEMA_signal_7958 ;
    wire new_AGEMA_signal_7959 ;
    wire new_AGEMA_signal_7960 ;
    wire new_AGEMA_signal_7961 ;
    wire new_AGEMA_signal_7962 ;
    wire new_AGEMA_signal_7963 ;
    wire new_AGEMA_signal_7964 ;
    wire new_AGEMA_signal_7965 ;
    wire new_AGEMA_signal_7966 ;
    wire new_AGEMA_signal_7967 ;
    wire new_AGEMA_signal_7968 ;
    wire new_AGEMA_signal_7969 ;
    wire new_AGEMA_signal_7970 ;
    wire new_AGEMA_signal_7971 ;
    wire new_AGEMA_signal_7972 ;
    wire new_AGEMA_signal_7973 ;
    wire new_AGEMA_signal_7974 ;
    wire new_AGEMA_signal_7975 ;
    wire new_AGEMA_signal_7976 ;
    wire new_AGEMA_signal_7977 ;
    wire new_AGEMA_signal_7978 ;
    wire new_AGEMA_signal_7979 ;
    wire new_AGEMA_signal_7980 ;
    wire new_AGEMA_signal_7981 ;
    wire new_AGEMA_signal_7982 ;
    wire new_AGEMA_signal_7983 ;
    wire new_AGEMA_signal_7984 ;
    wire new_AGEMA_signal_7985 ;
    wire new_AGEMA_signal_7986 ;
    wire new_AGEMA_signal_7987 ;
    wire new_AGEMA_signal_7988 ;
    wire new_AGEMA_signal_7989 ;
    wire new_AGEMA_signal_7990 ;
    wire new_AGEMA_signal_7991 ;
    wire new_AGEMA_signal_7992 ;
    wire new_AGEMA_signal_7993 ;
    wire new_AGEMA_signal_7994 ;
    wire new_AGEMA_signal_7995 ;
    wire new_AGEMA_signal_7996 ;
    wire new_AGEMA_signal_7997 ;
    wire new_AGEMA_signal_7998 ;
    wire new_AGEMA_signal_7999 ;
    wire new_AGEMA_signal_8000 ;
    wire new_AGEMA_signal_8001 ;
    wire new_AGEMA_signal_8002 ;
    wire new_AGEMA_signal_8003 ;
    wire new_AGEMA_signal_8004 ;
    wire new_AGEMA_signal_8005 ;
    wire new_AGEMA_signal_8006 ;
    wire new_AGEMA_signal_8007 ;
    wire new_AGEMA_signal_8008 ;
    wire new_AGEMA_signal_8009 ;
    wire new_AGEMA_signal_8010 ;
    wire new_AGEMA_signal_8011 ;
    wire new_AGEMA_signal_8012 ;
    wire new_AGEMA_signal_8013 ;
    wire new_AGEMA_signal_8014 ;
    wire new_AGEMA_signal_8015 ;
    wire new_AGEMA_signal_8016 ;
    wire new_AGEMA_signal_8017 ;
    wire new_AGEMA_signal_8018 ;
    wire new_AGEMA_signal_8019 ;
    wire new_AGEMA_signal_8020 ;
    wire new_AGEMA_signal_8021 ;
    wire new_AGEMA_signal_8022 ;
    wire new_AGEMA_signal_8023 ;
    wire new_AGEMA_signal_8024 ;
    wire new_AGEMA_signal_8025 ;
    wire new_AGEMA_signal_8026 ;
    wire new_AGEMA_signal_8027 ;
    wire new_AGEMA_signal_8028 ;
    wire new_AGEMA_signal_8029 ;
    wire new_AGEMA_signal_8030 ;
    wire new_AGEMA_signal_8031 ;
    wire new_AGEMA_signal_8032 ;
    wire new_AGEMA_signal_8033 ;
    wire new_AGEMA_signal_8034 ;
    wire new_AGEMA_signal_8035 ;
    wire new_AGEMA_signal_8036 ;
    wire new_AGEMA_signal_8037 ;
    wire new_AGEMA_signal_8038 ;
    wire new_AGEMA_signal_8039 ;
    wire new_AGEMA_signal_8040 ;
    wire new_AGEMA_signal_8041 ;
    wire new_AGEMA_signal_8042 ;
    wire new_AGEMA_signal_8043 ;
    wire new_AGEMA_signal_8044 ;
    wire new_AGEMA_signal_8045 ;
    wire new_AGEMA_signal_8046 ;
    wire new_AGEMA_signal_8047 ;
    wire new_AGEMA_signal_8048 ;
    wire new_AGEMA_signal_8049 ;
    wire new_AGEMA_signal_8050 ;
    wire new_AGEMA_signal_8051 ;
    wire new_AGEMA_signal_8052 ;
    wire new_AGEMA_signal_8053 ;
    wire new_AGEMA_signal_8054 ;
    wire new_AGEMA_signal_8055 ;
    wire new_AGEMA_signal_8056 ;
    wire new_AGEMA_signal_8057 ;
    wire new_AGEMA_signal_8058 ;
    wire new_AGEMA_signal_8059 ;
    wire new_AGEMA_signal_8060 ;
    wire new_AGEMA_signal_8061 ;
    wire new_AGEMA_signal_8062 ;
    wire new_AGEMA_signal_8063 ;
    wire new_AGEMA_signal_8064 ;
    wire new_AGEMA_signal_8065 ;
    wire new_AGEMA_signal_8066 ;
    wire new_AGEMA_signal_8067 ;
    wire new_AGEMA_signal_8068 ;
    wire new_AGEMA_signal_8069 ;
    wire new_AGEMA_signal_8070 ;
    wire new_AGEMA_signal_8071 ;
    wire new_AGEMA_signal_8072 ;
    wire new_AGEMA_signal_8073 ;
    wire new_AGEMA_signal_8074 ;
    wire new_AGEMA_signal_8075 ;
    wire new_AGEMA_signal_8076 ;
    wire new_AGEMA_signal_8077 ;
    wire new_AGEMA_signal_8078 ;
    wire new_AGEMA_signal_8079 ;
    wire new_AGEMA_signal_8080 ;
    wire new_AGEMA_signal_8081 ;
    wire new_AGEMA_signal_8082 ;
    wire new_AGEMA_signal_8083 ;
    wire new_AGEMA_signal_8084 ;
    wire new_AGEMA_signal_8085 ;
    wire new_AGEMA_signal_8086 ;
    wire new_AGEMA_signal_8087 ;
    wire new_AGEMA_signal_8088 ;
    wire new_AGEMA_signal_8089 ;
    wire new_AGEMA_signal_8090 ;
    wire new_AGEMA_signal_8091 ;
    wire new_AGEMA_signal_8092 ;
    wire new_AGEMA_signal_8093 ;
    wire new_AGEMA_signal_8094 ;
    wire new_AGEMA_signal_8095 ;
    wire new_AGEMA_signal_8096 ;
    wire new_AGEMA_signal_8097 ;
    wire new_AGEMA_signal_8098 ;
    wire new_AGEMA_signal_8099 ;
    wire new_AGEMA_signal_8100 ;
    wire new_AGEMA_signal_8101 ;
    wire new_AGEMA_signal_8102 ;
    wire new_AGEMA_signal_8103 ;
    wire new_AGEMA_signal_8104 ;
    wire new_AGEMA_signal_8105 ;
    wire new_AGEMA_signal_8106 ;
    wire new_AGEMA_signal_8107 ;
    wire new_AGEMA_signal_8108 ;
    wire new_AGEMA_signal_8109 ;
    wire new_AGEMA_signal_8110 ;
    wire new_AGEMA_signal_8111 ;
    wire new_AGEMA_signal_8112 ;
    wire new_AGEMA_signal_8113 ;
    wire new_AGEMA_signal_8114 ;
    wire new_AGEMA_signal_8115 ;
    wire new_AGEMA_signal_8116 ;
    wire new_AGEMA_signal_8117 ;
    wire new_AGEMA_signal_8118 ;
    wire new_AGEMA_signal_8119 ;
    wire new_AGEMA_signal_8120 ;
    wire new_AGEMA_signal_8121 ;
    wire new_AGEMA_signal_8122 ;
    wire new_AGEMA_signal_8123 ;
    wire new_AGEMA_signal_8124 ;
    wire new_AGEMA_signal_8125 ;
    wire new_AGEMA_signal_8126 ;
    wire new_AGEMA_signal_8127 ;
    wire new_AGEMA_signal_8128 ;
    wire new_AGEMA_signal_8129 ;
    wire new_AGEMA_signal_8130 ;
    wire new_AGEMA_signal_8131 ;
    wire new_AGEMA_signal_8132 ;
    wire new_AGEMA_signal_8133 ;
    wire new_AGEMA_signal_8134 ;
    wire new_AGEMA_signal_8135 ;
    wire new_AGEMA_signal_8136 ;
    wire new_AGEMA_signal_8137 ;
    wire new_AGEMA_signal_8138 ;
    wire new_AGEMA_signal_8139 ;
    wire new_AGEMA_signal_8140 ;
    wire new_AGEMA_signal_8141 ;
    wire new_AGEMA_signal_8142 ;
    wire new_AGEMA_signal_8143 ;
    wire new_AGEMA_signal_8144 ;
    wire new_AGEMA_signal_8145 ;
    wire new_AGEMA_signal_8146 ;
    wire new_AGEMA_signal_8147 ;
    wire new_AGEMA_signal_8148 ;
    wire new_AGEMA_signal_8149 ;
    wire new_AGEMA_signal_8150 ;
    wire new_AGEMA_signal_8151 ;
    wire new_AGEMA_signal_8152 ;
    wire new_AGEMA_signal_8153 ;
    wire new_AGEMA_signal_8154 ;
    wire new_AGEMA_signal_8155 ;
    wire new_AGEMA_signal_8156 ;
    wire new_AGEMA_signal_8157 ;
    wire new_AGEMA_signal_8158 ;
    wire new_AGEMA_signal_8159 ;
    wire new_AGEMA_signal_8160 ;
    wire new_AGEMA_signal_8161 ;
    wire new_AGEMA_signal_8162 ;
    wire new_AGEMA_signal_8163 ;
    wire new_AGEMA_signal_8164 ;
    wire new_AGEMA_signal_8165 ;
    wire new_AGEMA_signal_8166 ;
    wire new_AGEMA_signal_8167 ;
    wire new_AGEMA_signal_8168 ;
    wire new_AGEMA_signal_8169 ;
    wire new_AGEMA_signal_8170 ;
    wire new_AGEMA_signal_8171 ;
    wire new_AGEMA_signal_8172 ;
    wire new_AGEMA_signal_8173 ;
    wire new_AGEMA_signal_8174 ;
    wire new_AGEMA_signal_8175 ;
    wire new_AGEMA_signal_8176 ;
    wire new_AGEMA_signal_8177 ;
    wire new_AGEMA_signal_8178 ;
    wire new_AGEMA_signal_8179 ;
    wire new_AGEMA_signal_8180 ;
    wire new_AGEMA_signal_8181 ;
    wire new_AGEMA_signal_8182 ;
    wire new_AGEMA_signal_8183 ;
    wire new_AGEMA_signal_8184 ;
    wire new_AGEMA_signal_8185 ;
    wire new_AGEMA_signal_8186 ;
    wire new_AGEMA_signal_8187 ;
    wire new_AGEMA_signal_8188 ;
    wire new_AGEMA_signal_8189 ;
    wire new_AGEMA_signal_8190 ;
    wire new_AGEMA_signal_8191 ;
    wire new_AGEMA_signal_8192 ;
    wire new_AGEMA_signal_8193 ;
    wire new_AGEMA_signal_8194 ;
    wire new_AGEMA_signal_8195 ;
    wire new_AGEMA_signal_8196 ;
    wire new_AGEMA_signal_8197 ;
    wire new_AGEMA_signal_8198 ;
    wire new_AGEMA_signal_8199 ;
    wire new_AGEMA_signal_8200 ;
    wire new_AGEMA_signal_8201 ;
    wire new_AGEMA_signal_8202 ;
    wire new_AGEMA_signal_8203 ;
    wire new_AGEMA_signal_8204 ;
    wire new_AGEMA_signal_8205 ;
    wire new_AGEMA_signal_8206 ;
    wire new_AGEMA_signal_8207 ;
    wire new_AGEMA_signal_8208 ;
    wire new_AGEMA_signal_8209 ;
    wire new_AGEMA_signal_8210 ;
    wire new_AGEMA_signal_8211 ;
    wire new_AGEMA_signal_8212 ;
    wire new_AGEMA_signal_8213 ;
    wire new_AGEMA_signal_8214 ;
    wire new_AGEMA_signal_8215 ;
    wire new_AGEMA_signal_8216 ;
    wire new_AGEMA_signal_8217 ;
    wire new_AGEMA_signal_8218 ;
    wire new_AGEMA_signal_8219 ;
    wire new_AGEMA_signal_8220 ;
    wire new_AGEMA_signal_8221 ;
    wire new_AGEMA_signal_8222 ;
    wire new_AGEMA_signal_8223 ;
    wire new_AGEMA_signal_8224 ;
    wire new_AGEMA_signal_8225 ;
    wire new_AGEMA_signal_8226 ;
    wire new_AGEMA_signal_8227 ;
    wire new_AGEMA_signal_8228 ;
    wire new_AGEMA_signal_8229 ;
    wire new_AGEMA_signal_8230 ;
    wire new_AGEMA_signal_8231 ;
    wire new_AGEMA_signal_8232 ;
    wire new_AGEMA_signal_8233 ;
    wire new_AGEMA_signal_8234 ;
    wire new_AGEMA_signal_8235 ;
    wire new_AGEMA_signal_8236 ;
    wire new_AGEMA_signal_8237 ;
    wire new_AGEMA_signal_8238 ;
    wire new_AGEMA_signal_8239 ;
    wire new_AGEMA_signal_8240 ;
    wire new_AGEMA_signal_8241 ;
    wire new_AGEMA_signal_8242 ;
    wire new_AGEMA_signal_8243 ;
    wire new_AGEMA_signal_8244 ;
    wire new_AGEMA_signal_8245 ;
    wire new_AGEMA_signal_8246 ;
    wire new_AGEMA_signal_8247 ;
    wire new_AGEMA_signal_8248 ;
    wire new_AGEMA_signal_8249 ;
    wire new_AGEMA_signal_8250 ;
    wire new_AGEMA_signal_8251 ;
    wire new_AGEMA_signal_8252 ;
    wire new_AGEMA_signal_8253 ;
    wire new_AGEMA_signal_8254 ;
    wire new_AGEMA_signal_8255 ;
    wire new_AGEMA_signal_8256 ;
    wire new_AGEMA_signal_8257 ;
    wire new_AGEMA_signal_8258 ;
    wire new_AGEMA_signal_8259 ;
    wire new_AGEMA_signal_8260 ;
    wire new_AGEMA_signal_8261 ;
    wire new_AGEMA_signal_8262 ;
    wire new_AGEMA_signal_8263 ;
    wire new_AGEMA_signal_8264 ;
    wire new_AGEMA_signal_8265 ;
    wire new_AGEMA_signal_8266 ;
    wire new_AGEMA_signal_8267 ;
    wire new_AGEMA_signal_8268 ;
    wire new_AGEMA_signal_8269 ;
    wire new_AGEMA_signal_8270 ;
    wire new_AGEMA_signal_8271 ;
    wire new_AGEMA_signal_8272 ;
    wire new_AGEMA_signal_8273 ;
    wire new_AGEMA_signal_8274 ;
    wire new_AGEMA_signal_8275 ;
    wire new_AGEMA_signal_8276 ;
    wire new_AGEMA_signal_8277 ;
    wire new_AGEMA_signal_8278 ;
    wire new_AGEMA_signal_8279 ;
    wire new_AGEMA_signal_8280 ;
    wire new_AGEMA_signal_8281 ;
    wire new_AGEMA_signal_8282 ;
    wire new_AGEMA_signal_8283 ;
    wire new_AGEMA_signal_8284 ;
    wire new_AGEMA_signal_8285 ;
    wire new_AGEMA_signal_8286 ;
    wire new_AGEMA_signal_8287 ;
    wire new_AGEMA_signal_8288 ;
    wire new_AGEMA_signal_8289 ;
    wire new_AGEMA_signal_8290 ;
    wire new_AGEMA_signal_8291 ;
    wire new_AGEMA_signal_8292 ;
    wire new_AGEMA_signal_8293 ;
    wire new_AGEMA_signal_8294 ;
    wire new_AGEMA_signal_8295 ;
    wire new_AGEMA_signal_8296 ;
    wire new_AGEMA_signal_8297 ;
    wire new_AGEMA_signal_8298 ;
    wire new_AGEMA_signal_8299 ;
    wire new_AGEMA_signal_8300 ;
    wire new_AGEMA_signal_8301 ;
    wire new_AGEMA_signal_8302 ;
    wire new_AGEMA_signal_8303 ;
    wire new_AGEMA_signal_8304 ;
    wire new_AGEMA_signal_8305 ;
    wire new_AGEMA_signal_8306 ;
    wire new_AGEMA_signal_8307 ;
    wire new_AGEMA_signal_8308 ;
    wire new_AGEMA_signal_8309 ;
    wire new_AGEMA_signal_8310 ;
    wire new_AGEMA_signal_8311 ;
    wire new_AGEMA_signal_8312 ;
    wire new_AGEMA_signal_8313 ;
    wire new_AGEMA_signal_8314 ;
    wire new_AGEMA_signal_8315 ;
    wire new_AGEMA_signal_8316 ;
    wire new_AGEMA_signal_8317 ;
    wire new_AGEMA_signal_8318 ;
    wire new_AGEMA_signal_8319 ;
    wire new_AGEMA_signal_8320 ;
    wire new_AGEMA_signal_8321 ;
    wire new_AGEMA_signal_8322 ;
    wire new_AGEMA_signal_8323 ;
    wire new_AGEMA_signal_8324 ;
    wire new_AGEMA_signal_8325 ;
    wire new_AGEMA_signal_8326 ;
    wire new_AGEMA_signal_8327 ;
    wire new_AGEMA_signal_8328 ;
    wire new_AGEMA_signal_8329 ;
    wire new_AGEMA_signal_8330 ;
    wire new_AGEMA_signal_8331 ;
    wire new_AGEMA_signal_8332 ;
    wire new_AGEMA_signal_8333 ;
    wire new_AGEMA_signal_8334 ;
    wire new_AGEMA_signal_8335 ;
    wire new_AGEMA_signal_8336 ;
    wire new_AGEMA_signal_8337 ;
    wire new_AGEMA_signal_8338 ;
    wire new_AGEMA_signal_8339 ;
    wire new_AGEMA_signal_8340 ;
    wire new_AGEMA_signal_8341 ;
    wire new_AGEMA_signal_8342 ;
    wire new_AGEMA_signal_8343 ;
    wire new_AGEMA_signal_8344 ;
    wire new_AGEMA_signal_8345 ;
    wire new_AGEMA_signal_8346 ;
    wire new_AGEMA_signal_8347 ;
    wire new_AGEMA_signal_8348 ;
    wire new_AGEMA_signal_8349 ;
    wire new_AGEMA_signal_8350 ;
    wire new_AGEMA_signal_8351 ;
    wire new_AGEMA_signal_8352 ;
    wire new_AGEMA_signal_8353 ;
    wire new_AGEMA_signal_8354 ;
    wire new_AGEMA_signal_8355 ;
    wire new_AGEMA_signal_8356 ;
    wire new_AGEMA_signal_8357 ;
    wire new_AGEMA_signal_8358 ;
    wire new_AGEMA_signal_8359 ;
    wire new_AGEMA_signal_8360 ;
    wire new_AGEMA_signal_8361 ;
    wire new_AGEMA_signal_8362 ;
    wire new_AGEMA_signal_8363 ;
    wire new_AGEMA_signal_8364 ;
    wire new_AGEMA_signal_8365 ;
    wire new_AGEMA_signal_8366 ;
    wire new_AGEMA_signal_8367 ;
    wire new_AGEMA_signal_8368 ;
    wire new_AGEMA_signal_8369 ;
    wire new_AGEMA_signal_8370 ;
    wire new_AGEMA_signal_8371 ;
    wire new_AGEMA_signal_8372 ;
    wire new_AGEMA_signal_8373 ;
    wire new_AGEMA_signal_8374 ;
    wire new_AGEMA_signal_8375 ;
    wire new_AGEMA_signal_8376 ;
    wire new_AGEMA_signal_8377 ;
    wire new_AGEMA_signal_8378 ;
    wire new_AGEMA_signal_8379 ;
    wire new_AGEMA_signal_8380 ;
    wire new_AGEMA_signal_8381 ;
    wire new_AGEMA_signal_8382 ;
    wire new_AGEMA_signal_8383 ;
    wire new_AGEMA_signal_8384 ;
    wire new_AGEMA_signal_8385 ;
    wire new_AGEMA_signal_8386 ;
    wire new_AGEMA_signal_8387 ;
    wire new_AGEMA_signal_8388 ;
    wire new_AGEMA_signal_8389 ;
    wire new_AGEMA_signal_8390 ;
    wire new_AGEMA_signal_8391 ;
    wire new_AGEMA_signal_8392 ;
    wire new_AGEMA_signal_8393 ;
    wire new_AGEMA_signal_8394 ;
    wire new_AGEMA_signal_8395 ;
    wire new_AGEMA_signal_8396 ;
    wire new_AGEMA_signal_8397 ;
    wire new_AGEMA_signal_8398 ;
    wire new_AGEMA_signal_8399 ;
    wire new_AGEMA_signal_8400 ;
    wire new_AGEMA_signal_8401 ;
    wire new_AGEMA_signal_8402 ;
    wire new_AGEMA_signal_8403 ;
    wire new_AGEMA_signal_8404 ;
    wire new_AGEMA_signal_8405 ;
    wire new_AGEMA_signal_8406 ;
    wire new_AGEMA_signal_8407 ;
    wire new_AGEMA_signal_8408 ;
    wire new_AGEMA_signal_8409 ;
    wire new_AGEMA_signal_8410 ;
    wire new_AGEMA_signal_8411 ;
    wire new_AGEMA_signal_8412 ;
    wire new_AGEMA_signal_8413 ;
    wire new_AGEMA_signal_8414 ;
    wire new_AGEMA_signal_8415 ;
    wire new_AGEMA_signal_8416 ;
    wire new_AGEMA_signal_8417 ;
    wire new_AGEMA_signal_8418 ;
    wire new_AGEMA_signal_8419 ;
    wire new_AGEMA_signal_8420 ;
    wire new_AGEMA_signal_8421 ;
    wire new_AGEMA_signal_8422 ;
    wire new_AGEMA_signal_8423 ;
    wire new_AGEMA_signal_8424 ;
    wire new_AGEMA_signal_8425 ;
    wire new_AGEMA_signal_8426 ;
    wire new_AGEMA_signal_8427 ;
    wire new_AGEMA_signal_8428 ;
    wire new_AGEMA_signal_8429 ;
    wire new_AGEMA_signal_8430 ;
    wire new_AGEMA_signal_8431 ;
    wire new_AGEMA_signal_8432 ;
    wire new_AGEMA_signal_8433 ;
    wire new_AGEMA_signal_8434 ;
    wire new_AGEMA_signal_8435 ;
    wire new_AGEMA_signal_8436 ;
    wire new_AGEMA_signal_8437 ;
    wire new_AGEMA_signal_8438 ;
    wire new_AGEMA_signal_8439 ;
    wire new_AGEMA_signal_8440 ;
    wire new_AGEMA_signal_8441 ;
    wire new_AGEMA_signal_8442 ;
    wire new_AGEMA_signal_8443 ;
    wire new_AGEMA_signal_8444 ;
    wire new_AGEMA_signal_8445 ;
    wire new_AGEMA_signal_8446 ;
    wire new_AGEMA_signal_8447 ;
    wire new_AGEMA_signal_8448 ;
    wire new_AGEMA_signal_8449 ;
    wire new_AGEMA_signal_8450 ;
    wire new_AGEMA_signal_8451 ;
    wire new_AGEMA_signal_8452 ;
    wire new_AGEMA_signal_8453 ;
    wire new_AGEMA_signal_8454 ;
    wire new_AGEMA_signal_8455 ;
    wire new_AGEMA_signal_8456 ;
    wire new_AGEMA_signal_8457 ;
    wire new_AGEMA_signal_8458 ;
    wire new_AGEMA_signal_8459 ;
    wire new_AGEMA_signal_8460 ;
    wire new_AGEMA_signal_8461 ;
    wire new_AGEMA_signal_8462 ;
    wire new_AGEMA_signal_8463 ;
    wire new_AGEMA_signal_8464 ;
    wire new_AGEMA_signal_8465 ;
    wire new_AGEMA_signal_8466 ;
    wire new_AGEMA_signal_8467 ;
    wire new_AGEMA_signal_8468 ;
    wire new_AGEMA_signal_8469 ;
    wire new_AGEMA_signal_8470 ;
    wire new_AGEMA_signal_8471 ;
    wire new_AGEMA_signal_8472 ;
    wire new_AGEMA_signal_8473 ;
    wire new_AGEMA_signal_8474 ;
    wire new_AGEMA_signal_8475 ;
    wire new_AGEMA_signal_8476 ;
    wire new_AGEMA_signal_8477 ;
    wire new_AGEMA_signal_8478 ;
    wire new_AGEMA_signal_8479 ;
    wire new_AGEMA_signal_8480 ;
    wire new_AGEMA_signal_8481 ;
    wire new_AGEMA_signal_8482 ;
    wire new_AGEMA_signal_8483 ;
    wire new_AGEMA_signal_8484 ;
    wire new_AGEMA_signal_8485 ;
    wire new_AGEMA_signal_8486 ;
    wire new_AGEMA_signal_8487 ;
    wire new_AGEMA_signal_8488 ;
    wire new_AGEMA_signal_8489 ;
    wire new_AGEMA_signal_8490 ;
    wire new_AGEMA_signal_8491 ;
    wire new_AGEMA_signal_8492 ;
    wire new_AGEMA_signal_8493 ;
    wire new_AGEMA_signal_8494 ;
    wire new_AGEMA_signal_8495 ;
    wire new_AGEMA_signal_8496 ;
    wire new_AGEMA_signal_8497 ;
    wire new_AGEMA_signal_8498 ;
    wire new_AGEMA_signal_8499 ;
    wire new_AGEMA_signal_8500 ;
    wire new_AGEMA_signal_8501 ;
    wire new_AGEMA_signal_8502 ;
    wire new_AGEMA_signal_8503 ;
    wire new_AGEMA_signal_8504 ;
    wire new_AGEMA_signal_8505 ;
    wire new_AGEMA_signal_8506 ;
    wire new_AGEMA_signal_8507 ;
    wire new_AGEMA_signal_8508 ;
    wire new_AGEMA_signal_8509 ;
    wire new_AGEMA_signal_8510 ;
    wire new_AGEMA_signal_8511 ;
    wire new_AGEMA_signal_8512 ;
    wire new_AGEMA_signal_8513 ;
    wire new_AGEMA_signal_8514 ;
    wire new_AGEMA_signal_8515 ;
    wire new_AGEMA_signal_8516 ;
    wire new_AGEMA_signal_8517 ;
    wire new_AGEMA_signal_8518 ;
    wire new_AGEMA_signal_8519 ;
    wire new_AGEMA_signal_8520 ;
    wire new_AGEMA_signal_8521 ;
    wire new_AGEMA_signal_8522 ;
    wire new_AGEMA_signal_8523 ;
    wire new_AGEMA_signal_8524 ;
    wire new_AGEMA_signal_8525 ;
    wire new_AGEMA_signal_8526 ;
    wire new_AGEMA_signal_8527 ;
    wire new_AGEMA_signal_8528 ;
    wire new_AGEMA_signal_8529 ;
    wire new_AGEMA_signal_8530 ;
    wire new_AGEMA_signal_8531 ;
    wire new_AGEMA_signal_8532 ;
    wire new_AGEMA_signal_8533 ;
    wire new_AGEMA_signal_8534 ;
    wire new_AGEMA_signal_8535 ;
    wire new_AGEMA_signal_8536 ;
    wire new_AGEMA_signal_8537 ;
    wire new_AGEMA_signal_8538 ;
    wire new_AGEMA_signal_8539 ;
    wire new_AGEMA_signal_8540 ;
    wire new_AGEMA_signal_8541 ;
    wire new_AGEMA_signal_8542 ;
    wire new_AGEMA_signal_8543 ;
    wire new_AGEMA_signal_8544 ;
    wire new_AGEMA_signal_8545 ;
    wire new_AGEMA_signal_8546 ;
    wire new_AGEMA_signal_8547 ;
    wire new_AGEMA_signal_8548 ;
    wire new_AGEMA_signal_8549 ;
    wire new_AGEMA_signal_8550 ;
    wire new_AGEMA_signal_8551 ;
    wire new_AGEMA_signal_8552 ;
    wire new_AGEMA_signal_8553 ;
    wire new_AGEMA_signal_8554 ;
    wire new_AGEMA_signal_8555 ;
    wire new_AGEMA_signal_8556 ;
    wire new_AGEMA_signal_8557 ;
    wire new_AGEMA_signal_8558 ;
    wire new_AGEMA_signal_8559 ;
    wire new_AGEMA_signal_8560 ;
    wire new_AGEMA_signal_8561 ;
    wire new_AGEMA_signal_8562 ;
    wire new_AGEMA_signal_8563 ;
    wire new_AGEMA_signal_8564 ;
    wire new_AGEMA_signal_8565 ;
    wire new_AGEMA_signal_8566 ;
    wire new_AGEMA_signal_8567 ;
    wire new_AGEMA_signal_8568 ;
    wire new_AGEMA_signal_8569 ;
    wire new_AGEMA_signal_8570 ;
    wire new_AGEMA_signal_8571 ;
    wire new_AGEMA_signal_8572 ;
    wire new_AGEMA_signal_8573 ;
    wire new_AGEMA_signal_8574 ;
    wire new_AGEMA_signal_8575 ;
    wire new_AGEMA_signal_8576 ;
    wire new_AGEMA_signal_8577 ;
    wire new_AGEMA_signal_8578 ;
    wire new_AGEMA_signal_8579 ;
    wire new_AGEMA_signal_8580 ;
    wire new_AGEMA_signal_8581 ;
    wire new_AGEMA_signal_8582 ;
    wire new_AGEMA_signal_8583 ;
    wire new_AGEMA_signal_8584 ;
    wire new_AGEMA_signal_8585 ;
    wire new_AGEMA_signal_8586 ;
    wire new_AGEMA_signal_8587 ;
    wire new_AGEMA_signal_8588 ;
    wire new_AGEMA_signal_8589 ;
    wire new_AGEMA_signal_8590 ;
    wire new_AGEMA_signal_8591 ;
    wire new_AGEMA_signal_8592 ;
    wire new_AGEMA_signal_8593 ;
    wire new_AGEMA_signal_8594 ;
    wire new_AGEMA_signal_8595 ;
    wire new_AGEMA_signal_8596 ;
    wire new_AGEMA_signal_8597 ;
    wire new_AGEMA_signal_8598 ;
    wire new_AGEMA_signal_8599 ;
    wire new_AGEMA_signal_8600 ;
    wire new_AGEMA_signal_8601 ;
    wire new_AGEMA_signal_8602 ;
    wire new_AGEMA_signal_8603 ;
    wire new_AGEMA_signal_8604 ;
    wire new_AGEMA_signal_8605 ;
    wire new_AGEMA_signal_8606 ;
    wire new_AGEMA_signal_8607 ;
    wire new_AGEMA_signal_8608 ;
    wire new_AGEMA_signal_8609 ;
    wire new_AGEMA_signal_8610 ;
    wire new_AGEMA_signal_8611 ;
    wire new_AGEMA_signal_8612 ;
    wire new_AGEMA_signal_8613 ;
    wire new_AGEMA_signal_8614 ;
    wire new_AGEMA_signal_8615 ;
    wire new_AGEMA_signal_8616 ;
    wire new_AGEMA_signal_8617 ;
    wire new_AGEMA_signal_8618 ;
    wire new_AGEMA_signal_8619 ;
    wire new_AGEMA_signal_8620 ;
    wire new_AGEMA_signal_8621 ;
    wire new_AGEMA_signal_8622 ;
    wire new_AGEMA_signal_8623 ;
    wire new_AGEMA_signal_8624 ;
    wire new_AGEMA_signal_8625 ;
    wire new_AGEMA_signal_8626 ;
    wire new_AGEMA_signal_8627 ;
    wire new_AGEMA_signal_8628 ;
    wire new_AGEMA_signal_8629 ;
    wire new_AGEMA_signal_8630 ;
    wire new_AGEMA_signal_8631 ;
    wire new_AGEMA_signal_8632 ;
    wire new_AGEMA_signal_8633 ;
    wire new_AGEMA_signal_8634 ;
    wire new_AGEMA_signal_8635 ;
    wire new_AGEMA_signal_8636 ;
    wire new_AGEMA_signal_8637 ;
    wire new_AGEMA_signal_8638 ;
    wire new_AGEMA_signal_8639 ;
    wire new_AGEMA_signal_8640 ;
    wire new_AGEMA_signal_8641 ;
    wire new_AGEMA_signal_8642 ;
    wire new_AGEMA_signal_8643 ;
    wire new_AGEMA_signal_8644 ;
    wire new_AGEMA_signal_8645 ;
    wire new_AGEMA_signal_8646 ;
    wire new_AGEMA_signal_8647 ;
    wire new_AGEMA_signal_8648 ;
    wire new_AGEMA_signal_8649 ;
    wire new_AGEMA_signal_8650 ;
    wire new_AGEMA_signal_8651 ;
    wire new_AGEMA_signal_8652 ;
    wire new_AGEMA_signal_8653 ;
    wire new_AGEMA_signal_8654 ;
    wire new_AGEMA_signal_8655 ;
    wire new_AGEMA_signal_8656 ;
    wire new_AGEMA_signal_8657 ;
    wire new_AGEMA_signal_8658 ;
    wire new_AGEMA_signal_8659 ;
    wire new_AGEMA_signal_8660 ;
    wire new_AGEMA_signal_8661 ;
    wire new_AGEMA_signal_8662 ;
    wire new_AGEMA_signal_8663 ;
    wire new_AGEMA_signal_8664 ;
    wire new_AGEMA_signal_8665 ;
    wire new_AGEMA_signal_8666 ;
    wire new_AGEMA_signal_8667 ;
    wire new_AGEMA_signal_8668 ;
    wire new_AGEMA_signal_8669 ;
    wire new_AGEMA_signal_8670 ;
    wire new_AGEMA_signal_8671 ;
    wire new_AGEMA_signal_8672 ;
    wire new_AGEMA_signal_8673 ;
    wire new_AGEMA_signal_8674 ;
    wire new_AGEMA_signal_8675 ;
    wire new_AGEMA_signal_8676 ;
    wire new_AGEMA_signal_8677 ;
    wire new_AGEMA_signal_8678 ;
    wire new_AGEMA_signal_8679 ;
    wire new_AGEMA_signal_8680 ;
    wire new_AGEMA_signal_8681 ;
    wire new_AGEMA_signal_8682 ;
    wire new_AGEMA_signal_8683 ;
    wire new_AGEMA_signal_8684 ;
    wire new_AGEMA_signal_8685 ;
    wire new_AGEMA_signal_8686 ;
    wire new_AGEMA_signal_8687 ;
    wire new_AGEMA_signal_8688 ;
    wire new_AGEMA_signal_8689 ;
    wire new_AGEMA_signal_8690 ;
    wire new_AGEMA_signal_8691 ;
    wire new_AGEMA_signal_8692 ;
    wire new_AGEMA_signal_8693 ;
    wire new_AGEMA_signal_8694 ;
    wire new_AGEMA_signal_8695 ;
    wire new_AGEMA_signal_8696 ;
    wire new_AGEMA_signal_8697 ;
    wire new_AGEMA_signal_8698 ;
    wire new_AGEMA_signal_8699 ;
    wire new_AGEMA_signal_8700 ;
    wire new_AGEMA_signal_8701 ;
    wire new_AGEMA_signal_8702 ;
    wire new_AGEMA_signal_8703 ;
    wire new_AGEMA_signal_8704 ;
    wire new_AGEMA_signal_8705 ;
    wire new_AGEMA_signal_8706 ;
    wire new_AGEMA_signal_8707 ;
    wire new_AGEMA_signal_8708 ;
    wire new_AGEMA_signal_8709 ;
    wire new_AGEMA_signal_8710 ;
    wire new_AGEMA_signal_8711 ;
    wire new_AGEMA_signal_8712 ;
    wire new_AGEMA_signal_8713 ;
    wire new_AGEMA_signal_8714 ;
    wire new_AGEMA_signal_8715 ;
    wire new_AGEMA_signal_8716 ;
    wire new_AGEMA_signal_8717 ;
    wire new_AGEMA_signal_8718 ;
    wire new_AGEMA_signal_8719 ;
    wire new_AGEMA_signal_8720 ;
    wire new_AGEMA_signal_8721 ;
    wire new_AGEMA_signal_8722 ;
    wire new_AGEMA_signal_8723 ;
    wire new_AGEMA_signal_8724 ;
    wire new_AGEMA_signal_8725 ;
    wire new_AGEMA_signal_8726 ;
    wire new_AGEMA_signal_8727 ;
    wire new_AGEMA_signal_8728 ;
    wire new_AGEMA_signal_8729 ;
    wire new_AGEMA_signal_8730 ;
    wire new_AGEMA_signal_8731 ;
    wire new_AGEMA_signal_8732 ;
    wire new_AGEMA_signal_8733 ;
    wire new_AGEMA_signal_8734 ;
    wire new_AGEMA_signal_8735 ;
    wire new_AGEMA_signal_8736 ;
    wire new_AGEMA_signal_8737 ;
    wire new_AGEMA_signal_8738 ;
    wire new_AGEMA_signal_8739 ;
    wire new_AGEMA_signal_8740 ;
    wire new_AGEMA_signal_8741 ;
    wire new_AGEMA_signal_8742 ;
    wire new_AGEMA_signal_8743 ;
    wire new_AGEMA_signal_8744 ;
    wire new_AGEMA_signal_8745 ;
    wire new_AGEMA_signal_8746 ;
    wire new_AGEMA_signal_8747 ;
    wire new_AGEMA_signal_8748 ;
    wire new_AGEMA_signal_8749 ;
    wire new_AGEMA_signal_8750 ;
    wire new_AGEMA_signal_8751 ;
    wire new_AGEMA_signal_8752 ;
    wire new_AGEMA_signal_8753 ;
    wire new_AGEMA_signal_8754 ;
    wire new_AGEMA_signal_8755 ;
    wire new_AGEMA_signal_8756 ;
    wire new_AGEMA_signal_8757 ;
    wire new_AGEMA_signal_8758 ;
    wire new_AGEMA_signal_8759 ;
    wire new_AGEMA_signal_8760 ;
    wire new_AGEMA_signal_8761 ;
    wire new_AGEMA_signal_8762 ;
    wire new_AGEMA_signal_8763 ;
    wire new_AGEMA_signal_8764 ;
    wire new_AGEMA_signal_8765 ;
    wire new_AGEMA_signal_8766 ;
    wire new_AGEMA_signal_8767 ;
    wire new_AGEMA_signal_8768 ;
    wire new_AGEMA_signal_8769 ;
    wire new_AGEMA_signal_8770 ;
    wire new_AGEMA_signal_8771 ;
    wire new_AGEMA_signal_8772 ;
    wire new_AGEMA_signal_8773 ;
    wire new_AGEMA_signal_8774 ;
    wire new_AGEMA_signal_8775 ;
    wire new_AGEMA_signal_8776 ;
    wire new_AGEMA_signal_8777 ;
    wire new_AGEMA_signal_8778 ;
    wire new_AGEMA_signal_8779 ;
    wire new_AGEMA_signal_8780 ;
    wire new_AGEMA_signal_8781 ;
    wire new_AGEMA_signal_8782 ;
    wire new_AGEMA_signal_8783 ;
    wire new_AGEMA_signal_8784 ;
    wire new_AGEMA_signal_8785 ;
    wire new_AGEMA_signal_8786 ;
    wire new_AGEMA_signal_8787 ;
    wire new_AGEMA_signal_8788 ;
    wire new_AGEMA_signal_8789 ;
    wire new_AGEMA_signal_8790 ;
    wire new_AGEMA_signal_8791 ;
    wire new_AGEMA_signal_8792 ;
    wire new_AGEMA_signal_8793 ;
    wire new_AGEMA_signal_8794 ;
    wire new_AGEMA_signal_8795 ;
    wire new_AGEMA_signal_8796 ;
    wire new_AGEMA_signal_8797 ;
    wire new_AGEMA_signal_8798 ;
    wire new_AGEMA_signal_8799 ;
    wire new_AGEMA_signal_8800 ;
    wire new_AGEMA_signal_8801 ;
    wire new_AGEMA_signal_8802 ;
    wire new_AGEMA_signal_8803 ;
    wire new_AGEMA_signal_8804 ;
    wire new_AGEMA_signal_8805 ;
    wire new_AGEMA_signal_8806 ;
    wire new_AGEMA_signal_8807 ;
    wire new_AGEMA_signal_8808 ;
    wire new_AGEMA_signal_8809 ;
    wire new_AGEMA_signal_8810 ;
    wire new_AGEMA_signal_8811 ;
    wire new_AGEMA_signal_8812 ;
    wire new_AGEMA_signal_8813 ;
    wire new_AGEMA_signal_8814 ;
    wire new_AGEMA_signal_8815 ;
    wire new_AGEMA_signal_8816 ;
    wire new_AGEMA_signal_8817 ;
    wire new_AGEMA_signal_8818 ;
    wire new_AGEMA_signal_8819 ;
    wire new_AGEMA_signal_8820 ;
    wire new_AGEMA_signal_8821 ;
    wire new_AGEMA_signal_8822 ;
    wire new_AGEMA_signal_8823 ;
    wire new_AGEMA_signal_8824 ;
    wire new_AGEMA_signal_8825 ;
    wire new_AGEMA_signal_8826 ;
    wire new_AGEMA_signal_8827 ;
    wire new_AGEMA_signal_8828 ;
    wire new_AGEMA_signal_8829 ;
    wire new_AGEMA_signal_8830 ;
    wire new_AGEMA_signal_8831 ;
    wire new_AGEMA_signal_8832 ;
    wire new_AGEMA_signal_8833 ;
    wire new_AGEMA_signal_8834 ;
    wire new_AGEMA_signal_8835 ;
    wire new_AGEMA_signal_8836 ;
    wire new_AGEMA_signal_8837 ;
    wire new_AGEMA_signal_8838 ;
    wire new_AGEMA_signal_8839 ;
    wire new_AGEMA_signal_8840 ;
    wire new_AGEMA_signal_8841 ;
    wire new_AGEMA_signal_8842 ;
    wire new_AGEMA_signal_8843 ;
    wire new_AGEMA_signal_8844 ;
    wire new_AGEMA_signal_8845 ;
    wire new_AGEMA_signal_8846 ;
    wire new_AGEMA_signal_8847 ;
    wire new_AGEMA_signal_8848 ;
    wire new_AGEMA_signal_8849 ;
    wire new_AGEMA_signal_8850 ;
    wire new_AGEMA_signal_8851 ;
    wire new_AGEMA_signal_8852 ;
    wire new_AGEMA_signal_8853 ;
    wire new_AGEMA_signal_8854 ;
    wire new_AGEMA_signal_8855 ;
    wire new_AGEMA_signal_8856 ;
    wire new_AGEMA_signal_8857 ;
    wire new_AGEMA_signal_8858 ;
    wire new_AGEMA_signal_8859 ;
    wire new_AGEMA_signal_8860 ;
    wire new_AGEMA_signal_8861 ;
    wire new_AGEMA_signal_8862 ;
    wire new_AGEMA_signal_8863 ;
    wire new_AGEMA_signal_8864 ;
    wire new_AGEMA_signal_8865 ;
    wire new_AGEMA_signal_8866 ;
    wire new_AGEMA_signal_8867 ;
    wire new_AGEMA_signal_8868 ;
    wire new_AGEMA_signal_8869 ;
    wire new_AGEMA_signal_8870 ;
    wire new_AGEMA_signal_8871 ;
    wire new_AGEMA_signal_8872 ;
    wire new_AGEMA_signal_8873 ;
    wire new_AGEMA_signal_8874 ;
    wire new_AGEMA_signal_8875 ;
    wire new_AGEMA_signal_8876 ;
    wire new_AGEMA_signal_8877 ;
    wire new_AGEMA_signal_8878 ;
    wire new_AGEMA_signal_8879 ;
    wire new_AGEMA_signal_8880 ;
    wire new_AGEMA_signal_8881 ;
    wire new_AGEMA_signal_8882 ;
    wire new_AGEMA_signal_8883 ;
    wire new_AGEMA_signal_8884 ;
    wire new_AGEMA_signal_8885 ;
    wire new_AGEMA_signal_8886 ;
    wire new_AGEMA_signal_8887 ;
    wire new_AGEMA_signal_8888 ;
    wire new_AGEMA_signal_8889 ;
    wire new_AGEMA_signal_8890 ;
    wire new_AGEMA_signal_8891 ;
    wire new_AGEMA_signal_8892 ;
    wire new_AGEMA_signal_8893 ;
    wire new_AGEMA_signal_8894 ;
    wire new_AGEMA_signal_8895 ;
    wire new_AGEMA_signal_8896 ;
    wire new_AGEMA_signal_8897 ;
    wire new_AGEMA_signal_8898 ;
    wire new_AGEMA_signal_8899 ;
    wire new_AGEMA_signal_8900 ;
    wire new_AGEMA_signal_8901 ;
    wire new_AGEMA_signal_8902 ;
    wire new_AGEMA_signal_8903 ;
    wire new_AGEMA_signal_8904 ;
    wire new_AGEMA_signal_8905 ;
    wire new_AGEMA_signal_8906 ;
    wire new_AGEMA_signal_8907 ;
    wire new_AGEMA_signal_8908 ;
    wire new_AGEMA_signal_8909 ;
    wire new_AGEMA_signal_8910 ;
    wire new_AGEMA_signal_8911 ;
    wire new_AGEMA_signal_8912 ;
    wire new_AGEMA_signal_8913 ;
    wire new_AGEMA_signal_8914 ;
    wire new_AGEMA_signal_8915 ;
    wire new_AGEMA_signal_8916 ;
    wire new_AGEMA_signal_8917 ;
    wire new_AGEMA_signal_8918 ;
    wire new_AGEMA_signal_8919 ;
    wire new_AGEMA_signal_8920 ;
    wire new_AGEMA_signal_8921 ;
    wire new_AGEMA_signal_8922 ;
    wire new_AGEMA_signal_8923 ;
    wire new_AGEMA_signal_8924 ;
    wire new_AGEMA_signal_8925 ;
    wire new_AGEMA_signal_8926 ;
    wire new_AGEMA_signal_8927 ;
    wire new_AGEMA_signal_8928 ;
    wire new_AGEMA_signal_8929 ;
    wire new_AGEMA_signal_8930 ;
    wire new_AGEMA_signal_8931 ;
    wire new_AGEMA_signal_8932 ;
    wire new_AGEMA_signal_8933 ;
    wire new_AGEMA_signal_8934 ;
    wire new_AGEMA_signal_8935 ;
    wire new_AGEMA_signal_8936 ;
    wire new_AGEMA_signal_8937 ;
    wire new_AGEMA_signal_8938 ;
    wire new_AGEMA_signal_8939 ;
    wire new_AGEMA_signal_8940 ;
    wire new_AGEMA_signal_8941 ;
    wire new_AGEMA_signal_8942 ;
    wire new_AGEMA_signal_8943 ;
    wire new_AGEMA_signal_8944 ;
    wire new_AGEMA_signal_8945 ;
    wire new_AGEMA_signal_8946 ;
    wire new_AGEMA_signal_8947 ;
    wire new_AGEMA_signal_8948 ;
    wire new_AGEMA_signal_8949 ;
    wire new_AGEMA_signal_8950 ;
    wire new_AGEMA_signal_8951 ;
    wire new_AGEMA_signal_8952 ;
    wire new_AGEMA_signal_8953 ;
    wire new_AGEMA_signal_8954 ;
    wire new_AGEMA_signal_8955 ;
    wire new_AGEMA_signal_8956 ;
    wire new_AGEMA_signal_8957 ;
    wire new_AGEMA_signal_8958 ;
    wire new_AGEMA_signal_8959 ;
    wire new_AGEMA_signal_8960 ;
    wire new_AGEMA_signal_8961 ;
    wire new_AGEMA_signal_8962 ;
    wire new_AGEMA_signal_8963 ;
    wire new_AGEMA_signal_8964 ;
    wire new_AGEMA_signal_8965 ;
    wire new_AGEMA_signal_8966 ;
    wire new_AGEMA_signal_8967 ;
    wire new_AGEMA_signal_8968 ;
    wire new_AGEMA_signal_8969 ;
    wire new_AGEMA_signal_8970 ;
    wire new_AGEMA_signal_8971 ;
    wire new_AGEMA_signal_8972 ;
    wire new_AGEMA_signal_8973 ;
    wire new_AGEMA_signal_8974 ;
    wire new_AGEMA_signal_8975 ;
    wire new_AGEMA_signal_8976 ;
    wire new_AGEMA_signal_8977 ;
    wire new_AGEMA_signal_8978 ;
    wire new_AGEMA_signal_8979 ;
    wire new_AGEMA_signal_8980 ;
    wire new_AGEMA_signal_8981 ;
    wire new_AGEMA_signal_8982 ;
    wire new_AGEMA_signal_8983 ;
    wire new_AGEMA_signal_8984 ;
    wire new_AGEMA_signal_8985 ;
    wire new_AGEMA_signal_8986 ;
    wire new_AGEMA_signal_8987 ;
    wire new_AGEMA_signal_8988 ;
    wire new_AGEMA_signal_8989 ;
    wire new_AGEMA_signal_8990 ;
    wire new_AGEMA_signal_8991 ;
    wire new_AGEMA_signal_8992 ;
    wire new_AGEMA_signal_8993 ;
    wire new_AGEMA_signal_8994 ;
    wire new_AGEMA_signal_8995 ;
    wire new_AGEMA_signal_8996 ;
    wire new_AGEMA_signal_8997 ;
    wire new_AGEMA_signal_8998 ;
    wire new_AGEMA_signal_8999 ;
    wire new_AGEMA_signal_9000 ;
    wire new_AGEMA_signal_9001 ;
    wire new_AGEMA_signal_9002 ;
    wire new_AGEMA_signal_9003 ;
    wire new_AGEMA_signal_9004 ;
    wire new_AGEMA_signal_9005 ;
    wire new_AGEMA_signal_9006 ;
    wire new_AGEMA_signal_9007 ;
    wire new_AGEMA_signal_9008 ;
    wire new_AGEMA_signal_9009 ;
    wire new_AGEMA_signal_9010 ;
    wire new_AGEMA_signal_9011 ;
    wire new_AGEMA_signal_9012 ;
    wire new_AGEMA_signal_9013 ;
    wire new_AGEMA_signal_9014 ;
    wire new_AGEMA_signal_9015 ;
    wire new_AGEMA_signal_9016 ;
    wire new_AGEMA_signal_9017 ;
    wire new_AGEMA_signal_9018 ;
    wire new_AGEMA_signal_9019 ;
    wire new_AGEMA_signal_9020 ;
    wire new_AGEMA_signal_9021 ;
    wire new_AGEMA_signal_9022 ;
    wire new_AGEMA_signal_9023 ;
    wire new_AGEMA_signal_9024 ;
    wire new_AGEMA_signal_9025 ;
    wire new_AGEMA_signal_9026 ;
    wire new_AGEMA_signal_9027 ;
    wire new_AGEMA_signal_9028 ;
    wire new_AGEMA_signal_9029 ;
    wire new_AGEMA_signal_9030 ;
    wire new_AGEMA_signal_9031 ;
    wire new_AGEMA_signal_9032 ;
    wire new_AGEMA_signal_9033 ;
    wire new_AGEMA_signal_9034 ;
    wire new_AGEMA_signal_9035 ;
    wire new_AGEMA_signal_9036 ;
    wire new_AGEMA_signal_9037 ;
    wire new_AGEMA_signal_9038 ;
    wire new_AGEMA_signal_9039 ;
    wire new_AGEMA_signal_9040 ;
    wire new_AGEMA_signal_9041 ;
    wire new_AGEMA_signal_9042 ;
    wire new_AGEMA_signal_9043 ;
    wire new_AGEMA_signal_9044 ;
    wire new_AGEMA_signal_9045 ;
    wire new_AGEMA_signal_9046 ;
    wire new_AGEMA_signal_9047 ;
    wire new_AGEMA_signal_9048 ;
    wire new_AGEMA_signal_9049 ;
    wire new_AGEMA_signal_9050 ;
    wire new_AGEMA_signal_9051 ;
    wire new_AGEMA_signal_9052 ;
    wire new_AGEMA_signal_9053 ;
    wire new_AGEMA_signal_9054 ;
    wire new_AGEMA_signal_9055 ;
    wire new_AGEMA_signal_9056 ;
    wire new_AGEMA_signal_9057 ;
    wire new_AGEMA_signal_9058 ;
    wire new_AGEMA_signal_9059 ;
    wire new_AGEMA_signal_9060 ;
    wire new_AGEMA_signal_9061 ;
    wire new_AGEMA_signal_9062 ;
    wire new_AGEMA_signal_9063 ;
    wire new_AGEMA_signal_9064 ;
    wire new_AGEMA_signal_9065 ;
    wire new_AGEMA_signal_9066 ;
    wire new_AGEMA_signal_9067 ;
    wire new_AGEMA_signal_9068 ;
    wire new_AGEMA_signal_9069 ;
    wire new_AGEMA_signal_9070 ;
    wire new_AGEMA_signal_9071 ;
    wire new_AGEMA_signal_9072 ;
    wire new_AGEMA_signal_9073 ;
    wire new_AGEMA_signal_9074 ;
    wire new_AGEMA_signal_9075 ;
    wire new_AGEMA_signal_9076 ;
    wire new_AGEMA_signal_9077 ;
    wire new_AGEMA_signal_9078 ;
    wire new_AGEMA_signal_9079 ;
    wire new_AGEMA_signal_9080 ;
    wire new_AGEMA_signal_9081 ;
    wire new_AGEMA_signal_9082 ;
    wire new_AGEMA_signal_9083 ;
    wire new_AGEMA_signal_9084 ;
    wire new_AGEMA_signal_9085 ;
    wire new_AGEMA_signal_9086 ;
    wire new_AGEMA_signal_9087 ;
    wire new_AGEMA_signal_9088 ;
    wire new_AGEMA_signal_9089 ;
    wire new_AGEMA_signal_9090 ;
    wire new_AGEMA_signal_9091 ;
    wire new_AGEMA_signal_9092 ;
    wire new_AGEMA_signal_9093 ;
    wire new_AGEMA_signal_9094 ;
    wire new_AGEMA_signal_9095 ;
    wire new_AGEMA_signal_9096 ;
    wire new_AGEMA_signal_9097 ;
    wire new_AGEMA_signal_9098 ;
    wire new_AGEMA_signal_9099 ;
    wire new_AGEMA_signal_9100 ;
    wire new_AGEMA_signal_9101 ;
    wire new_AGEMA_signal_9102 ;
    wire new_AGEMA_signal_9103 ;
    wire new_AGEMA_signal_9104 ;
    wire new_AGEMA_signal_9105 ;
    wire new_AGEMA_signal_9106 ;
    wire new_AGEMA_signal_9107 ;
    wire new_AGEMA_signal_9108 ;
    wire new_AGEMA_signal_9109 ;
    wire new_AGEMA_signal_9110 ;
    wire new_AGEMA_signal_9111 ;
    wire new_AGEMA_signal_9112 ;
    wire new_AGEMA_signal_9113 ;
    wire new_AGEMA_signal_9114 ;
    wire new_AGEMA_signal_9115 ;
    wire new_AGEMA_signal_9116 ;
    wire new_AGEMA_signal_9117 ;
    wire new_AGEMA_signal_9118 ;
    wire new_AGEMA_signal_9119 ;
    wire new_AGEMA_signal_9120 ;
    wire new_AGEMA_signal_9121 ;
    wire new_AGEMA_signal_9122 ;
    wire new_AGEMA_signal_9123 ;
    wire new_AGEMA_signal_9124 ;
    wire new_AGEMA_signal_9125 ;
    wire new_AGEMA_signal_9126 ;
    wire new_AGEMA_signal_9127 ;
    wire new_AGEMA_signal_9128 ;
    wire new_AGEMA_signal_9129 ;
    wire new_AGEMA_signal_9130 ;
    wire new_AGEMA_signal_9131 ;
    wire new_AGEMA_signal_9132 ;
    wire new_AGEMA_signal_9133 ;
    wire new_AGEMA_signal_9134 ;
    wire new_AGEMA_signal_9135 ;
    wire new_AGEMA_signal_9136 ;
    wire new_AGEMA_signal_9137 ;
    wire new_AGEMA_signal_9138 ;
    wire new_AGEMA_signal_9139 ;
    wire new_AGEMA_signal_9140 ;
    wire new_AGEMA_signal_9141 ;
    wire new_AGEMA_signal_9142 ;
    wire new_AGEMA_signal_9143 ;
    wire new_AGEMA_signal_9144 ;
    wire new_AGEMA_signal_9145 ;
    wire new_AGEMA_signal_9146 ;
    wire new_AGEMA_signal_9147 ;
    wire new_AGEMA_signal_9148 ;
    wire new_AGEMA_signal_9149 ;
    wire new_AGEMA_signal_9150 ;
    wire new_AGEMA_signal_9151 ;
    wire new_AGEMA_signal_9152 ;
    wire new_AGEMA_signal_9153 ;
    wire new_AGEMA_signal_9154 ;
    wire new_AGEMA_signal_9155 ;
    wire new_AGEMA_signal_9156 ;
    wire new_AGEMA_signal_9157 ;
    wire new_AGEMA_signal_9158 ;
    wire new_AGEMA_signal_9159 ;
    wire new_AGEMA_signal_9160 ;
    wire new_AGEMA_signal_9161 ;
    wire new_AGEMA_signal_9162 ;
    wire new_AGEMA_signal_9163 ;
    wire new_AGEMA_signal_9164 ;
    wire new_AGEMA_signal_9165 ;
    wire new_AGEMA_signal_9166 ;
    wire new_AGEMA_signal_9167 ;
    wire new_AGEMA_signal_9168 ;
    wire new_AGEMA_signal_9169 ;
    wire new_AGEMA_signal_9170 ;
    wire new_AGEMA_signal_9171 ;
    wire new_AGEMA_signal_9172 ;
    wire new_AGEMA_signal_9173 ;
    wire new_AGEMA_signal_9174 ;
    wire new_AGEMA_signal_9175 ;
    wire new_AGEMA_signal_9176 ;
    wire new_AGEMA_signal_9177 ;
    wire new_AGEMA_signal_9178 ;
    wire new_AGEMA_signal_9179 ;
    wire new_AGEMA_signal_9180 ;
    wire new_AGEMA_signal_9181 ;
    wire new_AGEMA_signal_9182 ;
    wire new_AGEMA_signal_9183 ;
    wire new_AGEMA_signal_9184 ;
    wire new_AGEMA_signal_9185 ;
    wire new_AGEMA_signal_9186 ;
    wire new_AGEMA_signal_9187 ;
    wire new_AGEMA_signal_9188 ;
    wire new_AGEMA_signal_9189 ;
    wire new_AGEMA_signal_9190 ;
    wire new_AGEMA_signal_9191 ;
    wire new_AGEMA_signal_9192 ;
    wire new_AGEMA_signal_9193 ;
    wire new_AGEMA_signal_9194 ;
    wire new_AGEMA_signal_9195 ;
    wire new_AGEMA_signal_9196 ;
    wire new_AGEMA_signal_9197 ;
    wire new_AGEMA_signal_9198 ;
    wire new_AGEMA_signal_9199 ;
    wire new_AGEMA_signal_9200 ;
    wire new_AGEMA_signal_9201 ;
    wire new_AGEMA_signal_9202 ;
    wire new_AGEMA_signal_9203 ;
    wire new_AGEMA_signal_9204 ;
    wire new_AGEMA_signal_9205 ;
    wire new_AGEMA_signal_9206 ;
    wire new_AGEMA_signal_9207 ;
    wire new_AGEMA_signal_9208 ;
    wire new_AGEMA_signal_9209 ;
    wire new_AGEMA_signal_9210 ;
    wire new_AGEMA_signal_9211 ;
    wire new_AGEMA_signal_9212 ;
    wire new_AGEMA_signal_9213 ;
    wire new_AGEMA_signal_9214 ;
    wire new_AGEMA_signal_9215 ;
    wire new_AGEMA_signal_9216 ;
    wire new_AGEMA_signal_9217 ;
    wire new_AGEMA_signal_9218 ;
    wire new_AGEMA_signal_9219 ;
    wire new_AGEMA_signal_9220 ;
    wire new_AGEMA_signal_9221 ;
    wire new_AGEMA_signal_9222 ;
    wire new_AGEMA_signal_9223 ;
    wire new_AGEMA_signal_9224 ;
    wire new_AGEMA_signal_9225 ;
    wire new_AGEMA_signal_9226 ;
    wire new_AGEMA_signal_9227 ;
    wire new_AGEMA_signal_9228 ;
    wire new_AGEMA_signal_9229 ;
    wire new_AGEMA_signal_9230 ;
    wire new_AGEMA_signal_9231 ;
    wire new_AGEMA_signal_9232 ;
    wire new_AGEMA_signal_9233 ;
    wire new_AGEMA_signal_9234 ;
    wire new_AGEMA_signal_9235 ;
    wire new_AGEMA_signal_9236 ;
    wire new_AGEMA_signal_9237 ;
    wire new_AGEMA_signal_9238 ;
    wire new_AGEMA_signal_9239 ;
    wire new_AGEMA_signal_9240 ;
    wire new_AGEMA_signal_9241 ;
    wire new_AGEMA_signal_9242 ;
    wire new_AGEMA_signal_9243 ;
    wire new_AGEMA_signal_9244 ;
    wire new_AGEMA_signal_9245 ;
    wire new_AGEMA_signal_9246 ;
    wire new_AGEMA_signal_9247 ;
    wire new_AGEMA_signal_9248 ;
    wire new_AGEMA_signal_9249 ;
    wire new_AGEMA_signal_9250 ;
    wire new_AGEMA_signal_9251 ;
    wire new_AGEMA_signal_9252 ;
    wire new_AGEMA_signal_9253 ;
    wire new_AGEMA_signal_9254 ;
    wire new_AGEMA_signal_9255 ;
    wire new_AGEMA_signal_9256 ;
    wire new_AGEMA_signal_9257 ;
    wire new_AGEMA_signal_9258 ;
    wire new_AGEMA_signal_9259 ;
    wire new_AGEMA_signal_9260 ;
    wire new_AGEMA_signal_9261 ;
    wire new_AGEMA_signal_9262 ;
    wire new_AGEMA_signal_9263 ;
    wire new_AGEMA_signal_9264 ;
    wire new_AGEMA_signal_9265 ;
    wire new_AGEMA_signal_9266 ;
    wire new_AGEMA_signal_9267 ;
    wire new_AGEMA_signal_9268 ;
    wire new_AGEMA_signal_9269 ;
    wire new_AGEMA_signal_9270 ;
    wire new_AGEMA_signal_9271 ;
    wire new_AGEMA_signal_9272 ;
    wire new_AGEMA_signal_9273 ;
    wire new_AGEMA_signal_9274 ;
    wire new_AGEMA_signal_9275 ;
    wire new_AGEMA_signal_9276 ;
    wire new_AGEMA_signal_9277 ;
    wire new_AGEMA_signal_9278 ;
    wire new_AGEMA_signal_9279 ;
    wire new_AGEMA_signal_9280 ;
    wire new_AGEMA_signal_9281 ;
    wire new_AGEMA_signal_9282 ;
    wire new_AGEMA_signal_9283 ;
    wire new_AGEMA_signal_9284 ;
    wire new_AGEMA_signal_9285 ;
    wire new_AGEMA_signal_9286 ;
    wire new_AGEMA_signal_9287 ;
    wire new_AGEMA_signal_9288 ;
    wire new_AGEMA_signal_9289 ;
    wire new_AGEMA_signal_9290 ;
    wire new_AGEMA_signal_9291 ;
    wire new_AGEMA_signal_9292 ;
    wire new_AGEMA_signal_9293 ;
    wire new_AGEMA_signal_9294 ;
    wire new_AGEMA_signal_9295 ;
    wire new_AGEMA_signal_9296 ;
    wire new_AGEMA_signal_9297 ;
    wire new_AGEMA_signal_9298 ;
    wire new_AGEMA_signal_9299 ;
    wire new_AGEMA_signal_9300 ;
    wire new_AGEMA_signal_9301 ;
    wire new_AGEMA_signal_9302 ;
    wire new_AGEMA_signal_9303 ;
    wire new_AGEMA_signal_9304 ;
    wire new_AGEMA_signal_9305 ;
    wire new_AGEMA_signal_9306 ;
    wire new_AGEMA_signal_9307 ;
    wire new_AGEMA_signal_9308 ;
    wire new_AGEMA_signal_9309 ;
    wire new_AGEMA_signal_9310 ;
    wire new_AGEMA_signal_9311 ;
    wire new_AGEMA_signal_9312 ;
    wire new_AGEMA_signal_9313 ;
    wire new_AGEMA_signal_9314 ;
    wire new_AGEMA_signal_9315 ;
    wire new_AGEMA_signal_9316 ;
    wire new_AGEMA_signal_9317 ;
    wire new_AGEMA_signal_9318 ;
    wire new_AGEMA_signal_9319 ;
    wire new_AGEMA_signal_9320 ;
    wire new_AGEMA_signal_9321 ;
    wire new_AGEMA_signal_9322 ;
    wire new_AGEMA_signal_9323 ;
    wire new_AGEMA_signal_9324 ;
    wire new_AGEMA_signal_9325 ;
    wire new_AGEMA_signal_9326 ;
    wire new_AGEMA_signal_9327 ;
    wire new_AGEMA_signal_9328 ;
    wire new_AGEMA_signal_9329 ;
    wire new_AGEMA_signal_9330 ;
    wire new_AGEMA_signal_9331 ;
    wire new_AGEMA_signal_9332 ;
    wire new_AGEMA_signal_9333 ;
    wire new_AGEMA_signal_9334 ;
    wire new_AGEMA_signal_9335 ;
    wire new_AGEMA_signal_9336 ;
    wire new_AGEMA_signal_9337 ;
    wire new_AGEMA_signal_9338 ;
    wire new_AGEMA_signal_9339 ;
    wire new_AGEMA_signal_9340 ;
    wire new_AGEMA_signal_9341 ;
    wire new_AGEMA_signal_9342 ;
    wire new_AGEMA_signal_9343 ;
    wire new_AGEMA_signal_9344 ;
    wire new_AGEMA_signal_9345 ;
    wire new_AGEMA_signal_9346 ;
    wire new_AGEMA_signal_9347 ;
    wire new_AGEMA_signal_9348 ;
    wire new_AGEMA_signal_9349 ;
    wire new_AGEMA_signal_9350 ;
    wire new_AGEMA_signal_9351 ;
    wire new_AGEMA_signal_9352 ;
    wire new_AGEMA_signal_9353 ;
    wire new_AGEMA_signal_9354 ;
    wire new_AGEMA_signal_9355 ;
    wire new_AGEMA_signal_9356 ;
    wire new_AGEMA_signal_9357 ;
    wire new_AGEMA_signal_9358 ;
    wire new_AGEMA_signal_9359 ;
    wire new_AGEMA_signal_9360 ;
    wire new_AGEMA_signal_9361 ;
    wire new_AGEMA_signal_9362 ;
    wire new_AGEMA_signal_9363 ;
    wire new_AGEMA_signal_9364 ;
    wire new_AGEMA_signal_9365 ;
    wire new_AGEMA_signal_9366 ;
    wire new_AGEMA_signal_9367 ;
    wire new_AGEMA_signal_9368 ;
    wire new_AGEMA_signal_9369 ;
    wire new_AGEMA_signal_9370 ;
    wire new_AGEMA_signal_9371 ;
    wire new_AGEMA_signal_9372 ;
    wire new_AGEMA_signal_9373 ;
    wire new_AGEMA_signal_9374 ;
    wire new_AGEMA_signal_9375 ;
    wire new_AGEMA_signal_9376 ;
    wire new_AGEMA_signal_9377 ;
    wire new_AGEMA_signal_9378 ;
    wire new_AGEMA_signal_9379 ;
    wire new_AGEMA_signal_9380 ;
    wire new_AGEMA_signal_9381 ;
    wire new_AGEMA_signal_9382 ;
    wire new_AGEMA_signal_9383 ;
    wire new_AGEMA_signal_9384 ;
    wire new_AGEMA_signal_9385 ;
    wire new_AGEMA_signal_9386 ;
    wire new_AGEMA_signal_9387 ;
    wire new_AGEMA_signal_9388 ;
    wire new_AGEMA_signal_9389 ;
    wire new_AGEMA_signal_9390 ;
    wire new_AGEMA_signal_9391 ;
    wire new_AGEMA_signal_9392 ;
    wire new_AGEMA_signal_9393 ;
    wire new_AGEMA_signal_9394 ;
    wire new_AGEMA_signal_9395 ;
    wire new_AGEMA_signal_9396 ;
    wire new_AGEMA_signal_9397 ;
    wire new_AGEMA_signal_9398 ;
    wire new_AGEMA_signal_9399 ;
    wire new_AGEMA_signal_9400 ;
    wire new_AGEMA_signal_9401 ;
    wire new_AGEMA_signal_9402 ;
    wire new_AGEMA_signal_9403 ;
    wire new_AGEMA_signal_9404 ;
    wire new_AGEMA_signal_9405 ;
    wire new_AGEMA_signal_9406 ;
    wire new_AGEMA_signal_9407 ;
    wire new_AGEMA_signal_9408 ;
    wire new_AGEMA_signal_9409 ;
    wire new_AGEMA_signal_9410 ;
    wire new_AGEMA_signal_9411 ;
    wire new_AGEMA_signal_9412 ;
    wire new_AGEMA_signal_9413 ;
    wire new_AGEMA_signal_9414 ;
    wire new_AGEMA_signal_9415 ;
    wire new_AGEMA_signal_9416 ;
    wire new_AGEMA_signal_9417 ;
    wire new_AGEMA_signal_9418 ;
    wire new_AGEMA_signal_9419 ;
    wire new_AGEMA_signal_9420 ;
    wire new_AGEMA_signal_9421 ;
    wire new_AGEMA_signal_9422 ;
    wire new_AGEMA_signal_9423 ;
    wire new_AGEMA_signal_9424 ;
    wire new_AGEMA_signal_9425 ;
    wire new_AGEMA_signal_9426 ;
    wire new_AGEMA_signal_9427 ;
    wire new_AGEMA_signal_9428 ;
    wire new_AGEMA_signal_9429 ;
    wire new_AGEMA_signal_9430 ;
    wire new_AGEMA_signal_9431 ;
    wire new_AGEMA_signal_9432 ;
    wire new_AGEMA_signal_9433 ;
    wire new_AGEMA_signal_9434 ;
    wire new_AGEMA_signal_9435 ;
    wire new_AGEMA_signal_9436 ;
    wire new_AGEMA_signal_9437 ;
    wire new_AGEMA_signal_9438 ;
    wire new_AGEMA_signal_9439 ;
    wire new_AGEMA_signal_9440 ;
    wire new_AGEMA_signal_9441 ;
    wire new_AGEMA_signal_9442 ;
    wire new_AGEMA_signal_9443 ;
    wire new_AGEMA_signal_9444 ;
    wire new_AGEMA_signal_9445 ;
    wire new_AGEMA_signal_9446 ;
    wire new_AGEMA_signal_9447 ;
    wire new_AGEMA_signal_9448 ;
    wire new_AGEMA_signal_9449 ;
    wire new_AGEMA_signal_9450 ;
    wire new_AGEMA_signal_9451 ;
    wire new_AGEMA_signal_9452 ;
    wire new_AGEMA_signal_9453 ;
    wire new_AGEMA_signal_9454 ;
    wire new_AGEMA_signal_9455 ;
    wire new_AGEMA_signal_9456 ;
    wire new_AGEMA_signal_9457 ;
    wire new_AGEMA_signal_9458 ;
    wire new_AGEMA_signal_9459 ;
    wire new_AGEMA_signal_9460 ;
    wire new_AGEMA_signal_9461 ;
    wire new_AGEMA_signal_9462 ;
    wire new_AGEMA_signal_9463 ;
    wire new_AGEMA_signal_9464 ;
    wire new_AGEMA_signal_9465 ;
    wire new_AGEMA_signal_9466 ;
    wire new_AGEMA_signal_9467 ;
    wire new_AGEMA_signal_9468 ;
    wire new_AGEMA_signal_9469 ;
    wire new_AGEMA_signal_9470 ;
    wire new_AGEMA_signal_9471 ;
    wire new_AGEMA_signal_9472 ;
    wire new_AGEMA_signal_9473 ;
    wire new_AGEMA_signal_9474 ;
    wire new_AGEMA_signal_9475 ;
    wire new_AGEMA_signal_9476 ;
    wire new_AGEMA_signal_9477 ;
    wire new_AGEMA_signal_9478 ;
    wire new_AGEMA_signal_9479 ;
    wire new_AGEMA_signal_9480 ;
    wire new_AGEMA_signal_9481 ;
    wire new_AGEMA_signal_9482 ;
    wire new_AGEMA_signal_9483 ;
    wire new_AGEMA_signal_9484 ;
    wire new_AGEMA_signal_9485 ;
    wire new_AGEMA_signal_9486 ;
    wire new_AGEMA_signal_9487 ;
    wire new_AGEMA_signal_9488 ;
    wire new_AGEMA_signal_9489 ;
    wire new_AGEMA_signal_9490 ;
    wire new_AGEMA_signal_9491 ;
    wire new_AGEMA_signal_9492 ;
    wire new_AGEMA_signal_9493 ;
    wire new_AGEMA_signal_9494 ;
    wire new_AGEMA_signal_9495 ;
    wire new_AGEMA_signal_9496 ;
    wire new_AGEMA_signal_9497 ;
    wire new_AGEMA_signal_9498 ;
    wire new_AGEMA_signal_9499 ;
    wire new_AGEMA_signal_9500 ;
    wire new_AGEMA_signal_9501 ;
    wire new_AGEMA_signal_9502 ;
    wire new_AGEMA_signal_9503 ;
    wire new_AGEMA_signal_9504 ;
    wire new_AGEMA_signal_9505 ;
    wire new_AGEMA_signal_9506 ;
    wire new_AGEMA_signal_9507 ;
    wire new_AGEMA_signal_9508 ;
    wire new_AGEMA_signal_9509 ;
    wire new_AGEMA_signal_9510 ;
    wire new_AGEMA_signal_9511 ;
    wire new_AGEMA_signal_9512 ;
    wire new_AGEMA_signal_9513 ;
    wire new_AGEMA_signal_9514 ;
    wire new_AGEMA_signal_9515 ;
    wire new_AGEMA_signal_9516 ;
    wire new_AGEMA_signal_9517 ;
    wire new_AGEMA_signal_9518 ;
    wire new_AGEMA_signal_9519 ;
    wire new_AGEMA_signal_9520 ;
    wire new_AGEMA_signal_9521 ;
    wire new_AGEMA_signal_9522 ;
    wire new_AGEMA_signal_9523 ;
    wire new_AGEMA_signal_9524 ;
    wire new_AGEMA_signal_9525 ;
    wire new_AGEMA_signal_9526 ;
    wire new_AGEMA_signal_9527 ;
    wire new_AGEMA_signal_9528 ;
    wire new_AGEMA_signal_9529 ;
    wire new_AGEMA_signal_9530 ;
    wire new_AGEMA_signal_9531 ;
    wire new_AGEMA_signal_9532 ;
    wire new_AGEMA_signal_9533 ;
    wire new_AGEMA_signal_9534 ;
    wire new_AGEMA_signal_9535 ;
    wire new_AGEMA_signal_9536 ;
    wire new_AGEMA_signal_9537 ;
    wire new_AGEMA_signal_9538 ;
    wire new_AGEMA_signal_9539 ;
    wire new_AGEMA_signal_9540 ;
    wire new_AGEMA_signal_9541 ;
    wire new_AGEMA_signal_9542 ;
    wire new_AGEMA_signal_9543 ;
    wire new_AGEMA_signal_9544 ;
    wire new_AGEMA_signal_9545 ;
    wire new_AGEMA_signal_9546 ;
    wire new_AGEMA_signal_9547 ;
    wire new_AGEMA_signal_9548 ;
    wire new_AGEMA_signal_9549 ;
    wire new_AGEMA_signal_9550 ;
    wire new_AGEMA_signal_9551 ;
    wire new_AGEMA_signal_9552 ;
    wire new_AGEMA_signal_9553 ;
    wire new_AGEMA_signal_9554 ;
    wire new_AGEMA_signal_9555 ;
    wire new_AGEMA_signal_9556 ;
    wire new_AGEMA_signal_9557 ;
    wire new_AGEMA_signal_9558 ;
    wire new_AGEMA_signal_9559 ;
    wire new_AGEMA_signal_9560 ;
    wire new_AGEMA_signal_9561 ;
    wire new_AGEMA_signal_9562 ;
    wire new_AGEMA_signal_9563 ;
    wire new_AGEMA_signal_9564 ;
    wire new_AGEMA_signal_9565 ;
    wire new_AGEMA_signal_9566 ;
    wire new_AGEMA_signal_9567 ;
    wire new_AGEMA_signal_9568 ;
    wire new_AGEMA_signal_9569 ;
    wire new_AGEMA_signal_9570 ;
    wire new_AGEMA_signal_9571 ;
    wire new_AGEMA_signal_9572 ;
    wire new_AGEMA_signal_9573 ;
    wire new_AGEMA_signal_9574 ;
    wire new_AGEMA_signal_9575 ;
    wire new_AGEMA_signal_9576 ;
    wire new_AGEMA_signal_9577 ;
    wire new_AGEMA_signal_9578 ;
    wire new_AGEMA_signal_9579 ;
    wire new_AGEMA_signal_9580 ;
    wire new_AGEMA_signal_9581 ;
    wire new_AGEMA_signal_9582 ;
    wire new_AGEMA_signal_9583 ;
    wire new_AGEMA_signal_9584 ;
    wire new_AGEMA_signal_9585 ;
    wire new_AGEMA_signal_9586 ;
    wire new_AGEMA_signal_9587 ;
    wire new_AGEMA_signal_9588 ;
    wire new_AGEMA_signal_9589 ;
    wire new_AGEMA_signal_9590 ;
    wire new_AGEMA_signal_9591 ;
    wire new_AGEMA_signal_9592 ;
    wire new_AGEMA_signal_9593 ;
    wire new_AGEMA_signal_9594 ;
    wire new_AGEMA_signal_9595 ;
    wire new_AGEMA_signal_9596 ;
    wire new_AGEMA_signal_9597 ;
    wire new_AGEMA_signal_9598 ;
    wire new_AGEMA_signal_9599 ;
    wire new_AGEMA_signal_9600 ;
    wire new_AGEMA_signal_9601 ;
    wire new_AGEMA_signal_9602 ;
    wire new_AGEMA_signal_9603 ;
    wire new_AGEMA_signal_9604 ;
    wire new_AGEMA_signal_9605 ;
    wire new_AGEMA_signal_9606 ;
    wire new_AGEMA_signal_9607 ;
    wire new_AGEMA_signal_9608 ;
    wire new_AGEMA_signal_9609 ;
    wire new_AGEMA_signal_9610 ;
    wire new_AGEMA_signal_9611 ;
    wire new_AGEMA_signal_9612 ;
    wire new_AGEMA_signal_9613 ;
    wire new_AGEMA_signal_9614 ;
    wire new_AGEMA_signal_9615 ;
    wire new_AGEMA_signal_9616 ;
    wire new_AGEMA_signal_9617 ;
    wire new_AGEMA_signal_9618 ;
    wire new_AGEMA_signal_9619 ;
    wire new_AGEMA_signal_9620 ;
    wire new_AGEMA_signal_9621 ;
    wire new_AGEMA_signal_9622 ;
    wire new_AGEMA_signal_9623 ;
    wire new_AGEMA_signal_9624 ;
    wire new_AGEMA_signal_9625 ;
    wire new_AGEMA_signal_9626 ;
    wire new_AGEMA_signal_9627 ;
    wire new_AGEMA_signal_9628 ;
    wire new_AGEMA_signal_9629 ;
    wire new_AGEMA_signal_9630 ;
    wire new_AGEMA_signal_9631 ;
    wire new_AGEMA_signal_9632 ;
    wire new_AGEMA_signal_9633 ;
    wire new_AGEMA_signal_9634 ;
    wire new_AGEMA_signal_9635 ;
    wire new_AGEMA_signal_9636 ;
    wire new_AGEMA_signal_9637 ;
    wire new_AGEMA_signal_9638 ;
    wire new_AGEMA_signal_9639 ;
    wire new_AGEMA_signal_9640 ;
    wire new_AGEMA_signal_9641 ;
    wire new_AGEMA_signal_9642 ;
    wire new_AGEMA_signal_9643 ;
    wire new_AGEMA_signal_9644 ;
    wire new_AGEMA_signal_9645 ;
    wire new_AGEMA_signal_9646 ;
    wire new_AGEMA_signal_9647 ;
    wire new_AGEMA_signal_9648 ;
    wire new_AGEMA_signal_9649 ;
    wire new_AGEMA_signal_9650 ;
    wire new_AGEMA_signal_9651 ;
    wire new_AGEMA_signal_9652 ;
    wire new_AGEMA_signal_9653 ;
    wire new_AGEMA_signal_9654 ;
    wire new_AGEMA_signal_9655 ;
    wire new_AGEMA_signal_9656 ;
    wire new_AGEMA_signal_9657 ;
    wire new_AGEMA_signal_9658 ;
    wire new_AGEMA_signal_9659 ;
    wire new_AGEMA_signal_9660 ;
    wire new_AGEMA_signal_9661 ;
    wire new_AGEMA_signal_9662 ;
    wire new_AGEMA_signal_9663 ;
    wire new_AGEMA_signal_9664 ;
    wire new_AGEMA_signal_9665 ;
    wire new_AGEMA_signal_9666 ;
    wire new_AGEMA_signal_9667 ;
    wire new_AGEMA_signal_9668 ;
    wire new_AGEMA_signal_9669 ;
    wire new_AGEMA_signal_9670 ;
    wire new_AGEMA_signal_9671 ;
    wire new_AGEMA_signal_9672 ;
    wire new_AGEMA_signal_9673 ;
    wire new_AGEMA_signal_9674 ;
    wire new_AGEMA_signal_9675 ;
    wire new_AGEMA_signal_9676 ;
    wire new_AGEMA_signal_9677 ;
    wire new_AGEMA_signal_9678 ;
    wire new_AGEMA_signal_9679 ;
    wire new_AGEMA_signal_9680 ;
    wire new_AGEMA_signal_9681 ;
    wire new_AGEMA_signal_9682 ;
    wire new_AGEMA_signal_9683 ;
    wire new_AGEMA_signal_9684 ;
    wire new_AGEMA_signal_9685 ;
    wire new_AGEMA_signal_9686 ;
    wire new_AGEMA_signal_9687 ;
    wire new_AGEMA_signal_9688 ;
    wire new_AGEMA_signal_9689 ;
    wire new_AGEMA_signal_9690 ;
    wire new_AGEMA_signal_9691 ;
    wire new_AGEMA_signal_9692 ;
    wire new_AGEMA_signal_9693 ;
    wire new_AGEMA_signal_9694 ;
    wire new_AGEMA_signal_9695 ;
    wire new_AGEMA_signal_9696 ;
    wire new_AGEMA_signal_9697 ;
    wire new_AGEMA_signal_9698 ;
    wire new_AGEMA_signal_9699 ;
    wire new_AGEMA_signal_9700 ;
    wire new_AGEMA_signal_9701 ;
    wire new_AGEMA_signal_9702 ;
    wire new_AGEMA_signal_9703 ;
    wire new_AGEMA_signal_9704 ;
    wire new_AGEMA_signal_9705 ;
    wire new_AGEMA_signal_9706 ;
    wire new_AGEMA_signal_9707 ;
    wire new_AGEMA_signal_9708 ;
    wire new_AGEMA_signal_9709 ;
    wire new_AGEMA_signal_9710 ;
    wire new_AGEMA_signal_9711 ;
    wire new_AGEMA_signal_9712 ;
    wire new_AGEMA_signal_9713 ;
    wire new_AGEMA_signal_9714 ;
    wire new_AGEMA_signal_9715 ;
    wire new_AGEMA_signal_9716 ;
    wire new_AGEMA_signal_9717 ;
    wire new_AGEMA_signal_9718 ;
    wire new_AGEMA_signal_9719 ;
    wire new_AGEMA_signal_9720 ;
    wire new_AGEMA_signal_9721 ;
    wire new_AGEMA_signal_9722 ;
    wire new_AGEMA_signal_9723 ;
    wire new_AGEMA_signal_9724 ;
    wire new_AGEMA_signal_9725 ;
    wire new_AGEMA_signal_9726 ;
    wire new_AGEMA_signal_9727 ;
    wire new_AGEMA_signal_9728 ;
    wire new_AGEMA_signal_9729 ;
    wire new_AGEMA_signal_9730 ;
    wire new_AGEMA_signal_9731 ;
    wire new_AGEMA_signal_9732 ;
    wire new_AGEMA_signal_9733 ;
    wire new_AGEMA_signal_9734 ;
    wire new_AGEMA_signal_9735 ;
    wire new_AGEMA_signal_9736 ;
    wire new_AGEMA_signal_9737 ;
    wire new_AGEMA_signal_9738 ;
    wire new_AGEMA_signal_9739 ;
    wire new_AGEMA_signal_9740 ;
    wire new_AGEMA_signal_9741 ;
    wire new_AGEMA_signal_9742 ;
    wire new_AGEMA_signal_9743 ;
    wire new_AGEMA_signal_9744 ;
    wire new_AGEMA_signal_9745 ;
    wire new_AGEMA_signal_9746 ;
    wire new_AGEMA_signal_9747 ;
    wire new_AGEMA_signal_9748 ;
    wire new_AGEMA_signal_9749 ;
    wire new_AGEMA_signal_9750 ;
    wire new_AGEMA_signal_9751 ;
    wire new_AGEMA_signal_9752 ;
    wire new_AGEMA_signal_9753 ;
    wire new_AGEMA_signal_9754 ;
    wire new_AGEMA_signal_9755 ;
    wire new_AGEMA_signal_9756 ;
    wire new_AGEMA_signal_9757 ;
    wire new_AGEMA_signal_9758 ;
    wire new_AGEMA_signal_9759 ;
    wire new_AGEMA_signal_9760 ;
    wire new_AGEMA_signal_9761 ;
    wire new_AGEMA_signal_9762 ;
    wire new_AGEMA_signal_9763 ;
    wire new_AGEMA_signal_9764 ;
    wire new_AGEMA_signal_9765 ;
    wire new_AGEMA_signal_9766 ;
    wire new_AGEMA_signal_9767 ;
    wire new_AGEMA_signal_9768 ;
    wire new_AGEMA_signal_9769 ;
    wire new_AGEMA_signal_9770 ;
    wire new_AGEMA_signal_9771 ;
    wire new_AGEMA_signal_9772 ;
    wire new_AGEMA_signal_9773 ;
    wire new_AGEMA_signal_9774 ;
    wire new_AGEMA_signal_9775 ;
    wire new_AGEMA_signal_9776 ;
    wire new_AGEMA_signal_9777 ;
    wire new_AGEMA_signal_9778 ;
    wire new_AGEMA_signal_9779 ;
    wire new_AGEMA_signal_9780 ;
    wire new_AGEMA_signal_9781 ;
    wire new_AGEMA_signal_9782 ;
    wire new_AGEMA_signal_9783 ;
    wire new_AGEMA_signal_9784 ;
    wire new_AGEMA_signal_9785 ;
    wire new_AGEMA_signal_9786 ;
    wire new_AGEMA_signal_9787 ;
    wire new_AGEMA_signal_9788 ;
    wire new_AGEMA_signal_9789 ;
    wire new_AGEMA_signal_9790 ;
    wire new_AGEMA_signal_9791 ;
    wire new_AGEMA_signal_9792 ;
    wire new_AGEMA_signal_9793 ;
    wire new_AGEMA_signal_9794 ;
    wire new_AGEMA_signal_9795 ;
    wire new_AGEMA_signal_9796 ;
    wire new_AGEMA_signal_9797 ;
    wire new_AGEMA_signal_9798 ;
    wire new_AGEMA_signal_9799 ;
    wire new_AGEMA_signal_9800 ;
    wire new_AGEMA_signal_9801 ;
    wire new_AGEMA_signal_9802 ;
    wire new_AGEMA_signal_9803 ;
    wire new_AGEMA_signal_9804 ;
    wire new_AGEMA_signal_9805 ;
    wire new_AGEMA_signal_9806 ;
    wire new_AGEMA_signal_9807 ;
    wire new_AGEMA_signal_9808 ;
    wire new_AGEMA_signal_9809 ;
    wire new_AGEMA_signal_9810 ;
    wire new_AGEMA_signal_9811 ;
    wire new_AGEMA_signal_9812 ;
    wire new_AGEMA_signal_9813 ;
    wire new_AGEMA_signal_9814 ;
    wire new_AGEMA_signal_9815 ;
    wire new_AGEMA_signal_9816 ;
    wire new_AGEMA_signal_9817 ;
    wire new_AGEMA_signal_9818 ;
    wire new_AGEMA_signal_9819 ;
    wire new_AGEMA_signal_9820 ;
    wire new_AGEMA_signal_9821 ;
    wire new_AGEMA_signal_9822 ;
    wire new_AGEMA_signal_9823 ;
    wire new_AGEMA_signal_9824 ;
    wire new_AGEMA_signal_9825 ;
    wire new_AGEMA_signal_9826 ;
    wire new_AGEMA_signal_9827 ;
    wire new_AGEMA_signal_9828 ;
    wire new_AGEMA_signal_9829 ;
    wire new_AGEMA_signal_9830 ;
    wire new_AGEMA_signal_9831 ;
    wire new_AGEMA_signal_9832 ;
    wire new_AGEMA_signal_9833 ;
    wire new_AGEMA_signal_9834 ;
    wire new_AGEMA_signal_9835 ;
    wire new_AGEMA_signal_9836 ;
    wire new_AGEMA_signal_9837 ;
    wire new_AGEMA_signal_9838 ;
    wire new_AGEMA_signal_9839 ;
    wire new_AGEMA_signal_9840 ;
    wire new_AGEMA_signal_9841 ;
    wire new_AGEMA_signal_9842 ;
    wire new_AGEMA_signal_9843 ;
    wire new_AGEMA_signal_9844 ;
    wire new_AGEMA_signal_9845 ;
    wire new_AGEMA_signal_9846 ;
    wire new_AGEMA_signal_9847 ;
    wire new_AGEMA_signal_9848 ;
    wire new_AGEMA_signal_9849 ;
    wire new_AGEMA_signal_9850 ;
    wire new_AGEMA_signal_9851 ;
    wire new_AGEMA_signal_9852 ;
    wire new_AGEMA_signal_9853 ;
    wire new_AGEMA_signal_9854 ;
    wire new_AGEMA_signal_9855 ;
    wire new_AGEMA_signal_9856 ;
    wire new_AGEMA_signal_9857 ;
    wire new_AGEMA_signal_9858 ;
    wire new_AGEMA_signal_9859 ;
    wire new_AGEMA_signal_9860 ;
    wire new_AGEMA_signal_9861 ;
    wire new_AGEMA_signal_9862 ;
    wire new_AGEMA_signal_9863 ;
    wire new_AGEMA_signal_9864 ;
    wire new_AGEMA_signal_9865 ;
    wire new_AGEMA_signal_9866 ;
    wire new_AGEMA_signal_9867 ;
    wire new_AGEMA_signal_9868 ;
    wire new_AGEMA_signal_9869 ;
    wire new_AGEMA_signal_9870 ;
    wire new_AGEMA_signal_9871 ;
    wire new_AGEMA_signal_9872 ;
    wire new_AGEMA_signal_9873 ;
    wire new_AGEMA_signal_9874 ;
    wire new_AGEMA_signal_9875 ;
    wire new_AGEMA_signal_9876 ;
    wire new_AGEMA_signal_9877 ;
    wire new_AGEMA_signal_9878 ;
    wire new_AGEMA_signal_9879 ;
    wire new_AGEMA_signal_9880 ;
    wire new_AGEMA_signal_9881 ;
    wire new_AGEMA_signal_9882 ;
    wire new_AGEMA_signal_9883 ;
    wire new_AGEMA_signal_9884 ;
    wire new_AGEMA_signal_9885 ;
    wire new_AGEMA_signal_9886 ;
    wire new_AGEMA_signal_9887 ;
    wire new_AGEMA_signal_9888 ;
    wire new_AGEMA_signal_9889 ;
    wire new_AGEMA_signal_9890 ;
    wire new_AGEMA_signal_9891 ;
    wire new_AGEMA_signal_9892 ;
    wire new_AGEMA_signal_9893 ;
    wire new_AGEMA_signal_9894 ;
    wire new_AGEMA_signal_9895 ;
    wire new_AGEMA_signal_9896 ;
    wire new_AGEMA_signal_9897 ;
    wire new_AGEMA_signal_9898 ;
    wire new_AGEMA_signal_9899 ;
    wire new_AGEMA_signal_9900 ;
    wire new_AGEMA_signal_9901 ;
    wire new_AGEMA_signal_9902 ;
    wire new_AGEMA_signal_9903 ;
    wire new_AGEMA_signal_9904 ;
    wire new_AGEMA_signal_9905 ;
    wire new_AGEMA_signal_9906 ;
    wire new_AGEMA_signal_9907 ;
    wire new_AGEMA_signal_9908 ;
    wire new_AGEMA_signal_9909 ;
    wire new_AGEMA_signal_9910 ;
    wire new_AGEMA_signal_9911 ;
    wire new_AGEMA_signal_9912 ;
    wire new_AGEMA_signal_9913 ;
    wire new_AGEMA_signal_9914 ;
    wire new_AGEMA_signal_9915 ;
    wire new_AGEMA_signal_9916 ;
    wire new_AGEMA_signal_9917 ;
    wire new_AGEMA_signal_9918 ;
    wire new_AGEMA_signal_9919 ;
    wire new_AGEMA_signal_9920 ;
    wire new_AGEMA_signal_9921 ;
    wire new_AGEMA_signal_9922 ;
    wire new_AGEMA_signal_9923 ;
    wire new_AGEMA_signal_9924 ;
    wire new_AGEMA_signal_9925 ;
    wire new_AGEMA_signal_9926 ;
    wire new_AGEMA_signal_9927 ;
    wire new_AGEMA_signal_9928 ;
    wire new_AGEMA_signal_9929 ;
    wire new_AGEMA_signal_9930 ;
    wire new_AGEMA_signal_9931 ;
    wire new_AGEMA_signal_9932 ;
    wire new_AGEMA_signal_9933 ;
    wire new_AGEMA_signal_9934 ;
    wire new_AGEMA_signal_9935 ;
    wire new_AGEMA_signal_9936 ;
    wire new_AGEMA_signal_9937 ;
    wire new_AGEMA_signal_9938 ;
    wire new_AGEMA_signal_9939 ;
    wire new_AGEMA_signal_9940 ;
    wire new_AGEMA_signal_9941 ;
    wire new_AGEMA_signal_9942 ;
    wire new_AGEMA_signal_9943 ;
    wire new_AGEMA_signal_9944 ;
    wire new_AGEMA_signal_9945 ;
    wire new_AGEMA_signal_9946 ;
    wire new_AGEMA_signal_9947 ;
    wire new_AGEMA_signal_9948 ;
    wire new_AGEMA_signal_9949 ;
    wire new_AGEMA_signal_9950 ;
    wire new_AGEMA_signal_9951 ;
    wire new_AGEMA_signal_9952 ;
    wire new_AGEMA_signal_9953 ;
    wire new_AGEMA_signal_9954 ;
    wire new_AGEMA_signal_9955 ;
    wire new_AGEMA_signal_9956 ;
    wire new_AGEMA_signal_9957 ;
    wire new_AGEMA_signal_9958 ;
    wire new_AGEMA_signal_9959 ;
    wire new_AGEMA_signal_9960 ;
    wire new_AGEMA_signal_9961 ;
    wire new_AGEMA_signal_9962 ;
    wire new_AGEMA_signal_9963 ;
    wire new_AGEMA_signal_9964 ;
    wire new_AGEMA_signal_9965 ;
    wire new_AGEMA_signal_9966 ;
    wire new_AGEMA_signal_9967 ;
    wire new_AGEMA_signal_9968 ;
    wire new_AGEMA_signal_9969 ;
    wire new_AGEMA_signal_9970 ;
    wire new_AGEMA_signal_9971 ;
    wire new_AGEMA_signal_9972 ;
    wire new_AGEMA_signal_9973 ;
    wire new_AGEMA_signal_9974 ;
    wire new_AGEMA_signal_9975 ;
    wire new_AGEMA_signal_9976 ;
    wire new_AGEMA_signal_9977 ;
    wire new_AGEMA_signal_9978 ;
    wire new_AGEMA_signal_9979 ;
    wire new_AGEMA_signal_9980 ;
    wire new_AGEMA_signal_9981 ;
    wire new_AGEMA_signal_9982 ;
    wire new_AGEMA_signal_9983 ;
    wire new_AGEMA_signal_9984 ;
    wire new_AGEMA_signal_9985 ;
    wire new_AGEMA_signal_9986 ;
    wire new_AGEMA_signal_9987 ;
    wire new_AGEMA_signal_9988 ;
    wire new_AGEMA_signal_9989 ;
    wire new_AGEMA_signal_9990 ;
    wire new_AGEMA_signal_9991 ;
    wire new_AGEMA_signal_9992 ;
    wire new_AGEMA_signal_9993 ;
    wire new_AGEMA_signal_9994 ;
    wire new_AGEMA_signal_9995 ;
    wire new_AGEMA_signal_9996 ;
    wire new_AGEMA_signal_9997 ;
    wire new_AGEMA_signal_9998 ;
    wire new_AGEMA_signal_9999 ;
    wire new_AGEMA_signal_10000 ;
    wire new_AGEMA_signal_10001 ;
    wire new_AGEMA_signal_10002 ;
    wire new_AGEMA_signal_10003 ;
    wire new_AGEMA_signal_10004 ;
    wire new_AGEMA_signal_10005 ;
    wire new_AGEMA_signal_10006 ;
    wire new_AGEMA_signal_10007 ;
    wire new_AGEMA_signal_10008 ;
    wire new_AGEMA_signal_10009 ;
    wire new_AGEMA_signal_10010 ;
    wire new_AGEMA_signal_10011 ;
    wire new_AGEMA_signal_10012 ;
    wire new_AGEMA_signal_10013 ;
    wire new_AGEMA_signal_10014 ;
    wire new_AGEMA_signal_10015 ;
    wire new_AGEMA_signal_10016 ;
    wire new_AGEMA_signal_10017 ;
    wire new_AGEMA_signal_10018 ;
    wire new_AGEMA_signal_10019 ;
    wire new_AGEMA_signal_10020 ;
    wire new_AGEMA_signal_10021 ;
    wire new_AGEMA_signal_10022 ;
    wire new_AGEMA_signal_10023 ;
    wire new_AGEMA_signal_10024 ;
    wire new_AGEMA_signal_10025 ;
    wire new_AGEMA_signal_10026 ;
    wire new_AGEMA_signal_10027 ;
    wire new_AGEMA_signal_10028 ;
    wire new_AGEMA_signal_10029 ;
    wire new_AGEMA_signal_10030 ;
    wire new_AGEMA_signal_10031 ;
    wire new_AGEMA_signal_10032 ;
    wire new_AGEMA_signal_10033 ;
    wire new_AGEMA_signal_10034 ;
    wire new_AGEMA_signal_10035 ;
    wire new_AGEMA_signal_10036 ;
    wire new_AGEMA_signal_10037 ;
    wire new_AGEMA_signal_10038 ;
    wire new_AGEMA_signal_10039 ;
    wire new_AGEMA_signal_10040 ;
    wire new_AGEMA_signal_10041 ;
    wire new_AGEMA_signal_10042 ;
    wire new_AGEMA_signal_10043 ;
    wire new_AGEMA_signal_10044 ;
    wire new_AGEMA_signal_10045 ;
    wire new_AGEMA_signal_10046 ;
    wire new_AGEMA_signal_10047 ;
    wire new_AGEMA_signal_10048 ;
    wire new_AGEMA_signal_10049 ;
    wire new_AGEMA_signal_10050 ;
    wire new_AGEMA_signal_10051 ;
    wire new_AGEMA_signal_10052 ;
    wire new_AGEMA_signal_10053 ;
    wire new_AGEMA_signal_10054 ;
    wire new_AGEMA_signal_10055 ;
    wire new_AGEMA_signal_10056 ;
    wire new_AGEMA_signal_10057 ;
    wire new_AGEMA_signal_10058 ;
    wire new_AGEMA_signal_10059 ;
    wire new_AGEMA_signal_10060 ;
    wire new_AGEMA_signal_10061 ;
    wire new_AGEMA_signal_10062 ;
    wire new_AGEMA_signal_10063 ;
    wire new_AGEMA_signal_10064 ;
    wire new_AGEMA_signal_10065 ;
    wire new_AGEMA_signal_10066 ;
    wire new_AGEMA_signal_10067 ;
    wire new_AGEMA_signal_10068 ;
    wire new_AGEMA_signal_10069 ;
    wire new_AGEMA_signal_10070 ;
    wire new_AGEMA_signal_10071 ;
    wire new_AGEMA_signal_10072 ;
    wire new_AGEMA_signal_10073 ;
    wire new_AGEMA_signal_10074 ;
    wire new_AGEMA_signal_10075 ;
    wire new_AGEMA_signal_10076 ;
    wire new_AGEMA_signal_10077 ;
    wire new_AGEMA_signal_10078 ;
    wire new_AGEMA_signal_10079 ;
    wire new_AGEMA_signal_10080 ;
    wire new_AGEMA_signal_10081 ;
    wire new_AGEMA_signal_10082 ;
    wire new_AGEMA_signal_10083 ;
    wire new_AGEMA_signal_10084 ;
    wire new_AGEMA_signal_10085 ;
    wire new_AGEMA_signal_10086 ;
    wire new_AGEMA_signal_10087 ;
    wire new_AGEMA_signal_10088 ;
    wire new_AGEMA_signal_10089 ;
    wire new_AGEMA_signal_10090 ;
    wire new_AGEMA_signal_10091 ;
    wire new_AGEMA_signal_10092 ;
    wire new_AGEMA_signal_10093 ;
    wire new_AGEMA_signal_10094 ;
    wire new_AGEMA_signal_10095 ;
    wire new_AGEMA_signal_10096 ;
    wire new_AGEMA_signal_10097 ;
    wire new_AGEMA_signal_10098 ;
    wire new_AGEMA_signal_10099 ;
    wire new_AGEMA_signal_10100 ;
    wire new_AGEMA_signal_10101 ;
    wire new_AGEMA_signal_10102 ;
    wire new_AGEMA_signal_10103 ;
    wire new_AGEMA_signal_10104 ;
    wire new_AGEMA_signal_10105 ;
    wire new_AGEMA_signal_10106 ;
    wire new_AGEMA_signal_10107 ;
    wire new_AGEMA_signal_10108 ;
    wire new_AGEMA_signal_10109 ;
    wire new_AGEMA_signal_10110 ;
    wire new_AGEMA_signal_10111 ;
    wire new_AGEMA_signal_10112 ;
    wire new_AGEMA_signal_10113 ;
    wire new_AGEMA_signal_10114 ;
    wire new_AGEMA_signal_10115 ;
    wire new_AGEMA_signal_10116 ;
    wire new_AGEMA_signal_10117 ;
    wire new_AGEMA_signal_10118 ;
    wire new_AGEMA_signal_10119 ;
    wire new_AGEMA_signal_10120 ;
    wire new_AGEMA_signal_10121 ;
    wire new_AGEMA_signal_10122 ;
    wire new_AGEMA_signal_10123 ;
    wire new_AGEMA_signal_10124 ;
    wire new_AGEMA_signal_10125 ;
    wire new_AGEMA_signal_10126 ;
    wire new_AGEMA_signal_10127 ;
    wire new_AGEMA_signal_10128 ;
    wire new_AGEMA_signal_10129 ;
    wire new_AGEMA_signal_10130 ;
    wire new_AGEMA_signal_10131 ;
    wire new_AGEMA_signal_10132 ;
    wire new_AGEMA_signal_10133 ;
    wire new_AGEMA_signal_10134 ;
    wire new_AGEMA_signal_10135 ;
    wire new_AGEMA_signal_10136 ;
    wire new_AGEMA_signal_10137 ;
    wire new_AGEMA_signal_10138 ;
    wire new_AGEMA_signal_10139 ;
    wire new_AGEMA_signal_10140 ;
    wire new_AGEMA_signal_10141 ;
    wire new_AGEMA_signal_10142 ;
    wire new_AGEMA_signal_10143 ;
    wire new_AGEMA_signal_10144 ;
    wire new_AGEMA_signal_10145 ;
    wire new_AGEMA_signal_10146 ;
    wire new_AGEMA_signal_10147 ;
    wire new_AGEMA_signal_10148 ;
    wire new_AGEMA_signal_10149 ;
    wire new_AGEMA_signal_10150 ;
    wire new_AGEMA_signal_10151 ;
    wire new_AGEMA_signal_10152 ;
    wire new_AGEMA_signal_10153 ;
    wire new_AGEMA_signal_10154 ;
    wire new_AGEMA_signal_10155 ;
    wire new_AGEMA_signal_10156 ;
    wire new_AGEMA_signal_10157 ;
    wire new_AGEMA_signal_10158 ;
    wire new_AGEMA_signal_10159 ;
    wire new_AGEMA_signal_10160 ;
    wire new_AGEMA_signal_10161 ;
    wire new_AGEMA_signal_10162 ;
    wire new_AGEMA_signal_10163 ;
    wire new_AGEMA_signal_10164 ;
    wire new_AGEMA_signal_10165 ;
    wire new_AGEMA_signal_10166 ;
    wire new_AGEMA_signal_10167 ;
    wire new_AGEMA_signal_10168 ;
    wire new_AGEMA_signal_10169 ;
    wire new_AGEMA_signal_10170 ;
    wire new_AGEMA_signal_10171 ;
    wire new_AGEMA_signal_10172 ;
    wire new_AGEMA_signal_10173 ;
    wire new_AGEMA_signal_10174 ;
    wire new_AGEMA_signal_10175 ;
    wire new_AGEMA_signal_10176 ;
    wire new_AGEMA_signal_10177 ;
    wire new_AGEMA_signal_10178 ;
    wire new_AGEMA_signal_10179 ;
    wire new_AGEMA_signal_10180 ;
    wire new_AGEMA_signal_10181 ;
    wire new_AGEMA_signal_10182 ;
    wire new_AGEMA_signal_10183 ;
    wire new_AGEMA_signal_10184 ;
    wire new_AGEMA_signal_10185 ;
    wire new_AGEMA_signal_10186 ;
    wire new_AGEMA_signal_10187 ;
    wire new_AGEMA_signal_10188 ;
    wire new_AGEMA_signal_10189 ;
    wire new_AGEMA_signal_10190 ;
    wire new_AGEMA_signal_10191 ;
    wire new_AGEMA_signal_10192 ;
    wire new_AGEMA_signal_10193 ;
    wire new_AGEMA_signal_10194 ;
    wire new_AGEMA_signal_10195 ;
    wire new_AGEMA_signal_10196 ;
    wire new_AGEMA_signal_10197 ;
    wire new_AGEMA_signal_10198 ;
    wire new_AGEMA_signal_10199 ;
    wire new_AGEMA_signal_10200 ;
    wire new_AGEMA_signal_10201 ;
    wire new_AGEMA_signal_10202 ;
    wire new_AGEMA_signal_10203 ;
    wire new_AGEMA_signal_10204 ;
    wire new_AGEMA_signal_10205 ;
    wire new_AGEMA_signal_10206 ;
    wire new_AGEMA_signal_10207 ;
    wire new_AGEMA_signal_10208 ;
    wire new_AGEMA_signal_10209 ;
    wire new_AGEMA_signal_10210 ;
    wire new_AGEMA_signal_10211 ;
    wire new_AGEMA_signal_10212 ;
    wire new_AGEMA_signal_10213 ;
    wire new_AGEMA_signal_10214 ;
    wire new_AGEMA_signal_10215 ;
    wire new_AGEMA_signal_10216 ;
    wire new_AGEMA_signal_10217 ;
    wire new_AGEMA_signal_10218 ;
    wire new_AGEMA_signal_10219 ;
    wire new_AGEMA_signal_10220 ;
    wire new_AGEMA_signal_10221 ;
    wire new_AGEMA_signal_10222 ;
    wire new_AGEMA_signal_10223 ;
    wire new_AGEMA_signal_10224 ;
    wire new_AGEMA_signal_10225 ;
    wire new_AGEMA_signal_10226 ;
    wire new_AGEMA_signal_10227 ;
    wire new_AGEMA_signal_10228 ;
    wire new_AGEMA_signal_10229 ;
    wire new_AGEMA_signal_10230 ;
    wire new_AGEMA_signal_10231 ;
    wire new_AGEMA_signal_10232 ;
    wire new_AGEMA_signal_10233 ;
    wire new_AGEMA_signal_10234 ;
    wire new_AGEMA_signal_10235 ;
    wire new_AGEMA_signal_10236 ;
    wire new_AGEMA_signal_10237 ;
    wire new_AGEMA_signal_10238 ;
    wire new_AGEMA_signal_10239 ;
    wire new_AGEMA_signal_10240 ;
    wire new_AGEMA_signal_10241 ;
    wire new_AGEMA_signal_10242 ;
    wire new_AGEMA_signal_10243 ;
    wire new_AGEMA_signal_10244 ;
    wire new_AGEMA_signal_10245 ;
    wire new_AGEMA_signal_10246 ;
    wire new_AGEMA_signal_10247 ;
    wire new_AGEMA_signal_10248 ;
    wire new_AGEMA_signal_10249 ;
    wire new_AGEMA_signal_10250 ;
    wire new_AGEMA_signal_10251 ;
    wire new_AGEMA_signal_10252 ;
    wire new_AGEMA_signal_10253 ;
    wire new_AGEMA_signal_10254 ;
    wire new_AGEMA_signal_10255 ;
    wire new_AGEMA_signal_10256 ;
    wire new_AGEMA_signal_10257 ;
    wire new_AGEMA_signal_10258 ;
    wire new_AGEMA_signal_10259 ;
    wire new_AGEMA_signal_10260 ;
    wire new_AGEMA_signal_10261 ;
    wire new_AGEMA_signal_10262 ;
    wire new_AGEMA_signal_10263 ;
    wire new_AGEMA_signal_10264 ;
    wire new_AGEMA_signal_10265 ;
    wire new_AGEMA_signal_10266 ;
    wire new_AGEMA_signal_10267 ;
    wire new_AGEMA_signal_10268 ;
    wire new_AGEMA_signal_10269 ;
    wire new_AGEMA_signal_10270 ;
    wire new_AGEMA_signal_10271 ;
    wire new_AGEMA_signal_10272 ;
    wire new_AGEMA_signal_10273 ;
    wire new_AGEMA_signal_10274 ;
    wire new_AGEMA_signal_10275 ;
    wire new_AGEMA_signal_10276 ;
    wire new_AGEMA_signal_10277 ;
    wire new_AGEMA_signal_10278 ;
    wire new_AGEMA_signal_10279 ;
    wire new_AGEMA_signal_10280 ;
    wire new_AGEMA_signal_10281 ;
    wire new_AGEMA_signal_10282 ;
    wire new_AGEMA_signal_10283 ;
    wire new_AGEMA_signal_10284 ;
    wire new_AGEMA_signal_10285 ;
    wire new_AGEMA_signal_10286 ;
    wire new_AGEMA_signal_10287 ;
    wire new_AGEMA_signal_10288 ;
    wire new_AGEMA_signal_10289 ;
    wire new_AGEMA_signal_10290 ;
    wire new_AGEMA_signal_10291 ;
    wire new_AGEMA_signal_10292 ;
    wire new_AGEMA_signal_10293 ;
    wire new_AGEMA_signal_10294 ;
    wire new_AGEMA_signal_10295 ;
    wire new_AGEMA_signal_10296 ;
    wire new_AGEMA_signal_10297 ;
    wire new_AGEMA_signal_10298 ;
    wire new_AGEMA_signal_10299 ;
    wire new_AGEMA_signal_10300 ;
    wire new_AGEMA_signal_10301 ;
    wire new_AGEMA_signal_10302 ;
    wire new_AGEMA_signal_10303 ;
    wire new_AGEMA_signal_10304 ;
    wire new_AGEMA_signal_10305 ;
    wire new_AGEMA_signal_10306 ;
    wire new_AGEMA_signal_10307 ;
    wire new_AGEMA_signal_10308 ;
    wire new_AGEMA_signal_10309 ;
    wire new_AGEMA_signal_10310 ;
    wire new_AGEMA_signal_10311 ;
    wire new_AGEMA_signal_10312 ;
    wire new_AGEMA_signal_10313 ;
    wire new_AGEMA_signal_10314 ;
    wire new_AGEMA_signal_10315 ;
    wire new_AGEMA_signal_10316 ;
    wire new_AGEMA_signal_10317 ;
    wire new_AGEMA_signal_10318 ;
    wire new_AGEMA_signal_10319 ;
    wire new_AGEMA_signal_10320 ;
    wire new_AGEMA_signal_10321 ;
    wire new_AGEMA_signal_10322 ;
    wire new_AGEMA_signal_10323 ;
    wire new_AGEMA_signal_10324 ;
    wire new_AGEMA_signal_10325 ;
    wire new_AGEMA_signal_10326 ;
    wire new_AGEMA_signal_10327 ;
    wire new_AGEMA_signal_10328 ;
    wire new_AGEMA_signal_10329 ;
    wire new_AGEMA_signal_10330 ;
    wire new_AGEMA_signal_10331 ;
    wire new_AGEMA_signal_10332 ;
    wire new_AGEMA_signal_10333 ;
    wire new_AGEMA_signal_10334 ;
    wire new_AGEMA_signal_10335 ;
    wire new_AGEMA_signal_10336 ;
    wire new_AGEMA_signal_10337 ;
    wire new_AGEMA_signal_10338 ;
    wire new_AGEMA_signal_10339 ;
    wire new_AGEMA_signal_10340 ;
    wire new_AGEMA_signal_10341 ;
    wire new_AGEMA_signal_10342 ;
    wire new_AGEMA_signal_10343 ;
    wire new_AGEMA_signal_10344 ;
    wire new_AGEMA_signal_10345 ;
    wire new_AGEMA_signal_10346 ;
    wire new_AGEMA_signal_10347 ;
    wire new_AGEMA_signal_10348 ;
    wire new_AGEMA_signal_10349 ;
    wire new_AGEMA_signal_10350 ;
    wire new_AGEMA_signal_10351 ;
    wire new_AGEMA_signal_10352 ;
    wire new_AGEMA_signal_10353 ;
    wire new_AGEMA_signal_10354 ;
    wire new_AGEMA_signal_10355 ;
    wire new_AGEMA_signal_10356 ;
    wire new_AGEMA_signal_10357 ;
    wire new_AGEMA_signal_10358 ;
    wire new_AGEMA_signal_10359 ;
    wire new_AGEMA_signal_10360 ;
    wire new_AGEMA_signal_10361 ;
    wire new_AGEMA_signal_10362 ;
    wire new_AGEMA_signal_10363 ;
    wire new_AGEMA_signal_10364 ;
    wire new_AGEMA_signal_10365 ;
    wire new_AGEMA_signal_10366 ;
    wire new_AGEMA_signal_10367 ;
    wire new_AGEMA_signal_10368 ;
    wire new_AGEMA_signal_10369 ;
    wire new_AGEMA_signal_10370 ;
    wire new_AGEMA_signal_10371 ;
    wire new_AGEMA_signal_10372 ;
    wire new_AGEMA_signal_10373 ;
    wire new_AGEMA_signal_10374 ;
    wire new_AGEMA_signal_10375 ;
    wire new_AGEMA_signal_10376 ;
    wire new_AGEMA_signal_10377 ;
    wire new_AGEMA_signal_10378 ;
    wire new_AGEMA_signal_10379 ;
    wire new_AGEMA_signal_10380 ;
    wire new_AGEMA_signal_10381 ;
    wire new_AGEMA_signal_10382 ;
    wire new_AGEMA_signal_10383 ;
    wire new_AGEMA_signal_10384 ;
    wire new_AGEMA_signal_10385 ;
    wire new_AGEMA_signal_10386 ;
    wire new_AGEMA_signal_10387 ;
    wire new_AGEMA_signal_10388 ;
    wire new_AGEMA_signal_10389 ;
    wire new_AGEMA_signal_10390 ;
    wire new_AGEMA_signal_10391 ;
    wire new_AGEMA_signal_10392 ;
    wire new_AGEMA_signal_10393 ;
    wire new_AGEMA_signal_10394 ;
    wire new_AGEMA_signal_10395 ;
    wire new_AGEMA_signal_10396 ;
    wire new_AGEMA_signal_10397 ;
    wire new_AGEMA_signal_10398 ;
    wire new_AGEMA_signal_10399 ;
    wire new_AGEMA_signal_10400 ;
    wire new_AGEMA_signal_10401 ;
    wire new_AGEMA_signal_10402 ;
    wire new_AGEMA_signal_10403 ;
    wire new_AGEMA_signal_10404 ;
    wire new_AGEMA_signal_10405 ;
    wire new_AGEMA_signal_10406 ;
    wire new_AGEMA_signal_10407 ;
    wire new_AGEMA_signal_10408 ;
    wire new_AGEMA_signal_10409 ;
    wire new_AGEMA_signal_10410 ;
    wire new_AGEMA_signal_10411 ;
    wire new_AGEMA_signal_10412 ;
    wire new_AGEMA_signal_10413 ;
    wire new_AGEMA_signal_10414 ;
    wire new_AGEMA_signal_10415 ;
    wire new_AGEMA_signal_10416 ;
    wire new_AGEMA_signal_10417 ;
    wire new_AGEMA_signal_10418 ;
    wire new_AGEMA_signal_10419 ;
    wire new_AGEMA_signal_10420 ;
    wire new_AGEMA_signal_10421 ;
    wire new_AGEMA_signal_10422 ;
    wire new_AGEMA_signal_10423 ;
    wire new_AGEMA_signal_10424 ;
    wire new_AGEMA_signal_10425 ;
    wire new_AGEMA_signal_10426 ;
    wire new_AGEMA_signal_10427 ;
    wire new_AGEMA_signal_10428 ;
    wire new_AGEMA_signal_10429 ;
    wire new_AGEMA_signal_10430 ;
    wire new_AGEMA_signal_10431 ;
    wire new_AGEMA_signal_10432 ;
    wire new_AGEMA_signal_10433 ;
    wire new_AGEMA_signal_10434 ;
    wire new_AGEMA_signal_10435 ;
    wire new_AGEMA_signal_10436 ;
    wire new_AGEMA_signal_10437 ;
    wire new_AGEMA_signal_10438 ;
    wire new_AGEMA_signal_10439 ;
    wire new_AGEMA_signal_10440 ;
    wire new_AGEMA_signal_10441 ;
    wire new_AGEMA_signal_10442 ;
    wire new_AGEMA_signal_10443 ;
    wire new_AGEMA_signal_10444 ;
    wire new_AGEMA_signal_10445 ;
    wire new_AGEMA_signal_10446 ;
    wire new_AGEMA_signal_10447 ;
    wire new_AGEMA_signal_10448 ;
    wire new_AGEMA_signal_10449 ;
    wire new_AGEMA_signal_10450 ;
    wire new_AGEMA_signal_10451 ;
    wire new_AGEMA_signal_10452 ;
    wire new_AGEMA_signal_10453 ;
    wire new_AGEMA_signal_10454 ;
    wire new_AGEMA_signal_10455 ;
    wire new_AGEMA_signal_10456 ;
    wire new_AGEMA_signal_10457 ;
    wire new_AGEMA_signal_10458 ;
    wire new_AGEMA_signal_10459 ;
    wire new_AGEMA_signal_10460 ;
    wire new_AGEMA_signal_10461 ;
    wire new_AGEMA_signal_10462 ;
    wire new_AGEMA_signal_10463 ;
    wire new_AGEMA_signal_10464 ;
    wire new_AGEMA_signal_10465 ;
    wire new_AGEMA_signal_10466 ;
    wire new_AGEMA_signal_10467 ;
    wire new_AGEMA_signal_10468 ;
    wire new_AGEMA_signal_10469 ;
    wire new_AGEMA_signal_10470 ;
    wire new_AGEMA_signal_10471 ;
    wire new_AGEMA_signal_10472 ;
    wire new_AGEMA_signal_10473 ;
    wire new_AGEMA_signal_10474 ;
    wire new_AGEMA_signal_10475 ;
    wire new_AGEMA_signal_10476 ;
    wire new_AGEMA_signal_10477 ;
    wire new_AGEMA_signal_10478 ;
    wire new_AGEMA_signal_10479 ;
    wire new_AGEMA_signal_10480 ;
    wire new_AGEMA_signal_10481 ;
    wire new_AGEMA_signal_10482 ;
    wire new_AGEMA_signal_10483 ;
    wire new_AGEMA_signal_10484 ;
    wire new_AGEMA_signal_10485 ;
    wire new_AGEMA_signal_10486 ;
    wire new_AGEMA_signal_10487 ;
    wire new_AGEMA_signal_10488 ;
    wire new_AGEMA_signal_10489 ;
    wire new_AGEMA_signal_10490 ;
    wire new_AGEMA_signal_10491 ;
    wire new_AGEMA_signal_10492 ;
    wire new_AGEMA_signal_10493 ;
    wire new_AGEMA_signal_10494 ;
    wire new_AGEMA_signal_10495 ;
    wire new_AGEMA_signal_10496 ;
    wire new_AGEMA_signal_10497 ;
    wire new_AGEMA_signal_10498 ;
    wire new_AGEMA_signal_10499 ;
    wire new_AGEMA_signal_10500 ;
    wire new_AGEMA_signal_10501 ;
    wire new_AGEMA_signal_10502 ;
    wire new_AGEMA_signal_10503 ;
    wire new_AGEMA_signal_10504 ;
    wire new_AGEMA_signal_10505 ;
    wire new_AGEMA_signal_10506 ;
    wire new_AGEMA_signal_10507 ;
    wire new_AGEMA_signal_10508 ;
    wire new_AGEMA_signal_10509 ;
    wire new_AGEMA_signal_10510 ;
    wire new_AGEMA_signal_10511 ;
    wire new_AGEMA_signal_10512 ;
    wire new_AGEMA_signal_10513 ;
    wire new_AGEMA_signal_10514 ;
    wire new_AGEMA_signal_10515 ;
    wire new_AGEMA_signal_10516 ;
    wire new_AGEMA_signal_10517 ;
    wire new_AGEMA_signal_10518 ;
    wire new_AGEMA_signal_10519 ;
    wire new_AGEMA_signal_10520 ;
    wire new_AGEMA_signal_10521 ;
    wire new_AGEMA_signal_10522 ;
    wire new_AGEMA_signal_10523 ;
    wire new_AGEMA_signal_10524 ;
    wire new_AGEMA_signal_10525 ;
    wire new_AGEMA_signal_10526 ;
    wire new_AGEMA_signal_10527 ;
    wire new_AGEMA_signal_10528 ;
    wire new_AGEMA_signal_10529 ;
    wire new_AGEMA_signal_10530 ;
    wire new_AGEMA_signal_10531 ;
    wire new_AGEMA_signal_10532 ;
    wire new_AGEMA_signal_10533 ;
    wire new_AGEMA_signal_10534 ;
    wire new_AGEMA_signal_10535 ;
    wire new_AGEMA_signal_10536 ;
    wire new_AGEMA_signal_10537 ;
    wire new_AGEMA_signal_10538 ;
    wire new_AGEMA_signal_10539 ;
    wire new_AGEMA_signal_10540 ;
    wire new_AGEMA_signal_10541 ;
    wire new_AGEMA_signal_10542 ;
    wire new_AGEMA_signal_10543 ;
    wire new_AGEMA_signal_10544 ;
    wire new_AGEMA_signal_10545 ;
    wire new_AGEMA_signal_10546 ;
    wire new_AGEMA_signal_10547 ;
    wire new_AGEMA_signal_10548 ;
    wire new_AGEMA_signal_10549 ;
    wire new_AGEMA_signal_10550 ;
    wire new_AGEMA_signal_10551 ;
    wire new_AGEMA_signal_10552 ;
    wire new_AGEMA_signal_10553 ;
    wire new_AGEMA_signal_10554 ;
    wire new_AGEMA_signal_10555 ;
    wire new_AGEMA_signal_10556 ;
    wire new_AGEMA_signal_10557 ;
    wire new_AGEMA_signal_10558 ;
    wire new_AGEMA_signal_10559 ;
    wire new_AGEMA_signal_10560 ;
    wire new_AGEMA_signal_10561 ;
    wire new_AGEMA_signal_10562 ;
    wire new_AGEMA_signal_10563 ;
    wire new_AGEMA_signal_10564 ;
    wire new_AGEMA_signal_10565 ;
    wire new_AGEMA_signal_10566 ;
    wire new_AGEMA_signal_10567 ;
    wire new_AGEMA_signal_10568 ;
    wire new_AGEMA_signal_10569 ;
    wire new_AGEMA_signal_10570 ;
    wire new_AGEMA_signal_10571 ;
    wire new_AGEMA_signal_10572 ;
    wire new_AGEMA_signal_10573 ;
    wire new_AGEMA_signal_10574 ;
    wire new_AGEMA_signal_10575 ;
    wire new_AGEMA_signal_10576 ;
    wire new_AGEMA_signal_10577 ;
    wire new_AGEMA_signal_10578 ;
    wire new_AGEMA_signal_10579 ;
    wire new_AGEMA_signal_10580 ;
    wire new_AGEMA_signal_10581 ;
    wire new_AGEMA_signal_10582 ;
    wire new_AGEMA_signal_10583 ;
    wire new_AGEMA_signal_10584 ;
    wire new_AGEMA_signal_10585 ;
    wire new_AGEMA_signal_10586 ;
    wire new_AGEMA_signal_10587 ;
    wire new_AGEMA_signal_10588 ;
    wire new_AGEMA_signal_10589 ;
    wire new_AGEMA_signal_10590 ;
    wire new_AGEMA_signal_10591 ;
    wire new_AGEMA_signal_10592 ;
    wire new_AGEMA_signal_10593 ;
    wire new_AGEMA_signal_10594 ;
    wire new_AGEMA_signal_10595 ;
    wire new_AGEMA_signal_10596 ;
    wire new_AGEMA_signal_10597 ;
    wire new_AGEMA_signal_10598 ;
    wire new_AGEMA_signal_10599 ;
    wire new_AGEMA_signal_10600 ;
    wire new_AGEMA_signal_10601 ;
    wire new_AGEMA_signal_10602 ;
    wire new_AGEMA_signal_10603 ;
    wire new_AGEMA_signal_10604 ;
    wire new_AGEMA_signal_10605 ;
    wire new_AGEMA_signal_10606 ;
    wire new_AGEMA_signal_10607 ;
    wire new_AGEMA_signal_10608 ;
    wire new_AGEMA_signal_10609 ;
    wire new_AGEMA_signal_10610 ;
    wire new_AGEMA_signal_10611 ;
    wire new_AGEMA_signal_10612 ;
    wire new_AGEMA_signal_10613 ;
    wire new_AGEMA_signal_10614 ;
    wire new_AGEMA_signal_10615 ;
    wire new_AGEMA_signal_10616 ;
    wire new_AGEMA_signal_10617 ;
    wire new_AGEMA_signal_10618 ;
    wire new_AGEMA_signal_10619 ;
    wire new_AGEMA_signal_10620 ;
    wire new_AGEMA_signal_10621 ;
    wire new_AGEMA_signal_10622 ;
    wire new_AGEMA_signal_10623 ;
    wire new_AGEMA_signal_10624 ;
    wire new_AGEMA_signal_10625 ;
    wire new_AGEMA_signal_10626 ;
    wire new_AGEMA_signal_10627 ;
    wire new_AGEMA_signal_10628 ;
    wire new_AGEMA_signal_10629 ;
    wire new_AGEMA_signal_10630 ;
    wire new_AGEMA_signal_10631 ;
    wire new_AGEMA_signal_10632 ;
    wire new_AGEMA_signal_10633 ;
    wire new_AGEMA_signal_10634 ;
    wire new_AGEMA_signal_10635 ;
    wire new_AGEMA_signal_10636 ;
    wire new_AGEMA_signal_10637 ;
    wire new_AGEMA_signal_10638 ;
    wire new_AGEMA_signal_10639 ;
    wire new_AGEMA_signal_10640 ;
    wire new_AGEMA_signal_10641 ;
    wire new_AGEMA_signal_10642 ;
    wire new_AGEMA_signal_10643 ;
    wire new_AGEMA_signal_10644 ;
    wire new_AGEMA_signal_10645 ;
    wire new_AGEMA_signal_10646 ;
    wire new_AGEMA_signal_10647 ;
    wire new_AGEMA_signal_10648 ;
    wire new_AGEMA_signal_10649 ;
    wire new_AGEMA_signal_10650 ;
    wire new_AGEMA_signal_10651 ;
    wire new_AGEMA_signal_10652 ;
    wire new_AGEMA_signal_10653 ;
    wire new_AGEMA_signal_10654 ;
    wire new_AGEMA_signal_10655 ;
    wire new_AGEMA_signal_10656 ;
    wire new_AGEMA_signal_10657 ;
    wire new_AGEMA_signal_10658 ;
    wire new_AGEMA_signal_10659 ;
    wire new_AGEMA_signal_10660 ;
    wire new_AGEMA_signal_10661 ;
    wire new_AGEMA_signal_10662 ;
    wire new_AGEMA_signal_10663 ;
    wire new_AGEMA_signal_10664 ;
    wire new_AGEMA_signal_10665 ;
    wire new_AGEMA_signal_10666 ;
    wire new_AGEMA_signal_10667 ;
    wire new_AGEMA_signal_10668 ;
    wire new_AGEMA_signal_10669 ;
    wire new_AGEMA_signal_10670 ;
    wire new_AGEMA_signal_10671 ;
    wire new_AGEMA_signal_10672 ;
    wire new_AGEMA_signal_10673 ;
    wire new_AGEMA_signal_10674 ;
    wire new_AGEMA_signal_10675 ;
    wire new_AGEMA_signal_10676 ;
    wire new_AGEMA_signal_10677 ;
    wire new_AGEMA_signal_10678 ;
    wire new_AGEMA_signal_10679 ;
    wire new_AGEMA_signal_10680 ;
    wire new_AGEMA_signal_10681 ;
    wire new_AGEMA_signal_10682 ;
    wire new_AGEMA_signal_10683 ;
    wire new_AGEMA_signal_10684 ;
    wire new_AGEMA_signal_10685 ;
    wire new_AGEMA_signal_10686 ;
    wire new_AGEMA_signal_10687 ;
    wire new_AGEMA_signal_10688 ;
    wire new_AGEMA_signal_10689 ;
    wire new_AGEMA_signal_10690 ;
    wire new_AGEMA_signal_10691 ;
    wire new_AGEMA_signal_10692 ;
    wire new_AGEMA_signal_10693 ;
    wire new_AGEMA_signal_10694 ;
    wire new_AGEMA_signal_10695 ;
    wire new_AGEMA_signal_10696 ;
    wire new_AGEMA_signal_10697 ;
    wire new_AGEMA_signal_10698 ;
    wire new_AGEMA_signal_10699 ;
    wire new_AGEMA_signal_10700 ;
    wire new_AGEMA_signal_10701 ;
    wire new_AGEMA_signal_10702 ;
    wire new_AGEMA_signal_10703 ;
    wire new_AGEMA_signal_10704 ;
    wire new_AGEMA_signal_10705 ;
    wire new_AGEMA_signal_10706 ;
    wire new_AGEMA_signal_10707 ;
    wire new_AGEMA_signal_10708 ;
    wire new_AGEMA_signal_10709 ;
    wire new_AGEMA_signal_10710 ;
    wire new_AGEMA_signal_10711 ;
    wire new_AGEMA_signal_10712 ;
    wire new_AGEMA_signal_10713 ;
    wire new_AGEMA_signal_10714 ;
    wire new_AGEMA_signal_10715 ;
    wire new_AGEMA_signal_10716 ;
    wire new_AGEMA_signal_10717 ;
    wire new_AGEMA_signal_10718 ;
    wire new_AGEMA_signal_10719 ;
    wire new_AGEMA_signal_10720 ;
    wire new_AGEMA_signal_10721 ;
    wire new_AGEMA_signal_10722 ;
    wire new_AGEMA_signal_10723 ;
    wire new_AGEMA_signal_10724 ;
    wire new_AGEMA_signal_10725 ;
    wire new_AGEMA_signal_10726 ;
    wire new_AGEMA_signal_10727 ;
    wire new_AGEMA_signal_10728 ;
    wire new_AGEMA_signal_10729 ;
    wire new_AGEMA_signal_10730 ;
    wire new_AGEMA_signal_10731 ;
    wire new_AGEMA_signal_10732 ;
    wire new_AGEMA_signal_10733 ;
    wire new_AGEMA_signal_10734 ;
    wire new_AGEMA_signal_10735 ;
    wire new_AGEMA_signal_10736 ;
    wire new_AGEMA_signal_10737 ;
    wire new_AGEMA_signal_10738 ;
    wire new_AGEMA_signal_10739 ;
    wire new_AGEMA_signal_10740 ;
    wire new_AGEMA_signal_10741 ;
    wire new_AGEMA_signal_10742 ;
    wire new_AGEMA_signal_10743 ;
    wire new_AGEMA_signal_10744 ;
    wire new_AGEMA_signal_10745 ;
    wire new_AGEMA_signal_10746 ;
    wire new_AGEMA_signal_10747 ;
    wire new_AGEMA_signal_10748 ;
    wire new_AGEMA_signal_10749 ;
    wire new_AGEMA_signal_10750 ;
    wire new_AGEMA_signal_10751 ;
    wire new_AGEMA_signal_10752 ;
    wire new_AGEMA_signal_10753 ;
    wire new_AGEMA_signal_10754 ;
    wire new_AGEMA_signal_10755 ;
    wire new_AGEMA_signal_10756 ;
    wire new_AGEMA_signal_10757 ;
    wire new_AGEMA_signal_10758 ;
    wire new_AGEMA_signal_10759 ;
    wire new_AGEMA_signal_10760 ;
    wire new_AGEMA_signal_10761 ;
    wire new_AGEMA_signal_10762 ;
    wire new_AGEMA_signal_10763 ;
    wire new_AGEMA_signal_10764 ;
    wire new_AGEMA_signal_10765 ;
    wire new_AGEMA_signal_10766 ;
    wire new_AGEMA_signal_10767 ;
    wire new_AGEMA_signal_10768 ;
    wire new_AGEMA_signal_10769 ;
    wire new_AGEMA_signal_10770 ;
    wire new_AGEMA_signal_10771 ;
    wire new_AGEMA_signal_10772 ;
    wire new_AGEMA_signal_10773 ;
    wire new_AGEMA_signal_10774 ;
    wire new_AGEMA_signal_10775 ;
    wire new_AGEMA_signal_10776 ;
    wire new_AGEMA_signal_10777 ;
    wire new_AGEMA_signal_10778 ;
    wire new_AGEMA_signal_10779 ;
    wire new_AGEMA_signal_10780 ;
    wire new_AGEMA_signal_10781 ;
    wire new_AGEMA_signal_10782 ;
    wire new_AGEMA_signal_10783 ;
    wire new_AGEMA_signal_10784 ;
    wire new_AGEMA_signal_10785 ;
    wire new_AGEMA_signal_10786 ;
    wire new_AGEMA_signal_10787 ;
    wire new_AGEMA_signal_10788 ;
    wire new_AGEMA_signal_10789 ;
    wire new_AGEMA_signal_10790 ;
    wire new_AGEMA_signal_10791 ;
    wire new_AGEMA_signal_10792 ;
    wire new_AGEMA_signal_10793 ;
    wire new_AGEMA_signal_10794 ;
    wire new_AGEMA_signal_10795 ;
    wire new_AGEMA_signal_10796 ;
    wire new_AGEMA_signal_10797 ;
    wire new_AGEMA_signal_10798 ;
    wire new_AGEMA_signal_10799 ;
    wire new_AGEMA_signal_10800 ;
    wire new_AGEMA_signal_10801 ;
    wire new_AGEMA_signal_10802 ;
    wire new_AGEMA_signal_10803 ;
    wire new_AGEMA_signal_10804 ;
    wire new_AGEMA_signal_10805 ;
    wire new_AGEMA_signal_10806 ;
    wire new_AGEMA_signal_10807 ;
    wire new_AGEMA_signal_10808 ;
    wire new_AGEMA_signal_10809 ;
    wire new_AGEMA_signal_10810 ;
    wire new_AGEMA_signal_10811 ;
    wire new_AGEMA_signal_10812 ;
    wire new_AGEMA_signal_10813 ;
    wire new_AGEMA_signal_10814 ;
    wire new_AGEMA_signal_10815 ;
    wire new_AGEMA_signal_10816 ;
    wire new_AGEMA_signal_10817 ;
    wire new_AGEMA_signal_10818 ;
    wire new_AGEMA_signal_10819 ;
    wire new_AGEMA_signal_10820 ;
    wire new_AGEMA_signal_10821 ;
    wire new_AGEMA_signal_10822 ;
    wire new_AGEMA_signal_10823 ;
    wire new_AGEMA_signal_10824 ;
    wire new_AGEMA_signal_10825 ;
    wire new_AGEMA_signal_10826 ;
    wire new_AGEMA_signal_10827 ;
    wire new_AGEMA_signal_10828 ;
    wire new_AGEMA_signal_10829 ;
    wire new_AGEMA_signal_10830 ;
    wire new_AGEMA_signal_10831 ;
    wire new_AGEMA_signal_10832 ;
    wire new_AGEMA_signal_10833 ;
    wire new_AGEMA_signal_10834 ;
    wire new_AGEMA_signal_10835 ;
    wire new_AGEMA_signal_10836 ;
    wire new_AGEMA_signal_10837 ;
    wire new_AGEMA_signal_10838 ;
    wire new_AGEMA_signal_10839 ;
    wire new_AGEMA_signal_10840 ;
    wire new_AGEMA_signal_10841 ;
    wire new_AGEMA_signal_10842 ;
    wire new_AGEMA_signal_10843 ;
    wire new_AGEMA_signal_10844 ;
    wire new_AGEMA_signal_10845 ;
    wire new_AGEMA_signal_10846 ;
    wire new_AGEMA_signal_10847 ;
    wire new_AGEMA_signal_10848 ;
    wire new_AGEMA_signal_10849 ;
    wire new_AGEMA_signal_10850 ;
    wire new_AGEMA_signal_10851 ;
    wire new_AGEMA_signal_10852 ;
    wire new_AGEMA_signal_10853 ;
    wire new_AGEMA_signal_10854 ;
    wire new_AGEMA_signal_10855 ;
    wire new_AGEMA_signal_10856 ;
    wire new_AGEMA_signal_10857 ;
    wire new_AGEMA_signal_10858 ;
    wire new_AGEMA_signal_10859 ;
    wire new_AGEMA_signal_10860 ;
    wire new_AGEMA_signal_10861 ;
    wire new_AGEMA_signal_10862 ;
    wire new_AGEMA_signal_10863 ;
    wire new_AGEMA_signal_10864 ;
    wire new_AGEMA_signal_10865 ;
    wire new_AGEMA_signal_10866 ;
    wire new_AGEMA_signal_10867 ;
    wire new_AGEMA_signal_10868 ;
    wire new_AGEMA_signal_10869 ;
    wire new_AGEMA_signal_10870 ;
    wire new_AGEMA_signal_10871 ;
    wire new_AGEMA_signal_10872 ;
    wire new_AGEMA_signal_10873 ;
    wire new_AGEMA_signal_10874 ;
    wire new_AGEMA_signal_10875 ;
    wire new_AGEMA_signal_10876 ;
    wire new_AGEMA_signal_10877 ;
    wire new_AGEMA_signal_10878 ;
    wire new_AGEMA_signal_10879 ;
    wire new_AGEMA_signal_10880 ;
    wire new_AGEMA_signal_10881 ;
    wire new_AGEMA_signal_10882 ;
    wire new_AGEMA_signal_10883 ;
    wire new_AGEMA_signal_10884 ;
    wire new_AGEMA_signal_10885 ;
    wire new_AGEMA_signal_10886 ;
    wire new_AGEMA_signal_10887 ;
    wire new_AGEMA_signal_10888 ;
    wire new_AGEMA_signal_10889 ;
    wire new_AGEMA_signal_10890 ;
    wire new_AGEMA_signal_10891 ;
    wire new_AGEMA_signal_10892 ;
    wire new_AGEMA_signal_10893 ;
    wire new_AGEMA_signal_10894 ;
    wire new_AGEMA_signal_10895 ;
    wire new_AGEMA_signal_10896 ;
    wire new_AGEMA_signal_10897 ;
    wire new_AGEMA_signal_10898 ;
    wire new_AGEMA_signal_10899 ;
    wire new_AGEMA_signal_10900 ;
    wire new_AGEMA_signal_10901 ;
    wire new_AGEMA_signal_10902 ;
    wire new_AGEMA_signal_10903 ;
    wire new_AGEMA_signal_10904 ;
    wire new_AGEMA_signal_10905 ;
    wire new_AGEMA_signal_10906 ;
    wire new_AGEMA_signal_10907 ;
    wire new_AGEMA_signal_10908 ;
    wire new_AGEMA_signal_10909 ;
    wire new_AGEMA_signal_10910 ;
    wire new_AGEMA_signal_10911 ;
    wire new_AGEMA_signal_10912 ;
    wire new_AGEMA_signal_10913 ;
    wire new_AGEMA_signal_10914 ;
    wire new_AGEMA_signal_10915 ;
    wire new_AGEMA_signal_10916 ;
    wire new_AGEMA_signal_10917 ;
    wire new_AGEMA_signal_10918 ;
    wire new_AGEMA_signal_10919 ;
    wire new_AGEMA_signal_10920 ;
    wire new_AGEMA_signal_10921 ;
    wire new_AGEMA_signal_10922 ;
    wire new_AGEMA_signal_10923 ;
    wire new_AGEMA_signal_10924 ;
    wire new_AGEMA_signal_10925 ;
    wire new_AGEMA_signal_10926 ;
    wire new_AGEMA_signal_10927 ;
    wire new_AGEMA_signal_10928 ;
    wire new_AGEMA_signal_10929 ;
    wire new_AGEMA_signal_10930 ;
    wire new_AGEMA_signal_10931 ;
    wire new_AGEMA_signal_10932 ;
    wire new_AGEMA_signal_10933 ;
    wire new_AGEMA_signal_10934 ;
    wire new_AGEMA_signal_10935 ;
    wire new_AGEMA_signal_10936 ;
    wire new_AGEMA_signal_10937 ;
    wire new_AGEMA_signal_10938 ;
    wire new_AGEMA_signal_10939 ;
    wire new_AGEMA_signal_10940 ;
    wire new_AGEMA_signal_10941 ;
    wire new_AGEMA_signal_10942 ;
    wire new_AGEMA_signal_10943 ;
    wire new_AGEMA_signal_10944 ;
    wire new_AGEMA_signal_10945 ;
    wire new_AGEMA_signal_10946 ;
    wire new_AGEMA_signal_10947 ;
    wire new_AGEMA_signal_10948 ;
    wire new_AGEMA_signal_10949 ;
    wire new_AGEMA_signal_10950 ;
    wire new_AGEMA_signal_10951 ;
    wire new_AGEMA_signal_10952 ;
    wire new_AGEMA_signal_10953 ;
    wire new_AGEMA_signal_10954 ;
    wire new_AGEMA_signal_10955 ;
    wire new_AGEMA_signal_10956 ;
    wire new_AGEMA_signal_10957 ;
    wire new_AGEMA_signal_10958 ;
    wire new_AGEMA_signal_10959 ;
    wire new_AGEMA_signal_10960 ;
    wire new_AGEMA_signal_10961 ;
    wire new_AGEMA_signal_10962 ;
    wire new_AGEMA_signal_10963 ;
    wire new_AGEMA_signal_10964 ;
    wire new_AGEMA_signal_10965 ;
    wire new_AGEMA_signal_10966 ;
    wire new_AGEMA_signal_10967 ;
    wire new_AGEMA_signal_10968 ;
    wire new_AGEMA_signal_10969 ;
    wire new_AGEMA_signal_10970 ;
    wire new_AGEMA_signal_10971 ;
    wire new_AGEMA_signal_10972 ;
    wire new_AGEMA_signal_10973 ;
    wire new_AGEMA_signal_10974 ;
    wire new_AGEMA_signal_10975 ;
    wire new_AGEMA_signal_10976 ;
    wire new_AGEMA_signal_10977 ;
    wire new_AGEMA_signal_10978 ;
    wire new_AGEMA_signal_10979 ;
    wire new_AGEMA_signal_10980 ;
    wire new_AGEMA_signal_10981 ;
    wire new_AGEMA_signal_10982 ;
    wire new_AGEMA_signal_10983 ;
    wire new_AGEMA_signal_10984 ;
    wire new_AGEMA_signal_10985 ;
    wire new_AGEMA_signal_10986 ;
    wire new_AGEMA_signal_10987 ;
    wire new_AGEMA_signal_10988 ;
    wire new_AGEMA_signal_10989 ;
    wire new_AGEMA_signal_10990 ;
    wire new_AGEMA_signal_10991 ;
    wire new_AGEMA_signal_10992 ;
    wire new_AGEMA_signal_10993 ;
    wire new_AGEMA_signal_10994 ;
    wire new_AGEMA_signal_10995 ;
    wire new_AGEMA_signal_10996 ;
    wire new_AGEMA_signal_10997 ;
    wire new_AGEMA_signal_10998 ;
    wire new_AGEMA_signal_10999 ;
    wire new_AGEMA_signal_11000 ;
    wire new_AGEMA_signal_11001 ;
    wire new_AGEMA_signal_11002 ;
    wire new_AGEMA_signal_11003 ;
    wire new_AGEMA_signal_11004 ;
    wire new_AGEMA_signal_11005 ;
    wire new_AGEMA_signal_11006 ;
    wire new_AGEMA_signal_11007 ;
    wire new_AGEMA_signal_11008 ;
    wire new_AGEMA_signal_11009 ;
    wire new_AGEMA_signal_11010 ;
    wire new_AGEMA_signal_11011 ;
    wire new_AGEMA_signal_11012 ;
    wire new_AGEMA_signal_11013 ;
    wire new_AGEMA_signal_11014 ;
    wire new_AGEMA_signal_11015 ;
    wire new_AGEMA_signal_11016 ;
    wire new_AGEMA_signal_11017 ;
    wire new_AGEMA_signal_11018 ;
    wire new_AGEMA_signal_11019 ;
    wire new_AGEMA_signal_11020 ;
    wire new_AGEMA_signal_11021 ;
    wire new_AGEMA_signal_11022 ;
    wire new_AGEMA_signal_11023 ;
    wire new_AGEMA_signal_11024 ;
    wire new_AGEMA_signal_11025 ;
    wire new_AGEMA_signal_11026 ;
    wire new_AGEMA_signal_11027 ;
    wire new_AGEMA_signal_11028 ;
    wire new_AGEMA_signal_11029 ;
    wire new_AGEMA_signal_11030 ;
    wire new_AGEMA_signal_11031 ;
    wire new_AGEMA_signal_11032 ;
    wire new_AGEMA_signal_11033 ;
    wire new_AGEMA_signal_11034 ;
    wire new_AGEMA_signal_11035 ;
    wire new_AGEMA_signal_11036 ;
    wire new_AGEMA_signal_11037 ;
    wire new_AGEMA_signal_11038 ;
    wire new_AGEMA_signal_11039 ;
    wire new_AGEMA_signal_11040 ;
    wire new_AGEMA_signal_11041 ;
    wire new_AGEMA_signal_11042 ;
    wire new_AGEMA_signal_11043 ;
    wire new_AGEMA_signal_11044 ;
    wire new_AGEMA_signal_11045 ;
    wire new_AGEMA_signal_11046 ;
    wire new_AGEMA_signal_11047 ;
    wire new_AGEMA_signal_11048 ;
    wire new_AGEMA_signal_11049 ;
    wire new_AGEMA_signal_11050 ;
    wire new_AGEMA_signal_11051 ;
    wire new_AGEMA_signal_11052 ;
    wire new_AGEMA_signal_11053 ;
    wire new_AGEMA_signal_11054 ;
    wire new_AGEMA_signal_11055 ;
    wire new_AGEMA_signal_11056 ;
    wire new_AGEMA_signal_11057 ;
    wire new_AGEMA_signal_11058 ;
    wire new_AGEMA_signal_11059 ;
    wire new_AGEMA_signal_11060 ;
    wire new_AGEMA_signal_11061 ;
    wire new_AGEMA_signal_11062 ;
    wire new_AGEMA_signal_11063 ;
    wire new_AGEMA_signal_11064 ;
    wire new_AGEMA_signal_11065 ;
    wire new_AGEMA_signal_11066 ;
    wire new_AGEMA_signal_11067 ;
    wire new_AGEMA_signal_11068 ;
    wire new_AGEMA_signal_11069 ;
    wire new_AGEMA_signal_11070 ;
    wire new_AGEMA_signal_11071 ;
    wire new_AGEMA_signal_11072 ;
    wire new_AGEMA_signal_11073 ;
    wire new_AGEMA_signal_11074 ;
    wire new_AGEMA_signal_11075 ;
    wire new_AGEMA_signal_11076 ;
    wire new_AGEMA_signal_11077 ;
    wire new_AGEMA_signal_11078 ;
    wire new_AGEMA_signal_11079 ;
    wire new_AGEMA_signal_11080 ;
    wire new_AGEMA_signal_11081 ;
    wire new_AGEMA_signal_11082 ;
    wire new_AGEMA_signal_11083 ;
    wire new_AGEMA_signal_11084 ;
    wire new_AGEMA_signal_11085 ;
    wire new_AGEMA_signal_11086 ;
    wire new_AGEMA_signal_11087 ;
    wire new_AGEMA_signal_11088 ;
    wire new_AGEMA_signal_11089 ;
    wire new_AGEMA_signal_11090 ;
    wire new_AGEMA_signal_11091 ;
    wire new_AGEMA_signal_11092 ;
    wire new_AGEMA_signal_11093 ;
    wire new_AGEMA_signal_11094 ;
    wire new_AGEMA_signal_11095 ;
    wire new_AGEMA_signal_11096 ;
    wire new_AGEMA_signal_11097 ;
    wire new_AGEMA_signal_11098 ;
    wire new_AGEMA_signal_11099 ;
    wire new_AGEMA_signal_11100 ;
    wire new_AGEMA_signal_11101 ;
    wire new_AGEMA_signal_11102 ;
    wire new_AGEMA_signal_11103 ;
    wire new_AGEMA_signal_11104 ;
    wire new_AGEMA_signal_11105 ;
    wire new_AGEMA_signal_11106 ;
    wire new_AGEMA_signal_11107 ;
    wire new_AGEMA_signal_11108 ;
    wire new_AGEMA_signal_11109 ;
    wire new_AGEMA_signal_11110 ;
    wire new_AGEMA_signal_11111 ;
    wire new_AGEMA_signal_11112 ;
    wire new_AGEMA_signal_11113 ;
    wire new_AGEMA_signal_11114 ;
    wire new_AGEMA_signal_11115 ;
    wire new_AGEMA_signal_11116 ;
    wire new_AGEMA_signal_11117 ;
    wire new_AGEMA_signal_11118 ;
    wire new_AGEMA_signal_11119 ;
    wire new_AGEMA_signal_11120 ;
    wire new_AGEMA_signal_11121 ;
    wire new_AGEMA_signal_11122 ;
    wire new_AGEMA_signal_11123 ;
    wire new_AGEMA_signal_11124 ;
    wire new_AGEMA_signal_11125 ;
    wire new_AGEMA_signal_11126 ;
    wire new_AGEMA_signal_11127 ;
    wire new_AGEMA_signal_11128 ;
    wire new_AGEMA_signal_11129 ;
    wire new_AGEMA_signal_11130 ;
    wire new_AGEMA_signal_11131 ;
    wire new_AGEMA_signal_11132 ;
    wire new_AGEMA_signal_11133 ;
    wire new_AGEMA_signal_11134 ;
    wire new_AGEMA_signal_11135 ;
    wire new_AGEMA_signal_11136 ;
    wire new_AGEMA_signal_11137 ;
    wire new_AGEMA_signal_11138 ;
    wire new_AGEMA_signal_11139 ;
    wire new_AGEMA_signal_11140 ;
    wire new_AGEMA_signal_11141 ;
    wire new_AGEMA_signal_11142 ;
    wire new_AGEMA_signal_11143 ;
    wire new_AGEMA_signal_11144 ;
    wire new_AGEMA_signal_11145 ;
    wire new_AGEMA_signal_11146 ;
    wire new_AGEMA_signal_11147 ;
    wire new_AGEMA_signal_11148 ;
    wire new_AGEMA_signal_11149 ;
    wire new_AGEMA_signal_11150 ;
    wire new_AGEMA_signal_11151 ;
    wire new_AGEMA_signal_11152 ;
    wire new_AGEMA_signal_11153 ;
    wire new_AGEMA_signal_11154 ;
    wire new_AGEMA_signal_11155 ;
    wire new_AGEMA_signal_11156 ;
    wire new_AGEMA_signal_11157 ;
    wire new_AGEMA_signal_11158 ;
    wire new_AGEMA_signal_11159 ;
    wire new_AGEMA_signal_11160 ;
    wire new_AGEMA_signal_11161 ;
    wire new_AGEMA_signal_11162 ;
    wire new_AGEMA_signal_11163 ;
    wire new_AGEMA_signal_11164 ;
    wire new_AGEMA_signal_11165 ;
    wire new_AGEMA_signal_11166 ;
    wire new_AGEMA_signal_11167 ;
    wire new_AGEMA_signal_11168 ;
    wire new_AGEMA_signal_11169 ;
    wire new_AGEMA_signal_11170 ;
    wire new_AGEMA_signal_11171 ;
    wire new_AGEMA_signal_11172 ;
    wire new_AGEMA_signal_11173 ;
    wire new_AGEMA_signal_11174 ;
    wire new_AGEMA_signal_11175 ;
    wire new_AGEMA_signal_11176 ;
    wire new_AGEMA_signal_11177 ;
    wire new_AGEMA_signal_11178 ;
    wire new_AGEMA_signal_11179 ;
    wire new_AGEMA_signal_11180 ;
    wire new_AGEMA_signal_11181 ;
    wire new_AGEMA_signal_11182 ;
    wire new_AGEMA_signal_11183 ;
    wire new_AGEMA_signal_11184 ;
    wire new_AGEMA_signal_11185 ;
    wire new_AGEMA_signal_11186 ;
    wire new_AGEMA_signal_11187 ;
    wire new_AGEMA_signal_11188 ;
    wire new_AGEMA_signal_11189 ;
    wire new_AGEMA_signal_11190 ;
    wire new_AGEMA_signal_11191 ;
    wire new_AGEMA_signal_11192 ;
    wire new_AGEMA_signal_11193 ;
    wire new_AGEMA_signal_11194 ;
    wire new_AGEMA_signal_11195 ;
    wire new_AGEMA_signal_11196 ;
    wire new_AGEMA_signal_11197 ;
    wire new_AGEMA_signal_11198 ;
    wire new_AGEMA_signal_11199 ;
    wire new_AGEMA_signal_11200 ;
    wire new_AGEMA_signal_11201 ;
    wire new_AGEMA_signal_11202 ;
    wire new_AGEMA_signal_11203 ;
    wire new_AGEMA_signal_11204 ;
    wire new_AGEMA_signal_11205 ;
    wire new_AGEMA_signal_11206 ;
    wire new_AGEMA_signal_11207 ;
    wire new_AGEMA_signal_11208 ;
    wire new_AGEMA_signal_11209 ;
    wire new_AGEMA_signal_11210 ;
    wire new_AGEMA_signal_11211 ;
    wire new_AGEMA_signal_11212 ;
    wire new_AGEMA_signal_11213 ;
    wire new_AGEMA_signal_11214 ;
    wire new_AGEMA_signal_11215 ;
    wire new_AGEMA_signal_11216 ;
    wire new_AGEMA_signal_11217 ;
    wire new_AGEMA_signal_11218 ;
    wire new_AGEMA_signal_11219 ;
    wire new_AGEMA_signal_11220 ;
    wire new_AGEMA_signal_11221 ;
    wire new_AGEMA_signal_11222 ;
    wire new_AGEMA_signal_11223 ;
    wire new_AGEMA_signal_11224 ;
    wire new_AGEMA_signal_11225 ;
    wire new_AGEMA_signal_11226 ;
    wire new_AGEMA_signal_11227 ;
    wire new_AGEMA_signal_11228 ;
    wire new_AGEMA_signal_11229 ;
    wire new_AGEMA_signal_11230 ;
    wire new_AGEMA_signal_11231 ;
    wire new_AGEMA_signal_11232 ;
    wire new_AGEMA_signal_11233 ;
    wire new_AGEMA_signal_11234 ;
    wire new_AGEMA_signal_11235 ;
    wire new_AGEMA_signal_11236 ;
    wire new_AGEMA_signal_11237 ;
    wire new_AGEMA_signal_11238 ;
    wire new_AGEMA_signal_11239 ;
    wire new_AGEMA_signal_11240 ;
    wire new_AGEMA_signal_11241 ;
    wire new_AGEMA_signal_11242 ;
    wire new_AGEMA_signal_11243 ;
    wire new_AGEMA_signal_11244 ;
    wire new_AGEMA_signal_11245 ;
    wire new_AGEMA_signal_11246 ;
    wire new_AGEMA_signal_11247 ;
    wire new_AGEMA_signal_11248 ;
    wire new_AGEMA_signal_11249 ;
    wire new_AGEMA_signal_11250 ;
    wire new_AGEMA_signal_11251 ;
    wire new_AGEMA_signal_11252 ;
    wire new_AGEMA_signal_11253 ;
    wire new_AGEMA_signal_11254 ;
    wire new_AGEMA_signal_11255 ;
    wire new_AGEMA_signal_11256 ;
    wire new_AGEMA_signal_11257 ;
    wire new_AGEMA_signal_11258 ;
    wire new_AGEMA_signal_11259 ;
    wire new_AGEMA_signal_11260 ;
    wire new_AGEMA_signal_11261 ;
    wire new_AGEMA_signal_11262 ;
    wire new_AGEMA_signal_11263 ;
    wire new_AGEMA_signal_11264 ;
    wire new_AGEMA_signal_11265 ;
    wire new_AGEMA_signal_11266 ;
    wire new_AGEMA_signal_11267 ;
    wire new_AGEMA_signal_11268 ;
    wire new_AGEMA_signal_11269 ;
    wire new_AGEMA_signal_11270 ;
    wire new_AGEMA_signal_11271 ;
    wire new_AGEMA_signal_11272 ;
    wire new_AGEMA_signal_11273 ;
    wire new_AGEMA_signal_11274 ;
    wire new_AGEMA_signal_11275 ;
    wire new_AGEMA_signal_11276 ;
    wire new_AGEMA_signal_11277 ;
    wire new_AGEMA_signal_11278 ;
    wire new_AGEMA_signal_11279 ;
    wire new_AGEMA_signal_11280 ;
    wire new_AGEMA_signal_11281 ;
    wire new_AGEMA_signal_11282 ;
    wire new_AGEMA_signal_11283 ;
    wire new_AGEMA_signal_11284 ;
    wire new_AGEMA_signal_11285 ;
    wire new_AGEMA_signal_11286 ;
    wire new_AGEMA_signal_11287 ;
    wire new_AGEMA_signal_11288 ;
    wire new_AGEMA_signal_11289 ;
    wire new_AGEMA_signal_11290 ;
    wire new_AGEMA_signal_11291 ;
    wire new_AGEMA_signal_11292 ;
    wire new_AGEMA_signal_11293 ;
    wire new_AGEMA_signal_11294 ;
    wire new_AGEMA_signal_11295 ;
    wire new_AGEMA_signal_11296 ;
    wire new_AGEMA_signal_11297 ;
    wire new_AGEMA_signal_11298 ;
    wire new_AGEMA_signal_11299 ;
    wire new_AGEMA_signal_11300 ;
    wire new_AGEMA_signal_11301 ;
    wire new_AGEMA_signal_11302 ;
    wire new_AGEMA_signal_11303 ;
    wire new_AGEMA_signal_11304 ;
    wire new_AGEMA_signal_11305 ;
    wire new_AGEMA_signal_11306 ;
    wire new_AGEMA_signal_11307 ;
    wire new_AGEMA_signal_11308 ;
    wire new_AGEMA_signal_11309 ;
    wire new_AGEMA_signal_11310 ;
    wire new_AGEMA_signal_11311 ;
    wire new_AGEMA_signal_11312 ;
    wire new_AGEMA_signal_11313 ;
    wire new_AGEMA_signal_11314 ;
    wire new_AGEMA_signal_11315 ;
    wire new_AGEMA_signal_11316 ;
    wire new_AGEMA_signal_11317 ;
    wire new_AGEMA_signal_11318 ;
    wire new_AGEMA_signal_11319 ;
    wire new_AGEMA_signal_11320 ;
    wire new_AGEMA_signal_11321 ;
    wire new_AGEMA_signal_11322 ;
    wire new_AGEMA_signal_11323 ;
    wire new_AGEMA_signal_11324 ;
    wire new_AGEMA_signal_11325 ;
    wire new_AGEMA_signal_11326 ;
    wire new_AGEMA_signal_11327 ;
    wire new_AGEMA_signal_11328 ;
    wire new_AGEMA_signal_11329 ;
    wire new_AGEMA_signal_11330 ;
    wire new_AGEMA_signal_11331 ;
    wire new_AGEMA_signal_11332 ;
    wire new_AGEMA_signal_11333 ;
    wire new_AGEMA_signal_11334 ;
    wire new_AGEMA_signal_11335 ;
    wire new_AGEMA_signal_11336 ;
    wire new_AGEMA_signal_11337 ;
    wire new_AGEMA_signal_11338 ;
    wire new_AGEMA_signal_11339 ;
    wire new_AGEMA_signal_11340 ;
    wire new_AGEMA_signal_11341 ;
    wire new_AGEMA_signal_11342 ;
    wire new_AGEMA_signal_11343 ;
    wire new_AGEMA_signal_11344 ;
    wire new_AGEMA_signal_11345 ;
    wire new_AGEMA_signal_11346 ;
    wire new_AGEMA_signal_11347 ;
    wire new_AGEMA_signal_11348 ;
    wire new_AGEMA_signal_11349 ;
    wire new_AGEMA_signal_11350 ;
    wire new_AGEMA_signal_11351 ;
    wire new_AGEMA_signal_11352 ;
    wire new_AGEMA_signal_11353 ;
    wire new_AGEMA_signal_11354 ;
    wire new_AGEMA_signal_11355 ;
    wire new_AGEMA_signal_11356 ;
    wire new_AGEMA_signal_11357 ;
    wire new_AGEMA_signal_11358 ;
    wire new_AGEMA_signal_11359 ;
    wire new_AGEMA_signal_11360 ;
    wire new_AGEMA_signal_11361 ;
    wire new_AGEMA_signal_11362 ;
    wire new_AGEMA_signal_11363 ;
    wire new_AGEMA_signal_11364 ;
    wire new_AGEMA_signal_11365 ;
    wire new_AGEMA_signal_11366 ;
    wire new_AGEMA_signal_11367 ;
    wire new_AGEMA_signal_11368 ;
    wire new_AGEMA_signal_11369 ;
    wire new_AGEMA_signal_11370 ;
    wire new_AGEMA_signal_11371 ;
    wire new_AGEMA_signal_11372 ;
    wire new_AGEMA_signal_11373 ;
    wire new_AGEMA_signal_11374 ;
    wire new_AGEMA_signal_11375 ;
    wire new_AGEMA_signal_11376 ;
    wire new_AGEMA_signal_11377 ;
    wire new_AGEMA_signal_11378 ;
    wire new_AGEMA_signal_11379 ;
    wire new_AGEMA_signal_11380 ;
    wire new_AGEMA_signal_11381 ;
    wire new_AGEMA_signal_11382 ;
    wire new_AGEMA_signal_11383 ;
    wire new_AGEMA_signal_11384 ;
    wire new_AGEMA_signal_11385 ;
    wire new_AGEMA_signal_11386 ;
    wire new_AGEMA_signal_11387 ;
    wire new_AGEMA_signal_11388 ;
    wire new_AGEMA_signal_11389 ;
    wire new_AGEMA_signal_11390 ;
    wire new_AGEMA_signal_11391 ;
    wire new_AGEMA_signal_11392 ;
    wire new_AGEMA_signal_11393 ;
    wire new_AGEMA_signal_11394 ;
    wire new_AGEMA_signal_11395 ;
    wire new_AGEMA_signal_11396 ;
    wire new_AGEMA_signal_11397 ;
    wire new_AGEMA_signal_11398 ;
    wire new_AGEMA_signal_11399 ;
    wire new_AGEMA_signal_11400 ;
    wire new_AGEMA_signal_11401 ;
    wire new_AGEMA_signal_11402 ;
    wire new_AGEMA_signal_11403 ;
    wire new_AGEMA_signal_11404 ;
    wire new_AGEMA_signal_11405 ;
    wire new_AGEMA_signal_11406 ;
    wire new_AGEMA_signal_11407 ;
    wire new_AGEMA_signal_11408 ;
    wire new_AGEMA_signal_11409 ;
    wire new_AGEMA_signal_11410 ;
    wire new_AGEMA_signal_11411 ;
    wire new_AGEMA_signal_11412 ;
    wire new_AGEMA_signal_11413 ;
    wire new_AGEMA_signal_11414 ;
    wire new_AGEMA_signal_11415 ;
    wire new_AGEMA_signal_11416 ;
    wire new_AGEMA_signal_11417 ;
    wire new_AGEMA_signal_11418 ;
    wire new_AGEMA_signal_11419 ;
    wire new_AGEMA_signal_11420 ;
    wire new_AGEMA_signal_11421 ;
    wire new_AGEMA_signal_11422 ;
    wire new_AGEMA_signal_11423 ;
    wire new_AGEMA_signal_11424 ;
    wire new_AGEMA_signal_11425 ;
    wire new_AGEMA_signal_11426 ;
    wire new_AGEMA_signal_11427 ;
    wire new_AGEMA_signal_11428 ;
    wire new_AGEMA_signal_11429 ;
    wire new_AGEMA_signal_11430 ;
    wire new_AGEMA_signal_11431 ;
    wire new_AGEMA_signal_11432 ;
    wire new_AGEMA_signal_11433 ;
    wire new_AGEMA_signal_11434 ;
    wire new_AGEMA_signal_11435 ;
    wire new_AGEMA_signal_11436 ;
    wire new_AGEMA_signal_11437 ;
    wire new_AGEMA_signal_11438 ;
    wire new_AGEMA_signal_11439 ;
    wire new_AGEMA_signal_11440 ;
    wire new_AGEMA_signal_11441 ;
    wire new_AGEMA_signal_11442 ;
    wire new_AGEMA_signal_11443 ;
    wire new_AGEMA_signal_11444 ;
    wire new_AGEMA_signal_11445 ;
    wire new_AGEMA_signal_11446 ;
    wire new_AGEMA_signal_11447 ;
    wire new_AGEMA_signal_11448 ;
    wire new_AGEMA_signal_11449 ;
    wire new_AGEMA_signal_11450 ;
    wire new_AGEMA_signal_11451 ;
    wire new_AGEMA_signal_11452 ;
    wire new_AGEMA_signal_11453 ;
    wire new_AGEMA_signal_11454 ;
    wire new_AGEMA_signal_11455 ;
    wire new_AGEMA_signal_11456 ;
    wire new_AGEMA_signal_11457 ;
    wire new_AGEMA_signal_11458 ;
    wire new_AGEMA_signal_11459 ;
    wire new_AGEMA_signal_11460 ;
    wire new_AGEMA_signal_11461 ;
    wire new_AGEMA_signal_11462 ;
    wire new_AGEMA_signal_11463 ;
    wire new_AGEMA_signal_11464 ;
    wire new_AGEMA_signal_11465 ;
    wire new_AGEMA_signal_11466 ;
    wire new_AGEMA_signal_11467 ;
    wire new_AGEMA_signal_11468 ;
    wire new_AGEMA_signal_11469 ;
    wire new_AGEMA_signal_11470 ;
    wire new_AGEMA_signal_11471 ;
    wire new_AGEMA_signal_11472 ;
    wire new_AGEMA_signal_11473 ;
    wire new_AGEMA_signal_11474 ;
    wire new_AGEMA_signal_11475 ;
    wire new_AGEMA_signal_11476 ;
    wire new_AGEMA_signal_11477 ;
    wire new_AGEMA_signal_11478 ;
    wire new_AGEMA_signal_11479 ;
    wire new_AGEMA_signal_11480 ;
    wire new_AGEMA_signal_11481 ;
    wire new_AGEMA_signal_11482 ;
    wire new_AGEMA_signal_11483 ;
    wire new_AGEMA_signal_11484 ;
    wire new_AGEMA_signal_11485 ;
    wire new_AGEMA_signal_11486 ;
    wire new_AGEMA_signal_11487 ;
    wire new_AGEMA_signal_11488 ;
    wire new_AGEMA_signal_11489 ;
    wire new_AGEMA_signal_11490 ;
    wire new_AGEMA_signal_11491 ;
    wire new_AGEMA_signal_11492 ;
    wire new_AGEMA_signal_11493 ;
    wire new_AGEMA_signal_11494 ;
    wire new_AGEMA_signal_11495 ;
    wire new_AGEMA_signal_11496 ;
    wire new_AGEMA_signal_11497 ;
    wire new_AGEMA_signal_11498 ;
    wire new_AGEMA_signal_11499 ;
    wire new_AGEMA_signal_11500 ;
    wire new_AGEMA_signal_11501 ;
    wire new_AGEMA_signal_11502 ;
    wire new_AGEMA_signal_11503 ;
    wire new_AGEMA_signal_11504 ;
    wire new_AGEMA_signal_11505 ;
    wire new_AGEMA_signal_11506 ;
    wire new_AGEMA_signal_11507 ;
    wire new_AGEMA_signal_11508 ;
    wire new_AGEMA_signal_11509 ;
    wire new_AGEMA_signal_11510 ;
    wire new_AGEMA_signal_11511 ;
    wire new_AGEMA_signal_11512 ;
    wire new_AGEMA_signal_11513 ;
    wire new_AGEMA_signal_11514 ;
    wire new_AGEMA_signal_11515 ;
    wire new_AGEMA_signal_11516 ;
    wire new_AGEMA_signal_11517 ;
    wire new_AGEMA_signal_11518 ;
    wire new_AGEMA_signal_11519 ;
    wire new_AGEMA_signal_11520 ;
    wire new_AGEMA_signal_11521 ;
    wire new_AGEMA_signal_11522 ;
    wire new_AGEMA_signal_11523 ;
    wire new_AGEMA_signal_11524 ;
    wire new_AGEMA_signal_11525 ;
    wire new_AGEMA_signal_11526 ;
    wire new_AGEMA_signal_11527 ;
    wire new_AGEMA_signal_11528 ;
    wire new_AGEMA_signal_11529 ;
    wire new_AGEMA_signal_11530 ;
    wire new_AGEMA_signal_11531 ;
    wire new_AGEMA_signal_11532 ;
    wire new_AGEMA_signal_11533 ;
    wire new_AGEMA_signal_11534 ;
    wire new_AGEMA_signal_11535 ;
    wire new_AGEMA_signal_11536 ;
    wire new_AGEMA_signal_11537 ;
    wire new_AGEMA_signal_11538 ;
    wire new_AGEMA_signal_11539 ;
    wire new_AGEMA_signal_11540 ;
    wire new_AGEMA_signal_11541 ;
    wire new_AGEMA_signal_11542 ;
    wire new_AGEMA_signal_11543 ;
    wire new_AGEMA_signal_11544 ;
    wire new_AGEMA_signal_11545 ;
    wire new_AGEMA_signal_11546 ;
    wire new_AGEMA_signal_11547 ;
    wire new_AGEMA_signal_11548 ;
    wire new_AGEMA_signal_11549 ;
    wire new_AGEMA_signal_11550 ;
    wire new_AGEMA_signal_11551 ;
    wire new_AGEMA_signal_11552 ;
    wire new_AGEMA_signal_11553 ;
    wire new_AGEMA_signal_11554 ;
    wire new_AGEMA_signal_11555 ;
    wire new_AGEMA_signal_11556 ;
    wire new_AGEMA_signal_11557 ;
    wire new_AGEMA_signal_11558 ;
    wire new_AGEMA_signal_11559 ;
    wire new_AGEMA_signal_11560 ;
    wire new_AGEMA_signal_11561 ;
    wire new_AGEMA_signal_11562 ;
    wire new_AGEMA_signal_11563 ;
    wire new_AGEMA_signal_11564 ;
    wire new_AGEMA_signal_11565 ;
    wire new_AGEMA_signal_11566 ;
    wire new_AGEMA_signal_11567 ;
    wire new_AGEMA_signal_11568 ;
    wire new_AGEMA_signal_11569 ;
    wire new_AGEMA_signal_11570 ;
    wire new_AGEMA_signal_11571 ;
    wire new_AGEMA_signal_11572 ;
    wire new_AGEMA_signal_11573 ;
    wire new_AGEMA_signal_11574 ;
    wire new_AGEMA_signal_11575 ;
    wire new_AGEMA_signal_11576 ;
    wire new_AGEMA_signal_11577 ;
    wire new_AGEMA_signal_11578 ;
    wire new_AGEMA_signal_11579 ;
    wire new_AGEMA_signal_11580 ;
    wire new_AGEMA_signal_11581 ;
    wire new_AGEMA_signal_11582 ;
    wire new_AGEMA_signal_11583 ;
    wire new_AGEMA_signal_11584 ;
    wire new_AGEMA_signal_11585 ;
    wire new_AGEMA_signal_11586 ;
    wire new_AGEMA_signal_11587 ;
    wire new_AGEMA_signal_11588 ;
    wire new_AGEMA_signal_11589 ;
    wire new_AGEMA_signal_11590 ;
    wire new_AGEMA_signal_11591 ;
    wire new_AGEMA_signal_11592 ;
    wire new_AGEMA_signal_11593 ;
    wire new_AGEMA_signal_11594 ;
    wire new_AGEMA_signal_11595 ;
    wire new_AGEMA_signal_11596 ;
    wire new_AGEMA_signal_11597 ;
    wire new_AGEMA_signal_11598 ;
    wire new_AGEMA_signal_11599 ;
    wire new_AGEMA_signal_11600 ;
    wire new_AGEMA_signal_11601 ;
    wire new_AGEMA_signal_11602 ;
    wire new_AGEMA_signal_11603 ;
    wire new_AGEMA_signal_11604 ;
    wire new_AGEMA_signal_11605 ;
    wire new_AGEMA_signal_11606 ;
    wire new_AGEMA_signal_11607 ;
    wire new_AGEMA_signal_11608 ;
    wire new_AGEMA_signal_11609 ;
    wire new_AGEMA_signal_11610 ;
    wire new_AGEMA_signal_11611 ;
    wire new_AGEMA_signal_11612 ;
    wire new_AGEMA_signal_11613 ;
    wire new_AGEMA_signal_11614 ;
    wire new_AGEMA_signal_11615 ;
    wire new_AGEMA_signal_11616 ;
    wire new_AGEMA_signal_11617 ;
    wire new_AGEMA_signal_11618 ;
    wire new_AGEMA_signal_11619 ;
    wire new_AGEMA_signal_11620 ;
    wire new_AGEMA_signal_11621 ;
    wire new_AGEMA_signal_11622 ;
    wire new_AGEMA_signal_11623 ;
    wire new_AGEMA_signal_11624 ;
    wire new_AGEMA_signal_11625 ;
    wire new_AGEMA_signal_11626 ;
    wire new_AGEMA_signal_11627 ;
    wire new_AGEMA_signal_11628 ;
    wire new_AGEMA_signal_11629 ;
    wire new_AGEMA_signal_11630 ;
    wire new_AGEMA_signal_11631 ;
    wire new_AGEMA_signal_11632 ;
    wire new_AGEMA_signal_11633 ;
    wire new_AGEMA_signal_11634 ;
    wire new_AGEMA_signal_11635 ;
    wire new_AGEMA_signal_11636 ;
    wire new_AGEMA_signal_11637 ;
    wire new_AGEMA_signal_11638 ;
    wire new_AGEMA_signal_11639 ;
    wire new_AGEMA_signal_11640 ;
    wire new_AGEMA_signal_11641 ;
    wire new_AGEMA_signal_11642 ;
    wire new_AGEMA_signal_11643 ;
    wire new_AGEMA_signal_11644 ;
    wire new_AGEMA_signal_11645 ;
    wire new_AGEMA_signal_11646 ;
    wire new_AGEMA_signal_11647 ;
    wire new_AGEMA_signal_11648 ;
    wire new_AGEMA_signal_11649 ;
    wire new_AGEMA_signal_11650 ;
    wire new_AGEMA_signal_11651 ;
    wire new_AGEMA_signal_11652 ;
    wire new_AGEMA_signal_11653 ;
    wire new_AGEMA_signal_11654 ;
    wire new_AGEMA_signal_11655 ;
    wire new_AGEMA_signal_11656 ;
    wire new_AGEMA_signal_11657 ;
    wire new_AGEMA_signal_11658 ;
    wire new_AGEMA_signal_11659 ;
    wire new_AGEMA_signal_11660 ;
    wire new_AGEMA_signal_11661 ;
    wire new_AGEMA_signal_11662 ;
    wire new_AGEMA_signal_11663 ;
    wire new_AGEMA_signal_11664 ;
    wire new_AGEMA_signal_11665 ;
    wire new_AGEMA_signal_11666 ;
    wire new_AGEMA_signal_11667 ;
    wire new_AGEMA_signal_11668 ;
    wire new_AGEMA_signal_11669 ;
    wire new_AGEMA_signal_11670 ;
    wire new_AGEMA_signal_11671 ;
    wire new_AGEMA_signal_11672 ;
    wire new_AGEMA_signal_11673 ;
    wire new_AGEMA_signal_11674 ;
    wire new_AGEMA_signal_11675 ;
    wire new_AGEMA_signal_11676 ;
    wire new_AGEMA_signal_11677 ;
    wire new_AGEMA_signal_11678 ;
    wire new_AGEMA_signal_11679 ;
    wire new_AGEMA_signal_11680 ;
    wire new_AGEMA_signal_11681 ;
    wire new_AGEMA_signal_11682 ;
    wire new_AGEMA_signal_11683 ;
    wire new_AGEMA_signal_11684 ;
    wire new_AGEMA_signal_11685 ;
    wire new_AGEMA_signal_11686 ;
    wire new_AGEMA_signal_11687 ;
    wire new_AGEMA_signal_11688 ;
    wire new_AGEMA_signal_11689 ;
    wire new_AGEMA_signal_11690 ;
    wire new_AGEMA_signal_11691 ;
    wire new_AGEMA_signal_11692 ;
    wire new_AGEMA_signal_11693 ;
    wire new_AGEMA_signal_11694 ;
    wire new_AGEMA_signal_11695 ;
    wire new_AGEMA_signal_11696 ;
    wire new_AGEMA_signal_11697 ;
    wire new_AGEMA_signal_11698 ;
    wire new_AGEMA_signal_11699 ;
    wire new_AGEMA_signal_11700 ;
    wire new_AGEMA_signal_11701 ;
    wire new_AGEMA_signal_11702 ;
    wire new_AGEMA_signal_11703 ;
    wire new_AGEMA_signal_11704 ;
    wire new_AGEMA_signal_11705 ;
    wire new_AGEMA_signal_11706 ;
    wire new_AGEMA_signal_11707 ;
    wire new_AGEMA_signal_11708 ;
    wire new_AGEMA_signal_11709 ;
    wire new_AGEMA_signal_11710 ;
    wire new_AGEMA_signal_11711 ;
    wire new_AGEMA_signal_11712 ;
    wire new_AGEMA_signal_11713 ;
    wire new_AGEMA_signal_11714 ;
    wire new_AGEMA_signal_11715 ;
    wire new_AGEMA_signal_11716 ;
    wire new_AGEMA_signal_11717 ;
    wire new_AGEMA_signal_11718 ;
    wire new_AGEMA_signal_11719 ;
    wire new_AGEMA_signal_11720 ;
    wire new_AGEMA_signal_11721 ;
    wire new_AGEMA_signal_11722 ;
    wire new_AGEMA_signal_11723 ;
    wire new_AGEMA_signal_11724 ;
    wire new_AGEMA_signal_11725 ;
    wire new_AGEMA_signal_11726 ;
    wire new_AGEMA_signal_11727 ;
    wire new_AGEMA_signal_11728 ;
    wire new_AGEMA_signal_11729 ;
    wire new_AGEMA_signal_11730 ;
    wire new_AGEMA_signal_11731 ;
    wire new_AGEMA_signal_11732 ;
    wire new_AGEMA_signal_11733 ;
    wire new_AGEMA_signal_11734 ;
    wire new_AGEMA_signal_11735 ;
    wire new_AGEMA_signal_11736 ;
    wire new_AGEMA_signal_11737 ;
    wire new_AGEMA_signal_11738 ;
    wire new_AGEMA_signal_11739 ;
    wire new_AGEMA_signal_11740 ;
    wire new_AGEMA_signal_11741 ;
    wire new_AGEMA_signal_11742 ;
    wire new_AGEMA_signal_11743 ;
    wire new_AGEMA_signal_11744 ;
    wire new_AGEMA_signal_11745 ;
    wire new_AGEMA_signal_11746 ;
    wire new_AGEMA_signal_11747 ;
    wire new_AGEMA_signal_11748 ;
    wire new_AGEMA_signal_11749 ;
    wire new_AGEMA_signal_11750 ;
    wire new_AGEMA_signal_11751 ;
    wire new_AGEMA_signal_11752 ;
    wire new_AGEMA_signal_11753 ;
    wire new_AGEMA_signal_11754 ;
    wire new_AGEMA_signal_11755 ;
    wire new_AGEMA_signal_11756 ;
    wire new_AGEMA_signal_11757 ;
    wire new_AGEMA_signal_11758 ;
    wire new_AGEMA_signal_11759 ;
    wire new_AGEMA_signal_11760 ;
    wire new_AGEMA_signal_11761 ;
    wire new_AGEMA_signal_11762 ;
    wire new_AGEMA_signal_11763 ;
    wire new_AGEMA_signal_11764 ;
    wire new_AGEMA_signal_11765 ;
    wire new_AGEMA_signal_11766 ;
    wire new_AGEMA_signal_11767 ;
    wire new_AGEMA_signal_11768 ;
    wire new_AGEMA_signal_11769 ;
    wire new_AGEMA_signal_11770 ;
    wire new_AGEMA_signal_11771 ;
    wire new_AGEMA_signal_11772 ;
    wire new_AGEMA_signal_11773 ;
    wire new_AGEMA_signal_11774 ;
    wire new_AGEMA_signal_11775 ;
    wire new_AGEMA_signal_11776 ;
    wire new_AGEMA_signal_11777 ;
    wire new_AGEMA_signal_11778 ;
    wire new_AGEMA_signal_11779 ;
    wire new_AGEMA_signal_11780 ;
    wire new_AGEMA_signal_11781 ;
    wire new_AGEMA_signal_11782 ;
    wire new_AGEMA_signal_11783 ;
    wire new_AGEMA_signal_11784 ;
    wire new_AGEMA_signal_11785 ;
    wire new_AGEMA_signal_11786 ;
    wire new_AGEMA_signal_11787 ;
    wire new_AGEMA_signal_11788 ;
    wire new_AGEMA_signal_11789 ;
    wire new_AGEMA_signal_11790 ;
    wire new_AGEMA_signal_11791 ;
    wire new_AGEMA_signal_11792 ;
    wire new_AGEMA_signal_11793 ;
    wire new_AGEMA_signal_11794 ;
    wire new_AGEMA_signal_11795 ;
    wire new_AGEMA_signal_11796 ;
    wire new_AGEMA_signal_11797 ;
    wire new_AGEMA_signal_11798 ;
    wire new_AGEMA_signal_11799 ;
    wire new_AGEMA_signal_11800 ;
    wire new_AGEMA_signal_11801 ;
    wire new_AGEMA_signal_11802 ;
    wire new_AGEMA_signal_11803 ;
    wire new_AGEMA_signal_11804 ;
    wire new_AGEMA_signal_11805 ;
    wire new_AGEMA_signal_11806 ;
    wire new_AGEMA_signal_11807 ;
    wire new_AGEMA_signal_11808 ;
    wire new_AGEMA_signal_11809 ;
    wire new_AGEMA_signal_11810 ;
    wire new_AGEMA_signal_11811 ;
    wire new_AGEMA_signal_11812 ;
    wire new_AGEMA_signal_11813 ;
    wire new_AGEMA_signal_11814 ;
    wire new_AGEMA_signal_11815 ;
    wire new_AGEMA_signal_11816 ;
    wire new_AGEMA_signal_11817 ;
    wire new_AGEMA_signal_11818 ;
    wire new_AGEMA_signal_11819 ;
    wire new_AGEMA_signal_11820 ;
    wire new_AGEMA_signal_11821 ;
    wire new_AGEMA_signal_11822 ;
    wire new_AGEMA_signal_11823 ;
    wire new_AGEMA_signal_11824 ;
    wire new_AGEMA_signal_11825 ;
    wire new_AGEMA_signal_11826 ;
    wire new_AGEMA_signal_11827 ;
    wire new_AGEMA_signal_11828 ;
    wire new_AGEMA_signal_11829 ;
    wire new_AGEMA_signal_11830 ;
    wire new_AGEMA_signal_11831 ;
    wire new_AGEMA_signal_11832 ;
    wire new_AGEMA_signal_11833 ;
    wire new_AGEMA_signal_11834 ;
    wire new_AGEMA_signal_11835 ;
    wire new_AGEMA_signal_11836 ;
    wire new_AGEMA_signal_11837 ;
    wire new_AGEMA_signal_11838 ;
    wire new_AGEMA_signal_11839 ;
    wire new_AGEMA_signal_11840 ;
    wire new_AGEMA_signal_11841 ;
    wire new_AGEMA_signal_11842 ;
    wire new_AGEMA_signal_11843 ;
    wire new_AGEMA_signal_11844 ;
    wire new_AGEMA_signal_11845 ;
    wire new_AGEMA_signal_11846 ;
    wire new_AGEMA_signal_11847 ;
    wire new_AGEMA_signal_11848 ;
    wire new_AGEMA_signal_11849 ;
    wire new_AGEMA_signal_11850 ;
    wire new_AGEMA_signal_11851 ;
    wire new_AGEMA_signal_11852 ;
    wire new_AGEMA_signal_11853 ;
    wire new_AGEMA_signal_11854 ;
    wire new_AGEMA_signal_11855 ;
    wire new_AGEMA_signal_11856 ;
    wire new_AGEMA_signal_11857 ;
    wire new_AGEMA_signal_11858 ;
    wire new_AGEMA_signal_11859 ;
    wire new_AGEMA_signal_11860 ;
    wire new_AGEMA_signal_11861 ;
    wire new_AGEMA_signal_11862 ;
    wire new_AGEMA_signal_11863 ;
    wire new_AGEMA_signal_11864 ;
    wire new_AGEMA_signal_11865 ;
    wire new_AGEMA_signal_11866 ;
    wire new_AGEMA_signal_11867 ;
    wire new_AGEMA_signal_11868 ;
    wire new_AGEMA_signal_11869 ;
    wire new_AGEMA_signal_11870 ;
    wire new_AGEMA_signal_11871 ;
    wire new_AGEMA_signal_11872 ;
    wire new_AGEMA_signal_11873 ;
    wire new_AGEMA_signal_11874 ;
    wire new_AGEMA_signal_11875 ;
    wire new_AGEMA_signal_11876 ;
    wire new_AGEMA_signal_11877 ;
    wire new_AGEMA_signal_11878 ;
    wire new_AGEMA_signal_11879 ;
    wire new_AGEMA_signal_11880 ;
    wire new_AGEMA_signal_11881 ;
    wire new_AGEMA_signal_11882 ;
    wire new_AGEMA_signal_11883 ;
    wire new_AGEMA_signal_11884 ;
    wire new_AGEMA_signal_11885 ;
    wire new_AGEMA_signal_11886 ;
    wire new_AGEMA_signal_11887 ;
    wire new_AGEMA_signal_11888 ;
    wire new_AGEMA_signal_11889 ;
    wire new_AGEMA_signal_11890 ;
    wire new_AGEMA_signal_11891 ;
    wire new_AGEMA_signal_11892 ;
    wire new_AGEMA_signal_11893 ;
    wire new_AGEMA_signal_11894 ;
    wire new_AGEMA_signal_11895 ;
    wire new_AGEMA_signal_11896 ;
    wire new_AGEMA_signal_11897 ;
    wire new_AGEMA_signal_11898 ;
    wire new_AGEMA_signal_11899 ;
    wire new_AGEMA_signal_11900 ;
    wire new_AGEMA_signal_11901 ;
    wire new_AGEMA_signal_11902 ;
    wire new_AGEMA_signal_11903 ;
    wire new_AGEMA_signal_11904 ;
    wire new_AGEMA_signal_11905 ;
    wire new_AGEMA_signal_11906 ;
    wire new_AGEMA_signal_11907 ;
    wire new_AGEMA_signal_11908 ;
    wire new_AGEMA_signal_11909 ;
    wire new_AGEMA_signal_11910 ;
    wire new_AGEMA_signal_11911 ;
    wire new_AGEMA_signal_11912 ;
    wire new_AGEMA_signal_11913 ;
    wire new_AGEMA_signal_11914 ;
    wire new_AGEMA_signal_11915 ;
    wire new_AGEMA_signal_11916 ;
    wire new_AGEMA_signal_11917 ;
    wire new_AGEMA_signal_11918 ;
    wire new_AGEMA_signal_11919 ;
    wire new_AGEMA_signal_11920 ;
    wire new_AGEMA_signal_11921 ;
    wire new_AGEMA_signal_11922 ;
    wire new_AGEMA_signal_11923 ;
    wire new_AGEMA_signal_11924 ;
    wire new_AGEMA_signal_11925 ;
    wire new_AGEMA_signal_11926 ;
    wire new_AGEMA_signal_11927 ;
    wire new_AGEMA_signal_11928 ;
    wire new_AGEMA_signal_11929 ;
    wire new_AGEMA_signal_11930 ;
    wire new_AGEMA_signal_11931 ;
    wire new_AGEMA_signal_11932 ;
    wire new_AGEMA_signal_11933 ;
    wire new_AGEMA_signal_11934 ;
    wire new_AGEMA_signal_11935 ;
    wire new_AGEMA_signal_11936 ;
    wire new_AGEMA_signal_11937 ;
    wire new_AGEMA_signal_11938 ;
    wire new_AGEMA_signal_11939 ;
    wire new_AGEMA_signal_11940 ;
    wire new_AGEMA_signal_11941 ;
    wire new_AGEMA_signal_11942 ;
    wire new_AGEMA_signal_11943 ;
    wire new_AGEMA_signal_11944 ;
    wire new_AGEMA_signal_11945 ;
    wire new_AGEMA_signal_11946 ;
    wire new_AGEMA_signal_11947 ;
    wire new_AGEMA_signal_11948 ;
    wire new_AGEMA_signal_11949 ;
    wire new_AGEMA_signal_11950 ;
    wire new_AGEMA_signal_11951 ;
    wire new_AGEMA_signal_11952 ;
    wire new_AGEMA_signal_11953 ;
    wire new_AGEMA_signal_11954 ;
    wire new_AGEMA_signal_11955 ;
    wire new_AGEMA_signal_11956 ;
    wire new_AGEMA_signal_11957 ;
    wire new_AGEMA_signal_11958 ;
    wire new_AGEMA_signal_11959 ;
    wire new_AGEMA_signal_11960 ;
    wire new_AGEMA_signal_11961 ;
    wire new_AGEMA_signal_11962 ;
    wire new_AGEMA_signal_11963 ;
    wire new_AGEMA_signal_11964 ;
    wire new_AGEMA_signal_11965 ;
    wire new_AGEMA_signal_11966 ;
    wire new_AGEMA_signal_11967 ;
    wire new_AGEMA_signal_11968 ;
    wire new_AGEMA_signal_11969 ;
    wire new_AGEMA_signal_11970 ;
    wire new_AGEMA_signal_11971 ;
    wire new_AGEMA_signal_11972 ;
    wire new_AGEMA_signal_11973 ;
    wire new_AGEMA_signal_11974 ;
    wire new_AGEMA_signal_11975 ;
    wire new_AGEMA_signal_11976 ;
    wire new_AGEMA_signal_11977 ;
    wire new_AGEMA_signal_11978 ;
    wire new_AGEMA_signal_11979 ;
    wire new_AGEMA_signal_11980 ;
    wire new_AGEMA_signal_11981 ;
    wire new_AGEMA_signal_11982 ;
    wire new_AGEMA_signal_11983 ;
    wire new_AGEMA_signal_11984 ;
    wire new_AGEMA_signal_11985 ;
    wire new_AGEMA_signal_11986 ;
    wire new_AGEMA_signal_11987 ;
    wire new_AGEMA_signal_11988 ;
    wire new_AGEMA_signal_11989 ;
    wire new_AGEMA_signal_11990 ;
    wire new_AGEMA_signal_11991 ;
    wire new_AGEMA_signal_11992 ;
    wire new_AGEMA_signal_11993 ;
    wire new_AGEMA_signal_11994 ;
    wire new_AGEMA_signal_11995 ;
    wire new_AGEMA_signal_11996 ;
    wire new_AGEMA_signal_11997 ;
    wire new_AGEMA_signal_11998 ;
    wire new_AGEMA_signal_11999 ;
    wire new_AGEMA_signal_12000 ;
    wire new_AGEMA_signal_12001 ;
    wire new_AGEMA_signal_12002 ;
    wire new_AGEMA_signal_12003 ;
    wire new_AGEMA_signal_12004 ;
    wire new_AGEMA_signal_12005 ;
    wire new_AGEMA_signal_12006 ;
    wire new_AGEMA_signal_12007 ;
    wire new_AGEMA_signal_12008 ;
    wire new_AGEMA_signal_12009 ;
    wire new_AGEMA_signal_12010 ;
    wire new_AGEMA_signal_12011 ;
    wire new_AGEMA_signal_12012 ;
    wire new_AGEMA_signal_12013 ;
    wire new_AGEMA_signal_12014 ;
    wire new_AGEMA_signal_12015 ;
    wire new_AGEMA_signal_12016 ;
    wire new_AGEMA_signal_12017 ;
    wire new_AGEMA_signal_12018 ;
    wire new_AGEMA_signal_12019 ;
    wire new_AGEMA_signal_12020 ;
    wire new_AGEMA_signal_12021 ;
    wire new_AGEMA_signal_12022 ;
    wire new_AGEMA_signal_12023 ;
    wire new_AGEMA_signal_12024 ;
    wire new_AGEMA_signal_12025 ;
    wire new_AGEMA_signal_12026 ;
    wire new_AGEMA_signal_12027 ;
    wire new_AGEMA_signal_12028 ;
    wire new_AGEMA_signal_12029 ;
    wire new_AGEMA_signal_12030 ;
    wire new_AGEMA_signal_12031 ;
    wire new_AGEMA_signal_12032 ;
    wire new_AGEMA_signal_12033 ;
    wire new_AGEMA_signal_12034 ;
    wire new_AGEMA_signal_12035 ;
    wire new_AGEMA_signal_12036 ;
    wire new_AGEMA_signal_12037 ;
    wire new_AGEMA_signal_12038 ;
    wire new_AGEMA_signal_12039 ;
    wire new_AGEMA_signal_12040 ;
    wire new_AGEMA_signal_12041 ;
    wire new_AGEMA_signal_12042 ;
    wire new_AGEMA_signal_12043 ;
    wire new_AGEMA_signal_12044 ;
    wire new_AGEMA_signal_12045 ;
    wire new_AGEMA_signal_12046 ;
    wire new_AGEMA_signal_12047 ;
    wire new_AGEMA_signal_12048 ;
    wire new_AGEMA_signal_12049 ;
    wire new_AGEMA_signal_12050 ;
    wire new_AGEMA_signal_12051 ;
    wire new_AGEMA_signal_12052 ;
    wire new_AGEMA_signal_12053 ;
    wire new_AGEMA_signal_12054 ;
    wire new_AGEMA_signal_12055 ;
    wire new_AGEMA_signal_12056 ;
    wire new_AGEMA_signal_12057 ;
    wire new_AGEMA_signal_12058 ;
    wire new_AGEMA_signal_12059 ;
    wire new_AGEMA_signal_12060 ;
    wire new_AGEMA_signal_12061 ;
    wire new_AGEMA_signal_12062 ;
    wire new_AGEMA_signal_12063 ;
    wire new_AGEMA_signal_12064 ;
    wire new_AGEMA_signal_12065 ;
    wire new_AGEMA_signal_12066 ;
    wire new_AGEMA_signal_12067 ;
    wire new_AGEMA_signal_12068 ;
    wire new_AGEMA_signal_12069 ;
    wire new_AGEMA_signal_12070 ;
    wire new_AGEMA_signal_12071 ;
    wire new_AGEMA_signal_12072 ;
    wire new_AGEMA_signal_12073 ;
    wire new_AGEMA_signal_12074 ;
    wire new_AGEMA_signal_12075 ;
    wire new_AGEMA_signal_12076 ;
    wire new_AGEMA_signal_12077 ;
    wire new_AGEMA_signal_12078 ;
    wire new_AGEMA_signal_12079 ;
    wire new_AGEMA_signal_12080 ;
    wire new_AGEMA_signal_12081 ;
    wire new_AGEMA_signal_12082 ;
    wire new_AGEMA_signal_12083 ;
    wire new_AGEMA_signal_12084 ;
    wire new_AGEMA_signal_12085 ;
    wire new_AGEMA_signal_12086 ;
    wire new_AGEMA_signal_12087 ;
    wire new_AGEMA_signal_12088 ;
    wire new_AGEMA_signal_12089 ;
    wire new_AGEMA_signal_12090 ;
    wire new_AGEMA_signal_12091 ;
    wire new_AGEMA_signal_12092 ;
    wire new_AGEMA_signal_12093 ;
    wire new_AGEMA_signal_12094 ;
    wire new_AGEMA_signal_12095 ;
    wire new_AGEMA_signal_12096 ;
    wire new_AGEMA_signal_12097 ;
    wire new_AGEMA_signal_12098 ;
    wire new_AGEMA_signal_12099 ;
    wire new_AGEMA_signal_12100 ;
    wire new_AGEMA_signal_12101 ;
    wire new_AGEMA_signal_12102 ;
    wire new_AGEMA_signal_12103 ;
    wire new_AGEMA_signal_12104 ;
    wire new_AGEMA_signal_12105 ;
    wire new_AGEMA_signal_12106 ;
    wire new_AGEMA_signal_12107 ;
    wire new_AGEMA_signal_12108 ;
    wire new_AGEMA_signal_12109 ;
    wire new_AGEMA_signal_12110 ;
    wire new_AGEMA_signal_12111 ;
    wire new_AGEMA_signal_12112 ;
    wire new_AGEMA_signal_12113 ;
    wire new_AGEMA_signal_12114 ;
    wire new_AGEMA_signal_12115 ;
    wire new_AGEMA_signal_12116 ;
    wire new_AGEMA_signal_12117 ;
    wire new_AGEMA_signal_12118 ;
    wire new_AGEMA_signal_12119 ;
    wire new_AGEMA_signal_12120 ;
    wire new_AGEMA_signal_12121 ;
    wire new_AGEMA_signal_12122 ;
    wire new_AGEMA_signal_12123 ;
    wire new_AGEMA_signal_12124 ;
    wire new_AGEMA_signal_12125 ;
    wire new_AGEMA_signal_12126 ;
    wire new_AGEMA_signal_12127 ;
    wire new_AGEMA_signal_12128 ;
    wire new_AGEMA_signal_12129 ;
    wire new_AGEMA_signal_12130 ;
    wire new_AGEMA_signal_12131 ;
    wire new_AGEMA_signal_12132 ;
    wire new_AGEMA_signal_12133 ;
    wire new_AGEMA_signal_12134 ;
    wire new_AGEMA_signal_12135 ;
    wire new_AGEMA_signal_12136 ;
    wire new_AGEMA_signal_12137 ;
    wire new_AGEMA_signal_12138 ;
    wire new_AGEMA_signal_12139 ;
    wire new_AGEMA_signal_12140 ;
    wire new_AGEMA_signal_12141 ;
    wire new_AGEMA_signal_12142 ;
    wire new_AGEMA_signal_12143 ;
    wire new_AGEMA_signal_12144 ;
    wire new_AGEMA_signal_12145 ;
    wire new_AGEMA_signal_12146 ;
    wire new_AGEMA_signal_12147 ;
    wire new_AGEMA_signal_12148 ;
    wire new_AGEMA_signal_12149 ;
    wire new_AGEMA_signal_12150 ;
    wire new_AGEMA_signal_12151 ;
    wire new_AGEMA_signal_12152 ;
    wire new_AGEMA_signal_12153 ;
    wire new_AGEMA_signal_12154 ;
    wire new_AGEMA_signal_12155 ;
    wire new_AGEMA_signal_12156 ;
    wire new_AGEMA_signal_12157 ;
    wire new_AGEMA_signal_12158 ;
    wire new_AGEMA_signal_12159 ;
    wire new_AGEMA_signal_12160 ;
    wire new_AGEMA_signal_12161 ;
    wire new_AGEMA_signal_12162 ;
    wire new_AGEMA_signal_12163 ;
    wire new_AGEMA_signal_12164 ;
    wire new_AGEMA_signal_12165 ;
    wire new_AGEMA_signal_12166 ;
    wire new_AGEMA_signal_12167 ;
    wire new_AGEMA_signal_12168 ;
    wire new_AGEMA_signal_12169 ;
    wire new_AGEMA_signal_12170 ;
    wire new_AGEMA_signal_12171 ;
    wire new_AGEMA_signal_12172 ;
    wire new_AGEMA_signal_12173 ;
    wire new_AGEMA_signal_12174 ;
    wire new_AGEMA_signal_12175 ;
    wire new_AGEMA_signal_12176 ;
    wire new_AGEMA_signal_12177 ;
    wire new_AGEMA_signal_12178 ;
    wire new_AGEMA_signal_12179 ;
    wire new_AGEMA_signal_12180 ;
    wire new_AGEMA_signal_12181 ;
    wire new_AGEMA_signal_12182 ;
    wire new_AGEMA_signal_12183 ;
    wire new_AGEMA_signal_12184 ;
    wire new_AGEMA_signal_12185 ;
    wire new_AGEMA_signal_12186 ;
    wire new_AGEMA_signal_12187 ;
    wire new_AGEMA_signal_12188 ;
    wire new_AGEMA_signal_12189 ;
    wire new_AGEMA_signal_12190 ;
    wire new_AGEMA_signal_12191 ;
    wire new_AGEMA_signal_12192 ;
    wire new_AGEMA_signal_12193 ;
    wire new_AGEMA_signal_12194 ;
    wire new_AGEMA_signal_12195 ;
    wire new_AGEMA_signal_12196 ;
    wire new_AGEMA_signal_12197 ;
    wire new_AGEMA_signal_12198 ;
    wire new_AGEMA_signal_12199 ;
    wire new_AGEMA_signal_12200 ;
    wire new_AGEMA_signal_12201 ;
    wire new_AGEMA_signal_12202 ;
    wire new_AGEMA_signal_12203 ;
    wire new_AGEMA_signal_12204 ;
    wire new_AGEMA_signal_12205 ;
    wire new_AGEMA_signal_12206 ;
    wire new_AGEMA_signal_12207 ;
    wire new_AGEMA_signal_12208 ;
    wire new_AGEMA_signal_12209 ;
    wire new_AGEMA_signal_12210 ;
    wire new_AGEMA_signal_12211 ;
    wire new_AGEMA_signal_12212 ;
    wire new_AGEMA_signal_12213 ;
    wire new_AGEMA_signal_12214 ;
    wire new_AGEMA_signal_12215 ;
    wire new_AGEMA_signal_12216 ;
    wire new_AGEMA_signal_12217 ;
    wire new_AGEMA_signal_12218 ;
    wire new_AGEMA_signal_12219 ;
    wire new_AGEMA_signal_12220 ;
    wire new_AGEMA_signal_12221 ;
    wire new_AGEMA_signal_12222 ;
    wire new_AGEMA_signal_12223 ;
    wire new_AGEMA_signal_12224 ;
    wire new_AGEMA_signal_12225 ;
    wire new_AGEMA_signal_12226 ;
    wire new_AGEMA_signal_12227 ;
    wire new_AGEMA_signal_12228 ;
    wire new_AGEMA_signal_12229 ;
    wire new_AGEMA_signal_12230 ;
    wire new_AGEMA_signal_12231 ;
    wire new_AGEMA_signal_12232 ;
    wire new_AGEMA_signal_12233 ;
    wire new_AGEMA_signal_12234 ;
    wire new_AGEMA_signal_12235 ;
    wire new_AGEMA_signal_12236 ;
    wire new_AGEMA_signal_12237 ;
    wire new_AGEMA_signal_12238 ;
    wire new_AGEMA_signal_12239 ;
    wire new_AGEMA_signal_12240 ;
    wire new_AGEMA_signal_12241 ;
    wire new_AGEMA_signal_12242 ;
    wire new_AGEMA_signal_12243 ;
    wire new_AGEMA_signal_12244 ;
    wire new_AGEMA_signal_12245 ;
    wire new_AGEMA_signal_12246 ;
    wire new_AGEMA_signal_12247 ;
    wire new_AGEMA_signal_12248 ;
    wire new_AGEMA_signal_12249 ;
    wire new_AGEMA_signal_12250 ;
    wire new_AGEMA_signal_12251 ;
    wire new_AGEMA_signal_12252 ;
    wire new_AGEMA_signal_12253 ;
    wire new_AGEMA_signal_12254 ;
    wire new_AGEMA_signal_12255 ;
    wire new_AGEMA_signal_12256 ;
    wire new_AGEMA_signal_12257 ;
    wire new_AGEMA_signal_12258 ;
    wire new_AGEMA_signal_12259 ;
    wire new_AGEMA_signal_12260 ;
    wire new_AGEMA_signal_12261 ;
    wire new_AGEMA_signal_12262 ;
    wire new_AGEMA_signal_12263 ;
    wire new_AGEMA_signal_12264 ;
    wire new_AGEMA_signal_12265 ;
    wire new_AGEMA_signal_12266 ;
    wire new_AGEMA_signal_12267 ;
    wire new_AGEMA_signal_12268 ;
    wire new_AGEMA_signal_12269 ;
    wire new_AGEMA_signal_12270 ;
    wire new_AGEMA_signal_12271 ;
    wire new_AGEMA_signal_12272 ;
    wire new_AGEMA_signal_12273 ;
    wire new_AGEMA_signal_12274 ;
    wire new_AGEMA_signal_12275 ;
    wire new_AGEMA_signal_12276 ;
    wire new_AGEMA_signal_12277 ;
    wire new_AGEMA_signal_12278 ;
    wire new_AGEMA_signal_12279 ;
    wire new_AGEMA_signal_12280 ;
    wire new_AGEMA_signal_12281 ;
    wire new_AGEMA_signal_12282 ;
    wire new_AGEMA_signal_12283 ;
    wire new_AGEMA_signal_12284 ;
    wire new_AGEMA_signal_12285 ;
    wire new_AGEMA_signal_12286 ;
    wire new_AGEMA_signal_12287 ;
    wire new_AGEMA_signal_12288 ;
    wire new_AGEMA_signal_12289 ;
    wire new_AGEMA_signal_12290 ;
    wire new_AGEMA_signal_12291 ;
    wire new_AGEMA_signal_12292 ;
    wire new_AGEMA_signal_12293 ;
    wire new_AGEMA_signal_12294 ;
    wire new_AGEMA_signal_12295 ;
    wire new_AGEMA_signal_12296 ;
    wire new_AGEMA_signal_12297 ;
    wire new_AGEMA_signal_12298 ;
    wire new_AGEMA_signal_12299 ;
    wire new_AGEMA_signal_12300 ;
    wire new_AGEMA_signal_12301 ;
    wire new_AGEMA_signal_12302 ;
    wire new_AGEMA_signal_12303 ;
    wire new_AGEMA_signal_12304 ;
    wire new_AGEMA_signal_12305 ;
    wire new_AGEMA_signal_12306 ;
    wire new_AGEMA_signal_12307 ;
    wire new_AGEMA_signal_12308 ;
    wire new_AGEMA_signal_12309 ;
    wire new_AGEMA_signal_12310 ;
    wire new_AGEMA_signal_12311 ;
    wire new_AGEMA_signal_12312 ;
    wire new_AGEMA_signal_12313 ;
    wire new_AGEMA_signal_12314 ;
    wire new_AGEMA_signal_12315 ;
    wire new_AGEMA_signal_12316 ;
    wire new_AGEMA_signal_12317 ;
    wire new_AGEMA_signal_12318 ;
    wire new_AGEMA_signal_12319 ;
    wire new_AGEMA_signal_12320 ;
    wire new_AGEMA_signal_12321 ;
    wire new_AGEMA_signal_12322 ;
    wire new_AGEMA_signal_12323 ;
    wire new_AGEMA_signal_12324 ;
    wire new_AGEMA_signal_12325 ;
    wire new_AGEMA_signal_12326 ;
    wire new_AGEMA_signal_12327 ;
    wire new_AGEMA_signal_12328 ;
    wire new_AGEMA_signal_12329 ;
    wire new_AGEMA_signal_12330 ;
    wire new_AGEMA_signal_12331 ;
    wire new_AGEMA_signal_12332 ;
    wire new_AGEMA_signal_12333 ;
    wire new_AGEMA_signal_12334 ;
    wire new_AGEMA_signal_12335 ;
    wire new_AGEMA_signal_12336 ;
    wire new_AGEMA_signal_12337 ;
    wire new_AGEMA_signal_12338 ;
    wire new_AGEMA_signal_12339 ;
    wire new_AGEMA_signal_12340 ;
    wire new_AGEMA_signal_12341 ;
    wire new_AGEMA_signal_12342 ;
    wire new_AGEMA_signal_12343 ;
    wire new_AGEMA_signal_12344 ;
    wire new_AGEMA_signal_12345 ;
    wire new_AGEMA_signal_12346 ;
    wire new_AGEMA_signal_12347 ;
    wire new_AGEMA_signal_12348 ;
    wire new_AGEMA_signal_12349 ;
    wire new_AGEMA_signal_12350 ;
    wire new_AGEMA_signal_12351 ;
    wire new_AGEMA_signal_12352 ;
    wire new_AGEMA_signal_12353 ;
    wire new_AGEMA_signal_12354 ;
    wire new_AGEMA_signal_12355 ;
    wire new_AGEMA_signal_12356 ;
    wire new_AGEMA_signal_12357 ;
    wire new_AGEMA_signal_12358 ;
    wire new_AGEMA_signal_12359 ;
    wire new_AGEMA_signal_12360 ;
    wire new_AGEMA_signal_12361 ;
    wire new_AGEMA_signal_12362 ;
    wire new_AGEMA_signal_12363 ;
    wire new_AGEMA_signal_12364 ;
    wire new_AGEMA_signal_12365 ;
    wire new_AGEMA_signal_12366 ;
    wire new_AGEMA_signal_12367 ;
    wire new_AGEMA_signal_12368 ;
    wire new_AGEMA_signal_12369 ;
    wire new_AGEMA_signal_12370 ;
    wire new_AGEMA_signal_12371 ;
    wire new_AGEMA_signal_12372 ;
    wire new_AGEMA_signal_12373 ;
    wire new_AGEMA_signal_12374 ;
    wire new_AGEMA_signal_12375 ;
    wire new_AGEMA_signal_12376 ;
    wire new_AGEMA_signal_12377 ;
    wire new_AGEMA_signal_12378 ;
    wire new_AGEMA_signal_12379 ;
    wire new_AGEMA_signal_12380 ;
    wire new_AGEMA_signal_12381 ;
    wire new_AGEMA_signal_12382 ;
    wire new_AGEMA_signal_12383 ;
    wire new_AGEMA_signal_12384 ;
    wire new_AGEMA_signal_12385 ;
    wire new_AGEMA_signal_12386 ;
    wire new_AGEMA_signal_12387 ;
    wire new_AGEMA_signal_12388 ;
    wire new_AGEMA_signal_12389 ;
    wire new_AGEMA_signal_12390 ;
    wire new_AGEMA_signal_12391 ;
    wire new_AGEMA_signal_12392 ;
    wire new_AGEMA_signal_12393 ;
    wire new_AGEMA_signal_12394 ;
    wire new_AGEMA_signal_12395 ;
    wire new_AGEMA_signal_12396 ;
    wire new_AGEMA_signal_12397 ;
    wire new_AGEMA_signal_12398 ;
    wire new_AGEMA_signal_12399 ;
    wire new_AGEMA_signal_12400 ;
    wire new_AGEMA_signal_12401 ;
    wire new_AGEMA_signal_12402 ;
    wire new_AGEMA_signal_12403 ;
    wire new_AGEMA_signal_12404 ;
    wire new_AGEMA_signal_12405 ;
    wire new_AGEMA_signal_12406 ;
    wire new_AGEMA_signal_12407 ;
    wire new_AGEMA_signal_12408 ;
    wire new_AGEMA_signal_12409 ;
    wire new_AGEMA_signal_12410 ;
    wire new_AGEMA_signal_12411 ;
    wire new_AGEMA_signal_12412 ;
    wire new_AGEMA_signal_12413 ;
    wire new_AGEMA_signal_12414 ;
    wire new_AGEMA_signal_12415 ;
    wire new_AGEMA_signal_12416 ;
    wire new_AGEMA_signal_12417 ;
    wire new_AGEMA_signal_12418 ;
    wire new_AGEMA_signal_12419 ;
    wire new_AGEMA_signal_12420 ;
    wire new_AGEMA_signal_12421 ;
    wire new_AGEMA_signal_12422 ;
    wire new_AGEMA_signal_12423 ;
    wire new_AGEMA_signal_12424 ;
    wire new_AGEMA_signal_12425 ;
    wire new_AGEMA_signal_12426 ;
    wire new_AGEMA_signal_12427 ;
    wire new_AGEMA_signal_12428 ;
    wire new_AGEMA_signal_12429 ;
    wire new_AGEMA_signal_12430 ;
    wire new_AGEMA_signal_12431 ;
    wire new_AGEMA_signal_12432 ;
    wire new_AGEMA_signal_12433 ;
    wire new_AGEMA_signal_12434 ;
    wire new_AGEMA_signal_12435 ;
    wire new_AGEMA_signal_12436 ;
    wire new_AGEMA_signal_12437 ;
    wire new_AGEMA_signal_12438 ;
    wire new_AGEMA_signal_12439 ;
    wire new_AGEMA_signal_12440 ;
    wire new_AGEMA_signal_12441 ;
    wire new_AGEMA_signal_12442 ;
    wire new_AGEMA_signal_12443 ;
    wire new_AGEMA_signal_12444 ;
    wire new_AGEMA_signal_12445 ;
    wire new_AGEMA_signal_12446 ;
    wire new_AGEMA_signal_12447 ;
    wire new_AGEMA_signal_12448 ;
    wire new_AGEMA_signal_12449 ;
    wire new_AGEMA_signal_12450 ;
    wire new_AGEMA_signal_12451 ;
    wire new_AGEMA_signal_12452 ;
    wire new_AGEMA_signal_12453 ;
    wire new_AGEMA_signal_12454 ;
    wire new_AGEMA_signal_12455 ;
    wire new_AGEMA_signal_12456 ;
    wire new_AGEMA_signal_12457 ;
    wire new_AGEMA_signal_12458 ;
    wire new_AGEMA_signal_12459 ;
    wire new_AGEMA_signal_12460 ;
    wire new_AGEMA_signal_12461 ;
    wire new_AGEMA_signal_12462 ;
    wire new_AGEMA_signal_12463 ;
    wire new_AGEMA_signal_12464 ;
    wire new_AGEMA_signal_12465 ;
    wire new_AGEMA_signal_12466 ;
    wire new_AGEMA_signal_12467 ;
    wire new_AGEMA_signal_12468 ;
    wire new_AGEMA_signal_12469 ;
    wire new_AGEMA_signal_12470 ;
    wire new_AGEMA_signal_12471 ;
    wire new_AGEMA_signal_12472 ;
    wire new_AGEMA_signal_12473 ;
    wire new_AGEMA_signal_12474 ;
    wire new_AGEMA_signal_12475 ;
    wire new_AGEMA_signal_12476 ;
    wire new_AGEMA_signal_12477 ;
    wire new_AGEMA_signal_12478 ;
    wire new_AGEMA_signal_12479 ;
    wire new_AGEMA_signal_12480 ;
    wire new_AGEMA_signal_12481 ;
    wire new_AGEMA_signal_12482 ;
    wire new_AGEMA_signal_12483 ;
    wire new_AGEMA_signal_12484 ;
    wire new_AGEMA_signal_12485 ;
    wire new_AGEMA_signal_12486 ;
    wire new_AGEMA_signal_12487 ;
    wire new_AGEMA_signal_12488 ;
    wire new_AGEMA_signal_12489 ;
    wire new_AGEMA_signal_12490 ;
    wire new_AGEMA_signal_12491 ;
    wire new_AGEMA_signal_12492 ;
    wire new_AGEMA_signal_12493 ;
    wire new_AGEMA_signal_12494 ;
    wire new_AGEMA_signal_12495 ;
    wire new_AGEMA_signal_12496 ;
    wire new_AGEMA_signal_12497 ;
    wire new_AGEMA_signal_12498 ;
    wire new_AGEMA_signal_12499 ;
    wire new_AGEMA_signal_12500 ;
    wire new_AGEMA_signal_12501 ;
    wire new_AGEMA_signal_12502 ;
    wire new_AGEMA_signal_12503 ;
    wire new_AGEMA_signal_12504 ;
    wire new_AGEMA_signal_12505 ;
    wire new_AGEMA_signal_12506 ;
    wire new_AGEMA_signal_12507 ;
    wire new_AGEMA_signal_12508 ;
    wire new_AGEMA_signal_12509 ;
    wire new_AGEMA_signal_12510 ;
    wire new_AGEMA_signal_12511 ;
    wire new_AGEMA_signal_12512 ;
    wire new_AGEMA_signal_12513 ;
    wire new_AGEMA_signal_12514 ;
    wire new_AGEMA_signal_12515 ;
    wire new_AGEMA_signal_12516 ;
    wire new_AGEMA_signal_12517 ;
    wire new_AGEMA_signal_12518 ;
    wire new_AGEMA_signal_12519 ;
    wire new_AGEMA_signal_12520 ;
    wire new_AGEMA_signal_12521 ;
    wire new_AGEMA_signal_12522 ;
    wire new_AGEMA_signal_12523 ;
    wire new_AGEMA_signal_12524 ;
    wire new_AGEMA_signal_12525 ;
    wire new_AGEMA_signal_12526 ;
    wire new_AGEMA_signal_12527 ;
    wire new_AGEMA_signal_12528 ;
    wire new_AGEMA_signal_12529 ;
    wire new_AGEMA_signal_12530 ;
    wire new_AGEMA_signal_12531 ;
    wire new_AGEMA_signal_12532 ;
    wire new_AGEMA_signal_12533 ;
    wire new_AGEMA_signal_12534 ;
    wire new_AGEMA_signal_12535 ;
    wire new_AGEMA_signal_12536 ;
    wire new_AGEMA_signal_12537 ;
    wire new_AGEMA_signal_12538 ;
    wire new_AGEMA_signal_12539 ;
    wire new_AGEMA_signal_12540 ;
    wire new_AGEMA_signal_12541 ;
    wire new_AGEMA_signal_12542 ;
    wire new_AGEMA_signal_12543 ;
    wire new_AGEMA_signal_12544 ;
    wire new_AGEMA_signal_12545 ;
    wire new_AGEMA_signal_12546 ;
    wire new_AGEMA_signal_12547 ;
    wire new_AGEMA_signal_12548 ;
    wire new_AGEMA_signal_12549 ;
    wire new_AGEMA_signal_12550 ;
    wire new_AGEMA_signal_12551 ;
    wire new_AGEMA_signal_12552 ;
    wire new_AGEMA_signal_12553 ;
    wire new_AGEMA_signal_12554 ;
    wire new_AGEMA_signal_12555 ;
    wire new_AGEMA_signal_12556 ;
    wire new_AGEMA_signal_12557 ;
    wire new_AGEMA_signal_12558 ;
    wire new_AGEMA_signal_12559 ;
    wire new_AGEMA_signal_12560 ;
    wire new_AGEMA_signal_12561 ;
    wire new_AGEMA_signal_12562 ;
    wire new_AGEMA_signal_12563 ;
    wire new_AGEMA_signal_12564 ;
    wire new_AGEMA_signal_12565 ;
    wire new_AGEMA_signal_12566 ;
    wire new_AGEMA_signal_12567 ;
    wire new_AGEMA_signal_12568 ;
    wire new_AGEMA_signal_12569 ;
    wire new_AGEMA_signal_12570 ;
    wire new_AGEMA_signal_12571 ;
    wire new_AGEMA_signal_12572 ;
    wire new_AGEMA_signal_12573 ;
    wire new_AGEMA_signal_12574 ;
    wire new_AGEMA_signal_12575 ;
    wire new_AGEMA_signal_12576 ;
    wire new_AGEMA_signal_12577 ;
    wire new_AGEMA_signal_12578 ;
    wire new_AGEMA_signal_12579 ;
    wire new_AGEMA_signal_12580 ;
    wire new_AGEMA_signal_12581 ;
    wire new_AGEMA_signal_12582 ;
    wire new_AGEMA_signal_12583 ;
    wire new_AGEMA_signal_12584 ;
    wire new_AGEMA_signal_12585 ;
    wire new_AGEMA_signal_12586 ;
    wire new_AGEMA_signal_12587 ;
    wire new_AGEMA_signal_12588 ;
    wire new_AGEMA_signal_12589 ;
    wire new_AGEMA_signal_12590 ;
    wire new_AGEMA_signal_12591 ;
    wire new_AGEMA_signal_12592 ;
    wire new_AGEMA_signal_12593 ;
    wire new_AGEMA_signal_12594 ;
    wire new_AGEMA_signal_12595 ;
    wire new_AGEMA_signal_12596 ;
    wire new_AGEMA_signal_12597 ;
    wire new_AGEMA_signal_12598 ;
    wire new_AGEMA_signal_12599 ;
    wire new_AGEMA_signal_12600 ;
    wire new_AGEMA_signal_12601 ;
    wire new_AGEMA_signal_12602 ;
    wire new_AGEMA_signal_12603 ;
    wire new_AGEMA_signal_12604 ;
    wire new_AGEMA_signal_12605 ;
    wire new_AGEMA_signal_12606 ;
    wire new_AGEMA_signal_12607 ;
    wire new_AGEMA_signal_12608 ;
    wire new_AGEMA_signal_12609 ;
    wire new_AGEMA_signal_12610 ;
    wire new_AGEMA_signal_12611 ;
    wire new_AGEMA_signal_12612 ;
    wire new_AGEMA_signal_12613 ;
    wire new_AGEMA_signal_12614 ;
    wire new_AGEMA_signal_12615 ;
    wire new_AGEMA_signal_12616 ;
    wire new_AGEMA_signal_12617 ;
    wire new_AGEMA_signal_12618 ;
    wire new_AGEMA_signal_12619 ;
    wire new_AGEMA_signal_12620 ;
    wire new_AGEMA_signal_12621 ;
    wire new_AGEMA_signal_12622 ;
    wire new_AGEMA_signal_12623 ;
    wire new_AGEMA_signal_12624 ;
    wire new_AGEMA_signal_12625 ;
    wire new_AGEMA_signal_12626 ;
    wire new_AGEMA_signal_12627 ;
    wire new_AGEMA_signal_12628 ;
    wire new_AGEMA_signal_12629 ;
    wire new_AGEMA_signal_12630 ;
    wire new_AGEMA_signal_12631 ;
    wire new_AGEMA_signal_12632 ;
    wire new_AGEMA_signal_12633 ;
    wire new_AGEMA_signal_12634 ;
    wire new_AGEMA_signal_12635 ;
    wire new_AGEMA_signal_12636 ;
    wire new_AGEMA_signal_12637 ;
    wire new_AGEMA_signal_12638 ;
    wire new_AGEMA_signal_12639 ;
    wire new_AGEMA_signal_12640 ;
    wire new_AGEMA_signal_12641 ;
    wire new_AGEMA_signal_12642 ;
    wire new_AGEMA_signal_12643 ;
    wire new_AGEMA_signal_12644 ;
    wire new_AGEMA_signal_12645 ;
    wire new_AGEMA_signal_12646 ;
    wire new_AGEMA_signal_12647 ;
    wire new_AGEMA_signal_12648 ;
    wire new_AGEMA_signal_12649 ;
    wire new_AGEMA_signal_12650 ;
    wire new_AGEMA_signal_12651 ;
    wire new_AGEMA_signal_12652 ;
    wire new_AGEMA_signal_12653 ;
    wire new_AGEMA_signal_12654 ;
    wire new_AGEMA_signal_12655 ;
    wire new_AGEMA_signal_12656 ;
    wire new_AGEMA_signal_12657 ;
    wire new_AGEMA_signal_12658 ;
    wire new_AGEMA_signal_12659 ;
    wire new_AGEMA_signal_12660 ;
    wire new_AGEMA_signal_12661 ;
    wire new_AGEMA_signal_12662 ;
    wire new_AGEMA_signal_12663 ;
    wire new_AGEMA_signal_12664 ;
    wire new_AGEMA_signal_12665 ;
    wire new_AGEMA_signal_12666 ;
    wire new_AGEMA_signal_12667 ;
    wire new_AGEMA_signal_12668 ;
    wire new_AGEMA_signal_12669 ;
    wire new_AGEMA_signal_12670 ;
    wire new_AGEMA_signal_12671 ;
    wire new_AGEMA_signal_12672 ;
    wire new_AGEMA_signal_12673 ;
    wire new_AGEMA_signal_12674 ;
    wire new_AGEMA_signal_12675 ;
    wire new_AGEMA_signal_12676 ;
    wire new_AGEMA_signal_12677 ;
    wire new_AGEMA_signal_12678 ;
    wire new_AGEMA_signal_12679 ;
    wire new_AGEMA_signal_12680 ;
    wire new_AGEMA_signal_12681 ;
    wire new_AGEMA_signal_12682 ;
    wire new_AGEMA_signal_12683 ;
    wire new_AGEMA_signal_12684 ;
    wire new_AGEMA_signal_12685 ;
    wire new_AGEMA_signal_12686 ;
    wire new_AGEMA_signal_12687 ;
    wire new_AGEMA_signal_12688 ;
    wire new_AGEMA_signal_12689 ;
    wire new_AGEMA_signal_12690 ;
    wire new_AGEMA_signal_12691 ;
    wire new_AGEMA_signal_12692 ;
    wire new_AGEMA_signal_12693 ;
    wire new_AGEMA_signal_12694 ;
    wire new_AGEMA_signal_12695 ;
    wire new_AGEMA_signal_12696 ;
    wire new_AGEMA_signal_12697 ;
    wire new_AGEMA_signal_12698 ;
    wire new_AGEMA_signal_12699 ;
    wire new_AGEMA_signal_12700 ;
    wire new_AGEMA_signal_12701 ;
    wire new_AGEMA_signal_12702 ;
    wire new_AGEMA_signal_12703 ;
    wire new_AGEMA_signal_12704 ;
    wire new_AGEMA_signal_12705 ;
    wire new_AGEMA_signal_12706 ;
    wire new_AGEMA_signal_12707 ;
    wire new_AGEMA_signal_12708 ;
    wire new_AGEMA_signal_12709 ;
    wire new_AGEMA_signal_12710 ;
    wire new_AGEMA_signal_12711 ;
    wire new_AGEMA_signal_12712 ;
    wire new_AGEMA_signal_12713 ;
    wire new_AGEMA_signal_12714 ;
    wire new_AGEMA_signal_12715 ;
    wire new_AGEMA_signal_12716 ;
    wire new_AGEMA_signal_12717 ;
    wire new_AGEMA_signal_12718 ;
    wire new_AGEMA_signal_12719 ;
    wire new_AGEMA_signal_12720 ;
    wire new_AGEMA_signal_12721 ;
    wire new_AGEMA_signal_12722 ;
    wire new_AGEMA_signal_12723 ;
    wire new_AGEMA_signal_12724 ;
    wire new_AGEMA_signal_12725 ;
    wire new_AGEMA_signal_12726 ;
    wire new_AGEMA_signal_12727 ;
    wire new_AGEMA_signal_12728 ;
    wire new_AGEMA_signal_12729 ;
    wire new_AGEMA_signal_12730 ;
    wire new_AGEMA_signal_12731 ;
    wire new_AGEMA_signal_12732 ;
    wire new_AGEMA_signal_12733 ;
    wire new_AGEMA_signal_12734 ;
    wire new_AGEMA_signal_12735 ;
    wire new_AGEMA_signal_12736 ;
    wire new_AGEMA_signal_12737 ;
    wire new_AGEMA_signal_12738 ;
    wire new_AGEMA_signal_12739 ;
    wire new_AGEMA_signal_12740 ;
    wire new_AGEMA_signal_12741 ;
    wire new_AGEMA_signal_12742 ;
    wire new_AGEMA_signal_12743 ;
    wire new_AGEMA_signal_12744 ;
    wire new_AGEMA_signal_12745 ;
    wire new_AGEMA_signal_12746 ;
    wire new_AGEMA_signal_12747 ;
    wire new_AGEMA_signal_12748 ;
    wire new_AGEMA_signal_12749 ;
    wire new_AGEMA_signal_12750 ;
    wire new_AGEMA_signal_12751 ;
    wire new_AGEMA_signal_12752 ;
    wire new_AGEMA_signal_12753 ;
    wire new_AGEMA_signal_12754 ;
    wire new_AGEMA_signal_12755 ;
    wire new_AGEMA_signal_12756 ;
    wire new_AGEMA_signal_12757 ;
    wire new_AGEMA_signal_12758 ;
    wire new_AGEMA_signal_12759 ;
    wire new_AGEMA_signal_12760 ;
    wire new_AGEMA_signal_12761 ;
    wire new_AGEMA_signal_12762 ;
    wire new_AGEMA_signal_12763 ;
    wire new_AGEMA_signal_12764 ;
    wire new_AGEMA_signal_12765 ;
    wire new_AGEMA_signal_12766 ;
    wire new_AGEMA_signal_12767 ;
    wire new_AGEMA_signal_12768 ;
    wire new_AGEMA_signal_12769 ;
    wire new_AGEMA_signal_12770 ;
    wire new_AGEMA_signal_12771 ;
    wire new_AGEMA_signal_12772 ;
    wire new_AGEMA_signal_12773 ;
    wire new_AGEMA_signal_12774 ;
    wire new_AGEMA_signal_12775 ;
    wire new_AGEMA_signal_12776 ;
    wire new_AGEMA_signal_12777 ;
    wire new_AGEMA_signal_12778 ;
    wire new_AGEMA_signal_12779 ;
    wire new_AGEMA_signal_12780 ;
    wire new_AGEMA_signal_12781 ;
    wire new_AGEMA_signal_12782 ;
    wire new_AGEMA_signal_12783 ;
    wire new_AGEMA_signal_12784 ;
    wire new_AGEMA_signal_12785 ;
    wire new_AGEMA_signal_12786 ;
    wire new_AGEMA_signal_12787 ;
    wire new_AGEMA_signal_12788 ;
    wire new_AGEMA_signal_12789 ;
    wire new_AGEMA_signal_12790 ;
    wire new_AGEMA_signal_12791 ;
    wire new_AGEMA_signal_12792 ;
    wire new_AGEMA_signal_12793 ;
    wire new_AGEMA_signal_12794 ;
    wire new_AGEMA_signal_12795 ;
    wire new_AGEMA_signal_12796 ;
    wire new_AGEMA_signal_12797 ;
    wire new_AGEMA_signal_12798 ;
    wire new_AGEMA_signal_12799 ;
    wire new_AGEMA_signal_12800 ;
    wire new_AGEMA_signal_12801 ;
    wire new_AGEMA_signal_12802 ;
    wire new_AGEMA_signal_12803 ;
    wire new_AGEMA_signal_12804 ;
    wire new_AGEMA_signal_12805 ;
    wire new_AGEMA_signal_12806 ;
    wire new_AGEMA_signal_12807 ;
    wire new_AGEMA_signal_12808 ;
    wire new_AGEMA_signal_12809 ;
    wire new_AGEMA_signal_12810 ;
    wire new_AGEMA_signal_12811 ;
    wire new_AGEMA_signal_12812 ;
    wire new_AGEMA_signal_12813 ;
    wire new_AGEMA_signal_12814 ;
    wire new_AGEMA_signal_12815 ;
    wire new_AGEMA_signal_12816 ;
    wire new_AGEMA_signal_12817 ;
    wire new_AGEMA_signal_12818 ;
    wire new_AGEMA_signal_12819 ;
    wire new_AGEMA_signal_12820 ;
    wire new_AGEMA_signal_12821 ;
    wire new_AGEMA_signal_12822 ;
    wire new_AGEMA_signal_12823 ;
    wire new_AGEMA_signal_12824 ;
    wire new_AGEMA_signal_12825 ;
    wire new_AGEMA_signal_12826 ;
    wire new_AGEMA_signal_12827 ;
    wire new_AGEMA_signal_12828 ;
    wire new_AGEMA_signal_12829 ;
    wire new_AGEMA_signal_12830 ;
    wire new_AGEMA_signal_12831 ;
    wire new_AGEMA_signal_12832 ;
    wire new_AGEMA_signal_12833 ;
    wire new_AGEMA_signal_12834 ;
    wire new_AGEMA_signal_12835 ;
    wire new_AGEMA_signal_12836 ;
    wire new_AGEMA_signal_12837 ;
    wire new_AGEMA_signal_12838 ;
    wire new_AGEMA_signal_12839 ;
    wire new_AGEMA_signal_12840 ;
    wire new_AGEMA_signal_12841 ;
    wire new_AGEMA_signal_12842 ;
    wire new_AGEMA_signal_12843 ;
    wire new_AGEMA_signal_12844 ;
    wire new_AGEMA_signal_12845 ;
    wire new_AGEMA_signal_12846 ;
    wire new_AGEMA_signal_12847 ;
    wire new_AGEMA_signal_12848 ;
    wire new_AGEMA_signal_12849 ;
    wire new_AGEMA_signal_12850 ;
    wire new_AGEMA_signal_12851 ;
    wire new_AGEMA_signal_12852 ;
    wire new_AGEMA_signal_12853 ;
    wire new_AGEMA_signal_12854 ;
    wire new_AGEMA_signal_12855 ;
    wire new_AGEMA_signal_12856 ;
    wire new_AGEMA_signal_12857 ;
    wire new_AGEMA_signal_12858 ;
    wire new_AGEMA_signal_12859 ;
    wire new_AGEMA_signal_12860 ;
    wire new_AGEMA_signal_12861 ;
    wire new_AGEMA_signal_12862 ;
    wire new_AGEMA_signal_12863 ;
    wire new_AGEMA_signal_12864 ;
    wire new_AGEMA_signal_12865 ;
    wire new_AGEMA_signal_12866 ;
    wire new_AGEMA_signal_12867 ;
    wire new_AGEMA_signal_12868 ;
    wire new_AGEMA_signal_12869 ;
    wire new_AGEMA_signal_12870 ;
    wire new_AGEMA_signal_12871 ;
    wire new_AGEMA_signal_12872 ;
    wire new_AGEMA_signal_12873 ;
    wire new_AGEMA_signal_12874 ;
    wire new_AGEMA_signal_12875 ;
    wire new_AGEMA_signal_12876 ;
    wire new_AGEMA_signal_12877 ;
    wire new_AGEMA_signal_12878 ;
    wire new_AGEMA_signal_12879 ;
    wire new_AGEMA_signal_12880 ;
    wire new_AGEMA_signal_12881 ;
    wire new_AGEMA_signal_12882 ;
    wire new_AGEMA_signal_12883 ;
    wire new_AGEMA_signal_12884 ;
    wire new_AGEMA_signal_12885 ;
    wire new_AGEMA_signal_12886 ;
    wire new_AGEMA_signal_12887 ;
    wire new_AGEMA_signal_12888 ;
    wire new_AGEMA_signal_12889 ;
    wire new_AGEMA_signal_12890 ;
    wire new_AGEMA_signal_12891 ;
    wire new_AGEMA_signal_12892 ;
    wire new_AGEMA_signal_12893 ;
    wire new_AGEMA_signal_12894 ;
    wire new_AGEMA_signal_12895 ;
    wire new_AGEMA_signal_12896 ;
    wire new_AGEMA_signal_12897 ;
    wire new_AGEMA_signal_12898 ;
    wire new_AGEMA_signal_12899 ;
    wire new_AGEMA_signal_12900 ;
    wire new_AGEMA_signal_12901 ;
    wire new_AGEMA_signal_12902 ;
    wire new_AGEMA_signal_12903 ;
    wire new_AGEMA_signal_12904 ;
    wire new_AGEMA_signal_12905 ;
    wire new_AGEMA_signal_12906 ;
    wire new_AGEMA_signal_12907 ;
    wire new_AGEMA_signal_12908 ;
    wire new_AGEMA_signal_12909 ;
    wire new_AGEMA_signal_12910 ;
    wire new_AGEMA_signal_12911 ;
    wire new_AGEMA_signal_12912 ;
    wire new_AGEMA_signal_12913 ;
    wire new_AGEMA_signal_12914 ;
    wire new_AGEMA_signal_12915 ;
    wire new_AGEMA_signal_12916 ;
    wire new_AGEMA_signal_12917 ;
    wire new_AGEMA_signal_12918 ;
    wire new_AGEMA_signal_12919 ;
    wire new_AGEMA_signal_12920 ;
    wire new_AGEMA_signal_12921 ;
    wire new_AGEMA_signal_12922 ;
    wire new_AGEMA_signal_12923 ;
    wire new_AGEMA_signal_12924 ;
    wire new_AGEMA_signal_12925 ;
    wire new_AGEMA_signal_12926 ;
    wire new_AGEMA_signal_12927 ;
    wire new_AGEMA_signal_12928 ;
    wire new_AGEMA_signal_12929 ;
    wire new_AGEMA_signal_12930 ;
    wire new_AGEMA_signal_12931 ;
    wire new_AGEMA_signal_12932 ;
    wire new_AGEMA_signal_12933 ;
    wire new_AGEMA_signal_12934 ;
    wire new_AGEMA_signal_12935 ;
    wire new_AGEMA_signal_12936 ;
    wire new_AGEMA_signal_12937 ;
    wire new_AGEMA_signal_12938 ;
    wire new_AGEMA_signal_12939 ;
    wire new_AGEMA_signal_12940 ;
    wire new_AGEMA_signal_12941 ;
    wire new_AGEMA_signal_12942 ;
    wire new_AGEMA_signal_12943 ;
    wire new_AGEMA_signal_12944 ;
    wire new_AGEMA_signal_12945 ;
    wire new_AGEMA_signal_12946 ;
    wire new_AGEMA_signal_12947 ;
    wire new_AGEMA_signal_12948 ;
    wire new_AGEMA_signal_12949 ;
    wire new_AGEMA_signal_12950 ;
    wire new_AGEMA_signal_12951 ;
    wire new_AGEMA_signal_12952 ;
    wire new_AGEMA_signal_12953 ;
    wire new_AGEMA_signal_12954 ;
    wire new_AGEMA_signal_12955 ;
    wire new_AGEMA_signal_12956 ;
    wire new_AGEMA_signal_12957 ;
    wire new_AGEMA_signal_12958 ;
    wire new_AGEMA_signal_12959 ;
    wire new_AGEMA_signal_12960 ;
    wire new_AGEMA_signal_12961 ;
    wire new_AGEMA_signal_12962 ;
    wire new_AGEMA_signal_12963 ;
    wire new_AGEMA_signal_12964 ;
    wire new_AGEMA_signal_12965 ;
    wire new_AGEMA_signal_12966 ;
    wire new_AGEMA_signal_12967 ;
    wire new_AGEMA_signal_12968 ;
    wire new_AGEMA_signal_12969 ;
    wire new_AGEMA_signal_12970 ;
    wire new_AGEMA_signal_12971 ;
    wire new_AGEMA_signal_12972 ;
    wire new_AGEMA_signal_12973 ;
    wire new_AGEMA_signal_12974 ;
    wire new_AGEMA_signal_12975 ;
    wire new_AGEMA_signal_12976 ;
    wire new_AGEMA_signal_12977 ;
    wire new_AGEMA_signal_12978 ;
    wire new_AGEMA_signal_12979 ;
    wire new_AGEMA_signal_12980 ;
    wire new_AGEMA_signal_12981 ;
    wire new_AGEMA_signal_12982 ;
    wire new_AGEMA_signal_12983 ;
    wire new_AGEMA_signal_12984 ;
    wire new_AGEMA_signal_12985 ;
    wire new_AGEMA_signal_12986 ;
    wire new_AGEMA_signal_12987 ;
    wire new_AGEMA_signal_12988 ;
    wire new_AGEMA_signal_12989 ;
    wire new_AGEMA_signal_12990 ;
    wire new_AGEMA_signal_12991 ;
    wire new_AGEMA_signal_12992 ;
    wire new_AGEMA_signal_12993 ;
    wire new_AGEMA_signal_12994 ;
    wire new_AGEMA_signal_12995 ;
    wire new_AGEMA_signal_12996 ;
    wire new_AGEMA_signal_12997 ;
    wire new_AGEMA_signal_12998 ;
    wire new_AGEMA_signal_12999 ;
    wire new_AGEMA_signal_13000 ;
    wire new_AGEMA_signal_13001 ;
    wire new_AGEMA_signal_13002 ;
    wire new_AGEMA_signal_13003 ;
    wire new_AGEMA_signal_13004 ;
    wire new_AGEMA_signal_13005 ;
    wire new_AGEMA_signal_13006 ;
    wire new_AGEMA_signal_13007 ;
    wire new_AGEMA_signal_13008 ;
    wire new_AGEMA_signal_13009 ;
    wire new_AGEMA_signal_13010 ;
    wire new_AGEMA_signal_13011 ;
    wire new_AGEMA_signal_13012 ;
    wire new_AGEMA_signal_13013 ;
    wire new_AGEMA_signal_13014 ;
    wire new_AGEMA_signal_13015 ;
    wire new_AGEMA_signal_13016 ;
    wire new_AGEMA_signal_13017 ;
    wire new_AGEMA_signal_13018 ;
    wire new_AGEMA_signal_13019 ;
    wire new_AGEMA_signal_13020 ;
    wire new_AGEMA_signal_13021 ;
    wire new_AGEMA_signal_13022 ;
    wire new_AGEMA_signal_13023 ;
    wire new_AGEMA_signal_13024 ;
    wire new_AGEMA_signal_13025 ;
    wire new_AGEMA_signal_13026 ;
    wire new_AGEMA_signal_13027 ;
    wire new_AGEMA_signal_13028 ;
    wire new_AGEMA_signal_13029 ;
    wire new_AGEMA_signal_13030 ;
    wire new_AGEMA_signal_13031 ;
    wire new_AGEMA_signal_13032 ;
    wire new_AGEMA_signal_13033 ;
    wire new_AGEMA_signal_13034 ;
    wire new_AGEMA_signal_13035 ;
    wire new_AGEMA_signal_13036 ;
    wire new_AGEMA_signal_13037 ;
    wire new_AGEMA_signal_13038 ;
    wire new_AGEMA_signal_13039 ;
    wire new_AGEMA_signal_13040 ;
    wire new_AGEMA_signal_13041 ;
    wire new_AGEMA_signal_13042 ;
    wire new_AGEMA_signal_13043 ;
    wire new_AGEMA_signal_13044 ;
    wire new_AGEMA_signal_13045 ;
    wire new_AGEMA_signal_13046 ;
    wire new_AGEMA_signal_13047 ;
    wire new_AGEMA_signal_13048 ;
    wire new_AGEMA_signal_13049 ;
    wire new_AGEMA_signal_13050 ;
    wire new_AGEMA_signal_13051 ;
    wire new_AGEMA_signal_13052 ;
    wire new_AGEMA_signal_13053 ;
    wire new_AGEMA_signal_13054 ;
    wire new_AGEMA_signal_13055 ;
    wire new_AGEMA_signal_13056 ;
    wire new_AGEMA_signal_13057 ;
    wire new_AGEMA_signal_13058 ;
    wire new_AGEMA_signal_13059 ;
    wire new_AGEMA_signal_13060 ;
    wire new_AGEMA_signal_13061 ;
    wire new_AGEMA_signal_13062 ;
    wire new_AGEMA_signal_13063 ;
    wire new_AGEMA_signal_13064 ;
    wire new_AGEMA_signal_13065 ;
    wire new_AGEMA_signal_13066 ;
    wire new_AGEMA_signal_13067 ;
    wire new_AGEMA_signal_13068 ;
    wire new_AGEMA_signal_13069 ;
    wire new_AGEMA_signal_13070 ;
    wire new_AGEMA_signal_13071 ;
    wire new_AGEMA_signal_13072 ;
    wire new_AGEMA_signal_13073 ;
    wire new_AGEMA_signal_13074 ;
    wire new_AGEMA_signal_13075 ;
    wire new_AGEMA_signal_13076 ;
    wire new_AGEMA_signal_13077 ;
    wire new_AGEMA_signal_13078 ;
    wire new_AGEMA_signal_13079 ;
    wire new_AGEMA_signal_13080 ;
    wire new_AGEMA_signal_13081 ;
    wire new_AGEMA_signal_13082 ;
    wire new_AGEMA_signal_13083 ;
    wire new_AGEMA_signal_13084 ;
    wire new_AGEMA_signal_13085 ;
    wire new_AGEMA_signal_13086 ;
    wire new_AGEMA_signal_13087 ;
    wire new_AGEMA_signal_13088 ;
    wire new_AGEMA_signal_13089 ;
    wire new_AGEMA_signal_13090 ;
    wire new_AGEMA_signal_13091 ;
    wire new_AGEMA_signal_13092 ;
    wire new_AGEMA_signal_13093 ;
    wire new_AGEMA_signal_13094 ;
    wire new_AGEMA_signal_13095 ;
    wire new_AGEMA_signal_13096 ;
    wire new_AGEMA_signal_13097 ;
    wire new_AGEMA_signal_13098 ;
    wire new_AGEMA_signal_13099 ;
    wire new_AGEMA_signal_13100 ;
    wire new_AGEMA_signal_13101 ;
    wire new_AGEMA_signal_13102 ;
    wire new_AGEMA_signal_13103 ;
    wire new_AGEMA_signal_13104 ;
    wire new_AGEMA_signal_13105 ;
    wire new_AGEMA_signal_13106 ;
    wire new_AGEMA_signal_13107 ;
    wire new_AGEMA_signal_13108 ;
    wire new_AGEMA_signal_13109 ;
    wire new_AGEMA_signal_13110 ;
    wire new_AGEMA_signal_13111 ;
    wire new_AGEMA_signal_13112 ;
    wire new_AGEMA_signal_13113 ;
    wire new_AGEMA_signal_13114 ;
    wire new_AGEMA_signal_13115 ;
    wire new_AGEMA_signal_13116 ;
    wire new_AGEMA_signal_13117 ;
    wire new_AGEMA_signal_13118 ;
    wire new_AGEMA_signal_13119 ;
    wire new_AGEMA_signal_13120 ;
    wire new_AGEMA_signal_13121 ;
    wire new_AGEMA_signal_13122 ;
    wire new_AGEMA_signal_13123 ;
    wire new_AGEMA_signal_13124 ;
    wire new_AGEMA_signal_13125 ;
    wire new_AGEMA_signal_13126 ;
    wire new_AGEMA_signal_13127 ;
    wire new_AGEMA_signal_13128 ;
    wire new_AGEMA_signal_13129 ;
    wire new_AGEMA_signal_13130 ;
    wire new_AGEMA_signal_13131 ;
    wire new_AGEMA_signal_13132 ;
    wire new_AGEMA_signal_13133 ;
    wire new_AGEMA_signal_13134 ;
    wire new_AGEMA_signal_13135 ;
    wire new_AGEMA_signal_13136 ;
    wire new_AGEMA_signal_13137 ;
    wire new_AGEMA_signal_13138 ;
    wire new_AGEMA_signal_13139 ;
    wire new_AGEMA_signal_13140 ;
    wire new_AGEMA_signal_13141 ;
    wire new_AGEMA_signal_13142 ;
    wire new_AGEMA_signal_13143 ;
    wire new_AGEMA_signal_13144 ;
    wire new_AGEMA_signal_13145 ;
    wire new_AGEMA_signal_13146 ;
    wire new_AGEMA_signal_13147 ;
    wire new_AGEMA_signal_13148 ;
    wire new_AGEMA_signal_13149 ;
    wire new_AGEMA_signal_13150 ;
    wire new_AGEMA_signal_13151 ;
    wire new_AGEMA_signal_13152 ;
    wire new_AGEMA_signal_13153 ;
    wire new_AGEMA_signal_13154 ;
    wire new_AGEMA_signal_13155 ;
    wire new_AGEMA_signal_13156 ;
    wire new_AGEMA_signal_13157 ;
    wire new_AGEMA_signal_13158 ;
    wire new_AGEMA_signal_13159 ;
    wire new_AGEMA_signal_13160 ;
    wire new_AGEMA_signal_13161 ;
    wire new_AGEMA_signal_13162 ;
    wire new_AGEMA_signal_13163 ;
    wire new_AGEMA_signal_13164 ;
    wire new_AGEMA_signal_13165 ;
    wire new_AGEMA_signal_13166 ;
    wire new_AGEMA_signal_13167 ;
    wire new_AGEMA_signal_13168 ;
    wire new_AGEMA_signal_13169 ;
    wire new_AGEMA_signal_13170 ;
    wire new_AGEMA_signal_13171 ;
    wire new_AGEMA_signal_13172 ;
    wire new_AGEMA_signal_13173 ;
    wire new_AGEMA_signal_13174 ;
    wire new_AGEMA_signal_13175 ;
    wire new_AGEMA_signal_13176 ;
    wire new_AGEMA_signal_13177 ;
    wire new_AGEMA_signal_13178 ;
    wire new_AGEMA_signal_13179 ;
    wire new_AGEMA_signal_13180 ;
    wire new_AGEMA_signal_13181 ;
    wire new_AGEMA_signal_13182 ;
    wire new_AGEMA_signal_13183 ;
    wire new_AGEMA_signal_13184 ;
    wire new_AGEMA_signal_13185 ;
    wire new_AGEMA_signal_13186 ;
    wire new_AGEMA_signal_13187 ;
    wire new_AGEMA_signal_13188 ;
    wire new_AGEMA_signal_13189 ;
    wire new_AGEMA_signal_13190 ;
    wire new_AGEMA_signal_13191 ;
    wire new_AGEMA_signal_13192 ;
    wire new_AGEMA_signal_13193 ;
    wire new_AGEMA_signal_13194 ;
    wire new_AGEMA_signal_13195 ;
    wire new_AGEMA_signal_13196 ;
    wire new_AGEMA_signal_13197 ;
    wire new_AGEMA_signal_13198 ;
    wire new_AGEMA_signal_13199 ;
    wire new_AGEMA_signal_13200 ;
    wire new_AGEMA_signal_13201 ;
    wire new_AGEMA_signal_13202 ;
    wire new_AGEMA_signal_13203 ;
    wire new_AGEMA_signal_13204 ;
    wire new_AGEMA_signal_13205 ;
    wire new_AGEMA_signal_13206 ;
    wire new_AGEMA_signal_13207 ;
    wire new_AGEMA_signal_13208 ;
    wire new_AGEMA_signal_13209 ;
    wire new_AGEMA_signal_13210 ;
    wire new_AGEMA_signal_13211 ;
    wire new_AGEMA_signal_13212 ;
    wire new_AGEMA_signal_13213 ;
    wire new_AGEMA_signal_13214 ;
    wire new_AGEMA_signal_13215 ;
    wire new_AGEMA_signal_13216 ;
    wire new_AGEMA_signal_13217 ;
    wire new_AGEMA_signal_13218 ;
    wire new_AGEMA_signal_13219 ;
    wire new_AGEMA_signal_13220 ;
    wire new_AGEMA_signal_13221 ;
    wire new_AGEMA_signal_13222 ;
    wire new_AGEMA_signal_13223 ;
    wire new_AGEMA_signal_13224 ;
    wire new_AGEMA_signal_13225 ;
    wire new_AGEMA_signal_13226 ;
    wire new_AGEMA_signal_13227 ;
    wire new_AGEMA_signal_13228 ;
    wire new_AGEMA_signal_13229 ;
    wire new_AGEMA_signal_13230 ;
    wire new_AGEMA_signal_13231 ;
    wire new_AGEMA_signal_13232 ;
    wire new_AGEMA_signal_13233 ;
    wire new_AGEMA_signal_13234 ;
    wire new_AGEMA_signal_13235 ;
    wire new_AGEMA_signal_13236 ;
    wire new_AGEMA_signal_13237 ;
    wire new_AGEMA_signal_13238 ;
    wire new_AGEMA_signal_13239 ;
    wire new_AGEMA_signal_13240 ;
    wire new_AGEMA_signal_13241 ;
    wire new_AGEMA_signal_13242 ;
    wire new_AGEMA_signal_13243 ;
    wire new_AGEMA_signal_13244 ;
    wire new_AGEMA_signal_13245 ;
    wire new_AGEMA_signal_13246 ;
    wire new_AGEMA_signal_13247 ;
    wire new_AGEMA_signal_13248 ;
    wire new_AGEMA_signal_13249 ;
    wire new_AGEMA_signal_13250 ;
    wire new_AGEMA_signal_13251 ;
    wire new_AGEMA_signal_13252 ;
    wire new_AGEMA_signal_13253 ;
    wire new_AGEMA_signal_13254 ;
    wire new_AGEMA_signal_13255 ;
    wire new_AGEMA_signal_13256 ;
    wire new_AGEMA_signal_13257 ;
    wire new_AGEMA_signal_13258 ;
    wire new_AGEMA_signal_13259 ;
    wire new_AGEMA_signal_13260 ;
    wire new_AGEMA_signal_13261 ;
    wire new_AGEMA_signal_13262 ;
    wire new_AGEMA_signal_13263 ;
    wire new_AGEMA_signal_13264 ;
    wire new_AGEMA_signal_13265 ;
    wire new_AGEMA_signal_13266 ;
    wire new_AGEMA_signal_13267 ;
    wire new_AGEMA_signal_13268 ;
    wire new_AGEMA_signal_13269 ;
    wire new_AGEMA_signal_13270 ;
    wire new_AGEMA_signal_13271 ;
    wire new_AGEMA_signal_13272 ;
    wire new_AGEMA_signal_13273 ;
    wire new_AGEMA_signal_13274 ;
    wire new_AGEMA_signal_13275 ;
    wire new_AGEMA_signal_13276 ;
    wire new_AGEMA_signal_13277 ;
    wire new_AGEMA_signal_13278 ;
    wire new_AGEMA_signal_13279 ;
    wire new_AGEMA_signal_13280 ;
    wire new_AGEMA_signal_13281 ;
    wire new_AGEMA_signal_13282 ;
    wire new_AGEMA_signal_13283 ;
    wire new_AGEMA_signal_13284 ;
    wire new_AGEMA_signal_13285 ;
    wire new_AGEMA_signal_13286 ;
    wire new_AGEMA_signal_13287 ;
    wire new_AGEMA_signal_13288 ;
    wire new_AGEMA_signal_13289 ;
    wire new_AGEMA_signal_13290 ;
    wire new_AGEMA_signal_13291 ;
    wire new_AGEMA_signal_13292 ;
    wire new_AGEMA_signal_13293 ;
    wire new_AGEMA_signal_13294 ;
    wire new_AGEMA_signal_13295 ;
    wire new_AGEMA_signal_13296 ;
    wire new_AGEMA_signal_13297 ;
    wire new_AGEMA_signal_13298 ;
    wire new_AGEMA_signal_13299 ;
    wire new_AGEMA_signal_13300 ;
    wire new_AGEMA_signal_13301 ;
    wire new_AGEMA_signal_13302 ;
    wire new_AGEMA_signal_13303 ;
    wire new_AGEMA_signal_13304 ;
    wire new_AGEMA_signal_13305 ;
    wire new_AGEMA_signal_13306 ;
    wire new_AGEMA_signal_13307 ;
    wire new_AGEMA_signal_13308 ;
    wire new_AGEMA_signal_13309 ;
    wire new_AGEMA_signal_13310 ;
    wire new_AGEMA_signal_13311 ;
    wire new_AGEMA_signal_13312 ;
    wire new_AGEMA_signal_13313 ;
    wire new_AGEMA_signal_13314 ;
    wire new_AGEMA_signal_13315 ;
    wire new_AGEMA_signal_13316 ;
    wire new_AGEMA_signal_13317 ;
    wire new_AGEMA_signal_13318 ;
    wire new_AGEMA_signal_13319 ;
    wire new_AGEMA_signal_13320 ;
    wire new_AGEMA_signal_13321 ;
    wire new_AGEMA_signal_13322 ;
    wire new_AGEMA_signal_13323 ;
    wire new_AGEMA_signal_13324 ;
    wire new_AGEMA_signal_13325 ;
    wire new_AGEMA_signal_13326 ;
    wire new_AGEMA_signal_13327 ;
    wire new_AGEMA_signal_13328 ;
    wire new_AGEMA_signal_13329 ;
    wire new_AGEMA_signal_13330 ;
    wire new_AGEMA_signal_13331 ;
    wire new_AGEMA_signal_13332 ;
    wire new_AGEMA_signal_13333 ;
    wire new_AGEMA_signal_13334 ;
    wire new_AGEMA_signal_13335 ;
    wire new_AGEMA_signal_13336 ;
    wire new_AGEMA_signal_13337 ;
    wire new_AGEMA_signal_13338 ;
    wire new_AGEMA_signal_13339 ;
    wire new_AGEMA_signal_13340 ;
    wire new_AGEMA_signal_13341 ;
    wire new_AGEMA_signal_13342 ;
    wire new_AGEMA_signal_13343 ;
    wire new_AGEMA_signal_13344 ;
    wire new_AGEMA_signal_13345 ;
    wire new_AGEMA_signal_13346 ;
    wire new_AGEMA_signal_13347 ;
    wire new_AGEMA_signal_13348 ;
    wire new_AGEMA_signal_13349 ;
    wire new_AGEMA_signal_13350 ;
    wire new_AGEMA_signal_13351 ;
    wire new_AGEMA_signal_13352 ;
    wire new_AGEMA_signal_13353 ;
    wire new_AGEMA_signal_13354 ;
    wire new_AGEMA_signal_13355 ;
    wire new_AGEMA_signal_13356 ;
    wire new_AGEMA_signal_13357 ;
    wire new_AGEMA_signal_13358 ;
    wire new_AGEMA_signal_13359 ;
    wire new_AGEMA_signal_13360 ;
    wire new_AGEMA_signal_13361 ;
    wire new_AGEMA_signal_13362 ;
    wire new_AGEMA_signal_13363 ;
    wire new_AGEMA_signal_13364 ;
    wire new_AGEMA_signal_13365 ;
    wire new_AGEMA_signal_13366 ;
    wire new_AGEMA_signal_13367 ;
    wire new_AGEMA_signal_13368 ;
    wire new_AGEMA_signal_13369 ;
    wire new_AGEMA_signal_13370 ;
    wire new_AGEMA_signal_13371 ;
    wire new_AGEMA_signal_13372 ;
    wire new_AGEMA_signal_13373 ;
    wire new_AGEMA_signal_13374 ;
    wire new_AGEMA_signal_13375 ;
    wire new_AGEMA_signal_13376 ;
    wire new_AGEMA_signal_13377 ;
    wire new_AGEMA_signal_13378 ;
    wire new_AGEMA_signal_13379 ;
    wire new_AGEMA_signal_13380 ;
    wire new_AGEMA_signal_13381 ;
    wire new_AGEMA_signal_13382 ;
    wire new_AGEMA_signal_13383 ;
    wire new_AGEMA_signal_13384 ;
    wire new_AGEMA_signal_13385 ;
    wire new_AGEMA_signal_13386 ;
    wire new_AGEMA_signal_13387 ;
    wire new_AGEMA_signal_13388 ;
    wire new_AGEMA_signal_13389 ;
    wire new_AGEMA_signal_13390 ;
    wire new_AGEMA_signal_13391 ;
    wire new_AGEMA_signal_13392 ;
    wire new_AGEMA_signal_13396 ;
    wire new_AGEMA_signal_13397 ;
    wire new_AGEMA_signal_13398 ;
    wire new_AGEMA_signal_13402 ;
    wire new_AGEMA_signal_13403 ;
    wire new_AGEMA_signal_13404 ;
    wire new_AGEMA_signal_13408 ;
    wire new_AGEMA_signal_13409 ;
    wire new_AGEMA_signal_13410 ;
    wire new_AGEMA_signal_13411 ;
    wire new_AGEMA_signal_13412 ;
    wire new_AGEMA_signal_13413 ;
    wire new_AGEMA_signal_13414 ;
    wire new_AGEMA_signal_13415 ;
    wire new_AGEMA_signal_13416 ;
    wire new_AGEMA_signal_13417 ;
    wire new_AGEMA_signal_13418 ;
    wire new_AGEMA_signal_13419 ;
    wire new_AGEMA_signal_13420 ;
    wire new_AGEMA_signal_13421 ;
    wire new_AGEMA_signal_13422 ;
    wire new_AGEMA_signal_13423 ;
    wire new_AGEMA_signal_13424 ;
    wire new_AGEMA_signal_13425 ;
    wire new_AGEMA_signal_13426 ;
    wire new_AGEMA_signal_13427 ;
    wire new_AGEMA_signal_13428 ;
    wire new_AGEMA_signal_13429 ;
    wire new_AGEMA_signal_13430 ;
    wire new_AGEMA_signal_13431 ;
    wire new_AGEMA_signal_13432 ;
    wire new_AGEMA_signal_13433 ;
    wire new_AGEMA_signal_13434 ;
    wire new_AGEMA_signal_13435 ;
    wire new_AGEMA_signal_13436 ;
    wire new_AGEMA_signal_13437 ;
    wire new_AGEMA_signal_13438 ;
    wire new_AGEMA_signal_13439 ;
    wire new_AGEMA_signal_13440 ;
    wire new_AGEMA_signal_13441 ;
    wire new_AGEMA_signal_13442 ;
    wire new_AGEMA_signal_13443 ;
    wire new_AGEMA_signal_13444 ;
    wire new_AGEMA_signal_13445 ;
    wire new_AGEMA_signal_13446 ;
    wire new_AGEMA_signal_13447 ;
    wire new_AGEMA_signal_13448 ;
    wire new_AGEMA_signal_13449 ;
    wire new_AGEMA_signal_13450 ;
    wire new_AGEMA_signal_13451 ;
    wire new_AGEMA_signal_13452 ;
    wire new_AGEMA_signal_13453 ;
    wire new_AGEMA_signal_13454 ;
    wire new_AGEMA_signal_13455 ;
    wire new_AGEMA_signal_13456 ;
    wire new_AGEMA_signal_13457 ;
    wire new_AGEMA_signal_13458 ;
    wire new_AGEMA_signal_13459 ;
    wire new_AGEMA_signal_13460 ;
    wire new_AGEMA_signal_13461 ;
    wire new_AGEMA_signal_13462 ;
    wire new_AGEMA_signal_13463 ;
    wire new_AGEMA_signal_13464 ;
    wire new_AGEMA_signal_13465 ;
    wire new_AGEMA_signal_13466 ;
    wire new_AGEMA_signal_13467 ;
    wire new_AGEMA_signal_13468 ;
    wire new_AGEMA_signal_13469 ;
    wire new_AGEMA_signal_13470 ;
    wire new_AGEMA_signal_13471 ;
    wire new_AGEMA_signal_13472 ;
    wire new_AGEMA_signal_13473 ;
    wire new_AGEMA_signal_13474 ;
    wire new_AGEMA_signal_13475 ;
    wire new_AGEMA_signal_13476 ;
    wire new_AGEMA_signal_13477 ;
    wire new_AGEMA_signal_13478 ;
    wire new_AGEMA_signal_13479 ;
    wire new_AGEMA_signal_13480 ;
    wire new_AGEMA_signal_13481 ;
    wire new_AGEMA_signal_13482 ;
    wire new_AGEMA_signal_13483 ;
    wire new_AGEMA_signal_13484 ;
    wire new_AGEMA_signal_13485 ;
    wire new_AGEMA_signal_13486 ;
    wire new_AGEMA_signal_13487 ;
    wire new_AGEMA_signal_13488 ;
    wire new_AGEMA_signal_13489 ;
    wire new_AGEMA_signal_13490 ;
    wire new_AGEMA_signal_13491 ;
    wire new_AGEMA_signal_13492 ;
    wire new_AGEMA_signal_13493 ;
    wire new_AGEMA_signal_13494 ;
    wire new_AGEMA_signal_13495 ;
    wire new_AGEMA_signal_13496 ;
    wire new_AGEMA_signal_13497 ;
    wire new_AGEMA_signal_13498 ;
    wire new_AGEMA_signal_13499 ;
    wire new_AGEMA_signal_13500 ;
    wire new_AGEMA_signal_13501 ;
    wire new_AGEMA_signal_13502 ;
    wire new_AGEMA_signal_13503 ;
    wire new_AGEMA_signal_13504 ;
    wire new_AGEMA_signal_13505 ;
    wire new_AGEMA_signal_13506 ;
    wire new_AGEMA_signal_13507 ;
    wire new_AGEMA_signal_13508 ;
    wire new_AGEMA_signal_13509 ;
    wire new_AGEMA_signal_13510 ;
    wire new_AGEMA_signal_13511 ;
    wire new_AGEMA_signal_13512 ;
    wire new_AGEMA_signal_13513 ;
    wire new_AGEMA_signal_13514 ;
    wire new_AGEMA_signal_13515 ;
    wire new_AGEMA_signal_13516 ;
    wire new_AGEMA_signal_13517 ;
    wire new_AGEMA_signal_13518 ;
    wire new_AGEMA_signal_13519 ;
    wire new_AGEMA_signal_13520 ;
    wire new_AGEMA_signal_13521 ;
    wire new_AGEMA_signal_13522 ;
    wire new_AGEMA_signal_13523 ;
    wire new_AGEMA_signal_13524 ;
    wire new_AGEMA_signal_13525 ;
    wire new_AGEMA_signal_13526 ;
    wire new_AGEMA_signal_13527 ;
    wire new_AGEMA_signal_13528 ;
    wire new_AGEMA_signal_13529 ;
    wire new_AGEMA_signal_13530 ;
    wire new_AGEMA_signal_13531 ;
    wire new_AGEMA_signal_13532 ;
    wire new_AGEMA_signal_13533 ;
    wire new_AGEMA_signal_13534 ;
    wire new_AGEMA_signal_13535 ;
    wire new_AGEMA_signal_13536 ;
    wire new_AGEMA_signal_13537 ;
    wire new_AGEMA_signal_13538 ;
    wire new_AGEMA_signal_13539 ;
    wire new_AGEMA_signal_13540 ;
    wire new_AGEMA_signal_13541 ;
    wire new_AGEMA_signal_13542 ;
    wire new_AGEMA_signal_13543 ;
    wire new_AGEMA_signal_13544 ;
    wire new_AGEMA_signal_13545 ;
    wire new_AGEMA_signal_13546 ;
    wire new_AGEMA_signal_13547 ;
    wire new_AGEMA_signal_13548 ;
    wire new_AGEMA_signal_13549 ;
    wire new_AGEMA_signal_13550 ;
    wire new_AGEMA_signal_13551 ;
    wire new_AGEMA_signal_13552 ;
    wire new_AGEMA_signal_13553 ;
    wire new_AGEMA_signal_13554 ;
    wire new_AGEMA_signal_13555 ;
    wire new_AGEMA_signal_13556 ;
    wire new_AGEMA_signal_13557 ;
    wire new_AGEMA_signal_13558 ;
    wire new_AGEMA_signal_13559 ;
    wire new_AGEMA_signal_13560 ;
    wire new_AGEMA_signal_13561 ;
    wire new_AGEMA_signal_13562 ;
    wire new_AGEMA_signal_13563 ;
    wire new_AGEMA_signal_13564 ;
    wire new_AGEMA_signal_13565 ;
    wire new_AGEMA_signal_13566 ;
    wire new_AGEMA_signal_13567 ;
    wire new_AGEMA_signal_13568 ;
    wire new_AGEMA_signal_13569 ;
    wire new_AGEMA_signal_13570 ;
    wire new_AGEMA_signal_13571 ;
    wire new_AGEMA_signal_13572 ;
    wire new_AGEMA_signal_13573 ;
    wire new_AGEMA_signal_13574 ;
    wire new_AGEMA_signal_13575 ;
    wire new_AGEMA_signal_13576 ;
    wire new_AGEMA_signal_13577 ;
    wire new_AGEMA_signal_13578 ;
    wire new_AGEMA_signal_13579 ;
    wire new_AGEMA_signal_13580 ;
    wire new_AGEMA_signal_13581 ;
    wire new_AGEMA_signal_13582 ;
    wire new_AGEMA_signal_13583 ;
    wire new_AGEMA_signal_13584 ;
    wire new_AGEMA_signal_13585 ;
    wire new_AGEMA_signal_13586 ;
    wire new_AGEMA_signal_13587 ;
    wire new_AGEMA_signal_13588 ;
    wire new_AGEMA_signal_13589 ;
    wire new_AGEMA_signal_13590 ;
    wire new_AGEMA_signal_13591 ;
    wire new_AGEMA_signal_13592 ;
    wire new_AGEMA_signal_13593 ;
    wire new_AGEMA_signal_13594 ;
    wire new_AGEMA_signal_13595 ;
    wire new_AGEMA_signal_13596 ;
    wire new_AGEMA_signal_13597 ;
    wire new_AGEMA_signal_13598 ;
    wire new_AGEMA_signal_13599 ;
    wire new_AGEMA_signal_13600 ;
    wire new_AGEMA_signal_13601 ;
    wire new_AGEMA_signal_13602 ;
    wire new_AGEMA_signal_13603 ;
    wire new_AGEMA_signal_13604 ;
    wire new_AGEMA_signal_13605 ;
    wire new_AGEMA_signal_13606 ;
    wire new_AGEMA_signal_13607 ;
    wire new_AGEMA_signal_13608 ;
    wire new_AGEMA_signal_13609 ;
    wire new_AGEMA_signal_13610 ;
    wire new_AGEMA_signal_13611 ;
    wire new_AGEMA_signal_13612 ;
    wire new_AGEMA_signal_13613 ;
    wire new_AGEMA_signal_13614 ;
    wire new_AGEMA_signal_13615 ;
    wire new_AGEMA_signal_13616 ;
    wire new_AGEMA_signal_13617 ;
    wire new_AGEMA_signal_13618 ;
    wire new_AGEMA_signal_13619 ;
    wire new_AGEMA_signal_13620 ;
    wire new_AGEMA_signal_13621 ;
    wire new_AGEMA_signal_13622 ;
    wire new_AGEMA_signal_13623 ;
    wire new_AGEMA_signal_13624 ;
    wire new_AGEMA_signal_13625 ;
    wire new_AGEMA_signal_13626 ;
    wire new_AGEMA_signal_13627 ;
    wire new_AGEMA_signal_13628 ;
    wire new_AGEMA_signal_13629 ;
    wire new_AGEMA_signal_13630 ;
    wire new_AGEMA_signal_13631 ;
    wire new_AGEMA_signal_13632 ;
    wire new_AGEMA_signal_13633 ;
    wire new_AGEMA_signal_13634 ;
    wire new_AGEMA_signal_13635 ;
    wire new_AGEMA_signal_13636 ;
    wire new_AGEMA_signal_13637 ;
    wire new_AGEMA_signal_13638 ;
    wire new_AGEMA_signal_13639 ;
    wire new_AGEMA_signal_13640 ;
    wire new_AGEMA_signal_13641 ;
    wire new_AGEMA_signal_13642 ;
    wire new_AGEMA_signal_13643 ;
    wire new_AGEMA_signal_13644 ;
    wire new_AGEMA_signal_13645 ;
    wire new_AGEMA_signal_13646 ;
    wire new_AGEMA_signal_13647 ;
    wire new_AGEMA_signal_13648 ;
    wire new_AGEMA_signal_13649 ;
    wire new_AGEMA_signal_13650 ;
    wire new_AGEMA_signal_13651 ;
    wire new_AGEMA_signal_13652 ;
    wire new_AGEMA_signal_13653 ;
    wire new_AGEMA_signal_13654 ;
    wire new_AGEMA_signal_13655 ;
    wire new_AGEMA_signal_13656 ;
    wire new_AGEMA_signal_13657 ;
    wire new_AGEMA_signal_13658 ;
    wire new_AGEMA_signal_13659 ;
    wire new_AGEMA_signal_13660 ;
    wire new_AGEMA_signal_13661 ;
    wire new_AGEMA_signal_13662 ;
    wire new_AGEMA_signal_13663 ;
    wire new_AGEMA_signal_13664 ;
    wire new_AGEMA_signal_13665 ;
    wire new_AGEMA_signal_13666 ;
    wire new_AGEMA_signal_13667 ;
    wire new_AGEMA_signal_13668 ;
    wire new_AGEMA_signal_13669 ;
    wire new_AGEMA_signal_13670 ;
    wire new_AGEMA_signal_13671 ;
    wire new_AGEMA_signal_13672 ;
    wire new_AGEMA_signal_13673 ;
    wire new_AGEMA_signal_13674 ;
    wire new_AGEMA_signal_13675 ;
    wire new_AGEMA_signal_13676 ;
    wire new_AGEMA_signal_13677 ;
    wire new_AGEMA_signal_13678 ;
    wire new_AGEMA_signal_13679 ;
    wire new_AGEMA_signal_13680 ;
    wire new_AGEMA_signal_13681 ;
    wire new_AGEMA_signal_13682 ;
    wire new_AGEMA_signal_13683 ;
    wire new_AGEMA_signal_13684 ;
    wire new_AGEMA_signal_13685 ;
    wire new_AGEMA_signal_13686 ;
    wire new_AGEMA_signal_13687 ;
    wire new_AGEMA_signal_13688 ;
    wire new_AGEMA_signal_13689 ;
    wire new_AGEMA_signal_13690 ;
    wire new_AGEMA_signal_13691 ;
    wire new_AGEMA_signal_13692 ;
    wire new_AGEMA_signal_13693 ;
    wire new_AGEMA_signal_13694 ;
    wire new_AGEMA_signal_13695 ;
    wire new_AGEMA_signal_13696 ;
    wire new_AGEMA_signal_13697 ;
    wire new_AGEMA_signal_13698 ;
    wire new_AGEMA_signal_13699 ;
    wire new_AGEMA_signal_13700 ;
    wire new_AGEMA_signal_13701 ;
    wire new_AGEMA_signal_13702 ;
    wire new_AGEMA_signal_13703 ;
    wire new_AGEMA_signal_13704 ;
    wire new_AGEMA_signal_13705 ;
    wire new_AGEMA_signal_13706 ;
    wire new_AGEMA_signal_13707 ;
    wire new_AGEMA_signal_13708 ;
    wire new_AGEMA_signal_13709 ;
    wire new_AGEMA_signal_13710 ;
    wire new_AGEMA_signal_13711 ;
    wire new_AGEMA_signal_13712 ;
    wire new_AGEMA_signal_13713 ;
    wire new_AGEMA_signal_13714 ;
    wire new_AGEMA_signal_13715 ;
    wire new_AGEMA_signal_13716 ;
    wire new_AGEMA_signal_13717 ;
    wire new_AGEMA_signal_13718 ;
    wire new_AGEMA_signal_13719 ;
    wire new_AGEMA_signal_13720 ;
    wire new_AGEMA_signal_13721 ;
    wire new_AGEMA_signal_13722 ;
    wire new_AGEMA_signal_13723 ;
    wire new_AGEMA_signal_13724 ;
    wire new_AGEMA_signal_13725 ;
    wire new_AGEMA_signal_13726 ;
    wire new_AGEMA_signal_13727 ;
    wire new_AGEMA_signal_13728 ;
    wire new_AGEMA_signal_13729 ;
    wire new_AGEMA_signal_13730 ;
    wire new_AGEMA_signal_13731 ;
    wire new_AGEMA_signal_13732 ;
    wire new_AGEMA_signal_13733 ;
    wire new_AGEMA_signal_13734 ;
    wire new_AGEMA_signal_13735 ;
    wire new_AGEMA_signal_13736 ;
    wire new_AGEMA_signal_13737 ;
    wire new_AGEMA_signal_13738 ;
    wire new_AGEMA_signal_13739 ;
    wire new_AGEMA_signal_13740 ;
    wire new_AGEMA_signal_13741 ;
    wire new_AGEMA_signal_13742 ;
    wire new_AGEMA_signal_13743 ;
    wire new_AGEMA_signal_13744 ;
    wire new_AGEMA_signal_13745 ;
    wire new_AGEMA_signal_13746 ;
    wire new_AGEMA_signal_13747 ;
    wire new_AGEMA_signal_13748 ;
    wire new_AGEMA_signal_13749 ;
    wire new_AGEMA_signal_13750 ;
    wire new_AGEMA_signal_13751 ;
    wire new_AGEMA_signal_13752 ;
    wire new_AGEMA_signal_13753 ;
    wire new_AGEMA_signal_13754 ;
    wire new_AGEMA_signal_13755 ;
    wire new_AGEMA_signal_13756 ;
    wire new_AGEMA_signal_13757 ;
    wire new_AGEMA_signal_13758 ;
    wire new_AGEMA_signal_13759 ;
    wire new_AGEMA_signal_13760 ;
    wire new_AGEMA_signal_13761 ;
    wire new_AGEMA_signal_13762 ;
    wire new_AGEMA_signal_13763 ;
    wire new_AGEMA_signal_13764 ;
    wire new_AGEMA_signal_13765 ;
    wire new_AGEMA_signal_13766 ;
    wire new_AGEMA_signal_13767 ;
    wire new_AGEMA_signal_13768 ;
    wire new_AGEMA_signal_13769 ;
    wire new_AGEMA_signal_13770 ;
    wire new_AGEMA_signal_13771 ;
    wire new_AGEMA_signal_13772 ;
    wire new_AGEMA_signal_13773 ;
    wire new_AGEMA_signal_13774 ;
    wire new_AGEMA_signal_13775 ;
    wire new_AGEMA_signal_13776 ;
    wire new_AGEMA_signal_13777 ;
    wire new_AGEMA_signal_13778 ;
    wire new_AGEMA_signal_13779 ;
    wire new_AGEMA_signal_13780 ;
    wire new_AGEMA_signal_13781 ;
    wire new_AGEMA_signal_13782 ;
    wire new_AGEMA_signal_13783 ;
    wire new_AGEMA_signal_13784 ;
    wire new_AGEMA_signal_13785 ;
    wire new_AGEMA_signal_13786 ;
    wire new_AGEMA_signal_13787 ;
    wire new_AGEMA_signal_13788 ;
    wire new_AGEMA_signal_13789 ;
    wire new_AGEMA_signal_13790 ;
    wire new_AGEMA_signal_13791 ;
    wire new_AGEMA_signal_13792 ;
    wire new_AGEMA_signal_13793 ;
    wire new_AGEMA_signal_13794 ;
    wire new_AGEMA_signal_13795 ;
    wire new_AGEMA_signal_13796 ;
    wire new_AGEMA_signal_13797 ;
    wire new_AGEMA_signal_13798 ;
    wire new_AGEMA_signal_13799 ;
    wire new_AGEMA_signal_13800 ;
    wire new_AGEMA_signal_13801 ;
    wire new_AGEMA_signal_13802 ;
    wire new_AGEMA_signal_13803 ;
    wire new_AGEMA_signal_13804 ;
    wire new_AGEMA_signal_13805 ;
    wire new_AGEMA_signal_13806 ;
    wire new_AGEMA_signal_13807 ;
    wire new_AGEMA_signal_13808 ;
    wire new_AGEMA_signal_13809 ;
    wire new_AGEMA_signal_13810 ;
    wire new_AGEMA_signal_13811 ;
    wire new_AGEMA_signal_13812 ;
    wire new_AGEMA_signal_13813 ;
    wire new_AGEMA_signal_13814 ;
    wire new_AGEMA_signal_13815 ;
    wire new_AGEMA_signal_13816 ;
    wire new_AGEMA_signal_13817 ;
    wire new_AGEMA_signal_13818 ;
    wire new_AGEMA_signal_13819 ;
    wire new_AGEMA_signal_13820 ;
    wire new_AGEMA_signal_13821 ;
    wire new_AGEMA_signal_13822 ;
    wire new_AGEMA_signal_13823 ;
    wire new_AGEMA_signal_13824 ;
    wire new_AGEMA_signal_13825 ;
    wire new_AGEMA_signal_13826 ;
    wire new_AGEMA_signal_13827 ;
    wire new_AGEMA_signal_13828 ;
    wire new_AGEMA_signal_13829 ;
    wire new_AGEMA_signal_13830 ;
    wire new_AGEMA_signal_13831 ;
    wire new_AGEMA_signal_13832 ;
    wire new_AGEMA_signal_13833 ;
    wire new_AGEMA_signal_13834 ;
    wire new_AGEMA_signal_13835 ;
    wire new_AGEMA_signal_13836 ;
    wire new_AGEMA_signal_13837 ;
    wire new_AGEMA_signal_13838 ;
    wire new_AGEMA_signal_13839 ;
    wire new_AGEMA_signal_13840 ;
    wire new_AGEMA_signal_13841 ;
    wire new_AGEMA_signal_13842 ;
    wire new_AGEMA_signal_13843 ;
    wire new_AGEMA_signal_13844 ;
    wire new_AGEMA_signal_13845 ;
    wire new_AGEMA_signal_13846 ;
    wire new_AGEMA_signal_13847 ;
    wire new_AGEMA_signal_13848 ;
    wire new_AGEMA_signal_13849 ;
    wire new_AGEMA_signal_13850 ;
    wire new_AGEMA_signal_13851 ;
    wire new_AGEMA_signal_13852 ;
    wire new_AGEMA_signal_13853 ;
    wire new_AGEMA_signal_13854 ;
    wire new_AGEMA_signal_13855 ;
    wire new_AGEMA_signal_13856 ;
    wire new_AGEMA_signal_13857 ;
    wire new_AGEMA_signal_13858 ;
    wire new_AGEMA_signal_13859 ;
    wire new_AGEMA_signal_13860 ;
    wire new_AGEMA_signal_13861 ;
    wire new_AGEMA_signal_13862 ;
    wire new_AGEMA_signal_13863 ;
    wire new_AGEMA_signal_13864 ;
    wire new_AGEMA_signal_13865 ;
    wire new_AGEMA_signal_13866 ;
    wire new_AGEMA_signal_13867 ;
    wire new_AGEMA_signal_13868 ;
    wire new_AGEMA_signal_13869 ;
    wire new_AGEMA_signal_13870 ;
    wire new_AGEMA_signal_13871 ;
    wire new_AGEMA_signal_13872 ;
    wire new_AGEMA_signal_13873 ;
    wire new_AGEMA_signal_13874 ;
    wire new_AGEMA_signal_13875 ;
    wire new_AGEMA_signal_13876 ;
    wire new_AGEMA_signal_13877 ;
    wire new_AGEMA_signal_13878 ;
    wire new_AGEMA_signal_13879 ;
    wire new_AGEMA_signal_13880 ;
    wire new_AGEMA_signal_13881 ;
    wire new_AGEMA_signal_13882 ;
    wire new_AGEMA_signal_13883 ;
    wire new_AGEMA_signal_13884 ;
    wire new_AGEMA_signal_13885 ;
    wire new_AGEMA_signal_13886 ;
    wire new_AGEMA_signal_13887 ;
    wire new_AGEMA_signal_13888 ;
    wire new_AGEMA_signal_13889 ;
    wire new_AGEMA_signal_13890 ;
    wire new_AGEMA_signal_13894 ;
    wire new_AGEMA_signal_13895 ;
    wire new_AGEMA_signal_13896 ;
    wire new_AGEMA_signal_13900 ;
    wire new_AGEMA_signal_13901 ;
    wire new_AGEMA_signal_13902 ;
    wire new_AGEMA_signal_13906 ;
    wire new_AGEMA_signal_13907 ;
    wire new_AGEMA_signal_13908 ;
    wire new_AGEMA_signal_13912 ;
    wire new_AGEMA_signal_13913 ;
    wire new_AGEMA_signal_13914 ;
    wire new_AGEMA_signal_13918 ;
    wire new_AGEMA_signal_13919 ;
    wire new_AGEMA_signal_13920 ;
    wire new_AGEMA_signal_13924 ;
    wire new_AGEMA_signal_13925 ;
    wire new_AGEMA_signal_13926 ;
    wire new_AGEMA_signal_13930 ;
    wire new_AGEMA_signal_13931 ;
    wire new_AGEMA_signal_13932 ;
    wire new_AGEMA_signal_13936 ;
    wire new_AGEMA_signal_13937 ;
    wire new_AGEMA_signal_13938 ;
    wire new_AGEMA_signal_13942 ;
    wire new_AGEMA_signal_13943 ;
    wire new_AGEMA_signal_13944 ;
    wire new_AGEMA_signal_13948 ;
    wire new_AGEMA_signal_13949 ;
    wire new_AGEMA_signal_13950 ;
    wire new_AGEMA_signal_13954 ;
    wire new_AGEMA_signal_13955 ;
    wire new_AGEMA_signal_13956 ;
    wire new_AGEMA_signal_13960 ;
    wire new_AGEMA_signal_13961 ;
    wire new_AGEMA_signal_13962 ;
    wire new_AGEMA_signal_13966 ;
    wire new_AGEMA_signal_13967 ;
    wire new_AGEMA_signal_13968 ;
    wire new_AGEMA_signal_13972 ;
    wire new_AGEMA_signal_13973 ;
    wire new_AGEMA_signal_13974 ;
    wire new_AGEMA_signal_13978 ;
    wire new_AGEMA_signal_13979 ;
    wire new_AGEMA_signal_13980 ;
    wire new_AGEMA_signal_13984 ;
    wire new_AGEMA_signal_13985 ;
    wire new_AGEMA_signal_13986 ;
    wire new_AGEMA_signal_13990 ;
    wire new_AGEMA_signal_13991 ;
    wire new_AGEMA_signal_13992 ;
    wire new_AGEMA_signal_13996 ;
    wire new_AGEMA_signal_13997 ;
    wire new_AGEMA_signal_13998 ;
    wire new_AGEMA_signal_14002 ;
    wire new_AGEMA_signal_14003 ;
    wire new_AGEMA_signal_14004 ;
    wire new_AGEMA_signal_14008 ;
    wire new_AGEMA_signal_14009 ;
    wire new_AGEMA_signal_14010 ;
    wire new_AGEMA_signal_14014 ;
    wire new_AGEMA_signal_14015 ;
    wire new_AGEMA_signal_14016 ;
    wire new_AGEMA_signal_14020 ;
    wire new_AGEMA_signal_14021 ;
    wire new_AGEMA_signal_14022 ;
    wire new_AGEMA_signal_14026 ;
    wire new_AGEMA_signal_14027 ;
    wire new_AGEMA_signal_14028 ;
    wire new_AGEMA_signal_14032 ;
    wire new_AGEMA_signal_14033 ;
    wire new_AGEMA_signal_14034 ;
    wire new_AGEMA_signal_14038 ;
    wire new_AGEMA_signal_14039 ;
    wire new_AGEMA_signal_14040 ;
    wire new_AGEMA_signal_14041 ;
    wire new_AGEMA_signal_14042 ;
    wire new_AGEMA_signal_14043 ;
    wire new_AGEMA_signal_14044 ;
    wire new_AGEMA_signal_14045 ;
    wire new_AGEMA_signal_14046 ;
    wire new_AGEMA_signal_14047 ;
    wire new_AGEMA_signal_14048 ;
    wire new_AGEMA_signal_14049 ;
    wire new_AGEMA_signal_14050 ;
    wire new_AGEMA_signal_14051 ;
    wire new_AGEMA_signal_14052 ;
    wire new_AGEMA_signal_14053 ;
    wire new_AGEMA_signal_14054 ;
    wire new_AGEMA_signal_14055 ;
    wire new_AGEMA_signal_14056 ;
    wire new_AGEMA_signal_14057 ;
    wire new_AGEMA_signal_14058 ;
    wire new_AGEMA_signal_14059 ;
    wire new_AGEMA_signal_14060 ;
    wire new_AGEMA_signal_14061 ;
    wire new_AGEMA_signal_14062 ;
    wire new_AGEMA_signal_14063 ;
    wire new_AGEMA_signal_14064 ;
    wire new_AGEMA_signal_14065 ;
    wire new_AGEMA_signal_14066 ;
    wire new_AGEMA_signal_14067 ;
    wire new_AGEMA_signal_14068 ;
    wire new_AGEMA_signal_14069 ;
    wire new_AGEMA_signal_14070 ;
    wire new_AGEMA_signal_14071 ;
    wire new_AGEMA_signal_14072 ;
    wire new_AGEMA_signal_14073 ;
    wire new_AGEMA_signal_14074 ;
    wire new_AGEMA_signal_14075 ;
    wire new_AGEMA_signal_14076 ;
    wire new_AGEMA_signal_14077 ;
    wire new_AGEMA_signal_14078 ;
    wire new_AGEMA_signal_14079 ;
    wire new_AGEMA_signal_14080 ;
    wire new_AGEMA_signal_14081 ;
    wire new_AGEMA_signal_14082 ;
    wire new_AGEMA_signal_14083 ;
    wire new_AGEMA_signal_14084 ;
    wire new_AGEMA_signal_14085 ;
    wire new_AGEMA_signal_14086 ;
    wire new_AGEMA_signal_14087 ;
    wire new_AGEMA_signal_14088 ;
    wire new_AGEMA_signal_14089 ;
    wire new_AGEMA_signal_14090 ;
    wire new_AGEMA_signal_14091 ;
    wire new_AGEMA_signal_14092 ;
    wire new_AGEMA_signal_14093 ;
    wire new_AGEMA_signal_14094 ;
    wire new_AGEMA_signal_14095 ;
    wire new_AGEMA_signal_14096 ;
    wire new_AGEMA_signal_14097 ;
    wire new_AGEMA_signal_14098 ;
    wire new_AGEMA_signal_14099 ;
    wire new_AGEMA_signal_14100 ;
    wire new_AGEMA_signal_14101 ;
    wire new_AGEMA_signal_14102 ;
    wire new_AGEMA_signal_14103 ;
    wire new_AGEMA_signal_14104 ;
    wire new_AGEMA_signal_14105 ;
    wire new_AGEMA_signal_14106 ;
    wire new_AGEMA_signal_14107 ;
    wire new_AGEMA_signal_14108 ;
    wire new_AGEMA_signal_14109 ;
    wire new_AGEMA_signal_14110 ;
    wire new_AGEMA_signal_14111 ;
    wire new_AGEMA_signal_14112 ;
    wire new_AGEMA_signal_14113 ;
    wire new_AGEMA_signal_14114 ;
    wire new_AGEMA_signal_14115 ;
    wire new_AGEMA_signal_14116 ;
    wire new_AGEMA_signal_14117 ;
    wire new_AGEMA_signal_14118 ;
    wire new_AGEMA_signal_14119 ;
    wire new_AGEMA_signal_14120 ;
    wire new_AGEMA_signal_14121 ;
    wire new_AGEMA_signal_14122 ;
    wire new_AGEMA_signal_14123 ;
    wire new_AGEMA_signal_14124 ;
    wire new_AGEMA_signal_14125 ;
    wire new_AGEMA_signal_14126 ;
    wire new_AGEMA_signal_14127 ;
    wire new_AGEMA_signal_14128 ;
    wire new_AGEMA_signal_14129 ;
    wire new_AGEMA_signal_14130 ;
    wire new_AGEMA_signal_14131 ;
    wire new_AGEMA_signal_14132 ;
    wire new_AGEMA_signal_14133 ;
    wire new_AGEMA_signal_14134 ;
    wire new_AGEMA_signal_14135 ;
    wire new_AGEMA_signal_14136 ;
    wire new_AGEMA_signal_14137 ;
    wire new_AGEMA_signal_14138 ;
    wire new_AGEMA_signal_14139 ;
    wire new_AGEMA_signal_14140 ;
    wire new_AGEMA_signal_14141 ;
    wire new_AGEMA_signal_14142 ;
    wire new_AGEMA_signal_14143 ;
    wire new_AGEMA_signal_14144 ;
    wire new_AGEMA_signal_14145 ;
    wire new_AGEMA_signal_14146 ;
    wire new_AGEMA_signal_14147 ;
    wire new_AGEMA_signal_14148 ;
    wire new_AGEMA_signal_14149 ;
    wire new_AGEMA_signal_14150 ;
    wire new_AGEMA_signal_14151 ;
    wire new_AGEMA_signal_14152 ;
    wire new_AGEMA_signal_14153 ;
    wire new_AGEMA_signal_14154 ;
    wire new_AGEMA_signal_14155 ;
    wire new_AGEMA_signal_14156 ;
    wire new_AGEMA_signal_14157 ;
    wire new_AGEMA_signal_14158 ;
    wire new_AGEMA_signal_14159 ;
    wire new_AGEMA_signal_14160 ;
    wire new_AGEMA_signal_14161 ;
    wire new_AGEMA_signal_14162 ;
    wire new_AGEMA_signal_14163 ;
    wire new_AGEMA_signal_14164 ;
    wire new_AGEMA_signal_14165 ;
    wire new_AGEMA_signal_14166 ;
    wire new_AGEMA_signal_14167 ;
    wire new_AGEMA_signal_14168 ;
    wire new_AGEMA_signal_14169 ;
    wire new_AGEMA_signal_14170 ;
    wire new_AGEMA_signal_14171 ;
    wire new_AGEMA_signal_14172 ;
    wire new_AGEMA_signal_14173 ;
    wire new_AGEMA_signal_14174 ;
    wire new_AGEMA_signal_14175 ;
    wire new_AGEMA_signal_14176 ;
    wire new_AGEMA_signal_14177 ;
    wire new_AGEMA_signal_14178 ;
    wire new_AGEMA_signal_14179 ;
    wire new_AGEMA_signal_14180 ;
    wire new_AGEMA_signal_14181 ;
    wire new_AGEMA_signal_14182 ;
    wire new_AGEMA_signal_14183 ;
    wire new_AGEMA_signal_14184 ;
    wire new_AGEMA_signal_14185 ;
    wire new_AGEMA_signal_14186 ;
    wire new_AGEMA_signal_14187 ;
    wire new_AGEMA_signal_14188 ;
    wire new_AGEMA_signal_14189 ;
    wire new_AGEMA_signal_14190 ;
    wire new_AGEMA_signal_14191 ;
    wire new_AGEMA_signal_14192 ;
    wire new_AGEMA_signal_14193 ;
    wire new_AGEMA_signal_14194 ;
    wire new_AGEMA_signal_14195 ;
    wire new_AGEMA_signal_14196 ;
    wire new_AGEMA_signal_14197 ;
    wire new_AGEMA_signal_14198 ;
    wire new_AGEMA_signal_14199 ;
    wire new_AGEMA_signal_14200 ;
    wire new_AGEMA_signal_14201 ;
    wire new_AGEMA_signal_14202 ;
    wire new_AGEMA_signal_14203 ;
    wire new_AGEMA_signal_14204 ;
    wire new_AGEMA_signal_14205 ;
    wire new_AGEMA_signal_14206 ;
    wire new_AGEMA_signal_14207 ;
    wire new_AGEMA_signal_14208 ;
    wire new_AGEMA_signal_14209 ;
    wire new_AGEMA_signal_14210 ;
    wire new_AGEMA_signal_14211 ;
    wire new_AGEMA_signal_14212 ;
    wire new_AGEMA_signal_14213 ;
    wire new_AGEMA_signal_14214 ;
    wire new_AGEMA_signal_14215 ;
    wire new_AGEMA_signal_14216 ;
    wire new_AGEMA_signal_14217 ;
    wire new_AGEMA_signal_14218 ;
    wire new_AGEMA_signal_14219 ;
    wire new_AGEMA_signal_14220 ;
    wire new_AGEMA_signal_14221 ;
    wire new_AGEMA_signal_14222 ;
    wire new_AGEMA_signal_14223 ;
    wire new_AGEMA_signal_14224 ;
    wire new_AGEMA_signal_14225 ;
    wire new_AGEMA_signal_14226 ;
    wire new_AGEMA_signal_14227 ;
    wire new_AGEMA_signal_14228 ;
    wire new_AGEMA_signal_14229 ;
    wire new_AGEMA_signal_14230 ;
    wire new_AGEMA_signal_14231 ;
    wire new_AGEMA_signal_14232 ;
    wire new_AGEMA_signal_14233 ;
    wire new_AGEMA_signal_14234 ;
    wire new_AGEMA_signal_14235 ;
    wire new_AGEMA_signal_14236 ;
    wire new_AGEMA_signal_14237 ;
    wire new_AGEMA_signal_14238 ;
    wire new_AGEMA_signal_14239 ;
    wire new_AGEMA_signal_14240 ;
    wire new_AGEMA_signal_14241 ;
    wire new_AGEMA_signal_14242 ;
    wire new_AGEMA_signal_14243 ;
    wire new_AGEMA_signal_14244 ;
    wire new_AGEMA_signal_14245 ;
    wire new_AGEMA_signal_14246 ;
    wire new_AGEMA_signal_14247 ;
    wire new_AGEMA_signal_14248 ;
    wire new_AGEMA_signal_14249 ;
    wire new_AGEMA_signal_14250 ;
    wire new_AGEMA_signal_14251 ;
    wire new_AGEMA_signal_14252 ;
    wire new_AGEMA_signal_14253 ;
    wire new_AGEMA_signal_14254 ;
    wire new_AGEMA_signal_14255 ;
    wire new_AGEMA_signal_14256 ;
    wire new_AGEMA_signal_14257 ;
    wire new_AGEMA_signal_14258 ;
    wire new_AGEMA_signal_14259 ;
    wire new_AGEMA_signal_14260 ;
    wire new_AGEMA_signal_14261 ;
    wire new_AGEMA_signal_14262 ;
    wire new_AGEMA_signal_14263 ;
    wire new_AGEMA_signal_14264 ;
    wire new_AGEMA_signal_14265 ;
    wire new_AGEMA_signal_14266 ;
    wire new_AGEMA_signal_14267 ;
    wire new_AGEMA_signal_14268 ;
    wire new_AGEMA_signal_14269 ;
    wire new_AGEMA_signal_14270 ;
    wire new_AGEMA_signal_14271 ;
    wire new_AGEMA_signal_14272 ;
    wire new_AGEMA_signal_14273 ;
    wire new_AGEMA_signal_14274 ;
    wire new_AGEMA_signal_14275 ;
    wire new_AGEMA_signal_14276 ;
    wire new_AGEMA_signal_14277 ;
    wire new_AGEMA_signal_14278 ;
    wire new_AGEMA_signal_14279 ;
    wire new_AGEMA_signal_14280 ;
    wire new_AGEMA_signal_14281 ;
    wire new_AGEMA_signal_14282 ;
    wire new_AGEMA_signal_14283 ;
    wire new_AGEMA_signal_14284 ;
    wire new_AGEMA_signal_14285 ;
    wire new_AGEMA_signal_14286 ;
    wire new_AGEMA_signal_14287 ;
    wire new_AGEMA_signal_14288 ;
    wire new_AGEMA_signal_14289 ;
    wire new_AGEMA_signal_14290 ;
    wire new_AGEMA_signal_14291 ;
    wire new_AGEMA_signal_14292 ;
    wire new_AGEMA_signal_14293 ;
    wire new_AGEMA_signal_14294 ;
    wire new_AGEMA_signal_14295 ;
    wire new_AGEMA_signal_14296 ;
    wire new_AGEMA_signal_14297 ;
    wire new_AGEMA_signal_14298 ;
    wire new_AGEMA_signal_14299 ;
    wire new_AGEMA_signal_14300 ;
    wire new_AGEMA_signal_14301 ;
    wire new_AGEMA_signal_14302 ;
    wire new_AGEMA_signal_14303 ;
    wire new_AGEMA_signal_14304 ;
    wire new_AGEMA_signal_14305 ;
    wire new_AGEMA_signal_14306 ;
    wire new_AGEMA_signal_14307 ;
    wire new_AGEMA_signal_14308 ;
    wire new_AGEMA_signal_14309 ;
    wire new_AGEMA_signal_14310 ;
    wire new_AGEMA_signal_14311 ;
    wire new_AGEMA_signal_14312 ;
    wire new_AGEMA_signal_14313 ;
    wire new_AGEMA_signal_14314 ;
    wire new_AGEMA_signal_14315 ;
    wire new_AGEMA_signal_14316 ;
    wire new_AGEMA_signal_14317 ;
    wire new_AGEMA_signal_14318 ;
    wire new_AGEMA_signal_14319 ;
    wire new_AGEMA_signal_14320 ;
    wire new_AGEMA_signal_14321 ;
    wire new_AGEMA_signal_14322 ;
    wire new_AGEMA_signal_14323 ;
    wire new_AGEMA_signal_14324 ;
    wire new_AGEMA_signal_14325 ;
    wire new_AGEMA_signal_14326 ;
    wire new_AGEMA_signal_14327 ;
    wire new_AGEMA_signal_14328 ;
    wire new_AGEMA_signal_14329 ;
    wire new_AGEMA_signal_14330 ;
    wire new_AGEMA_signal_14331 ;
    wire new_AGEMA_signal_14332 ;
    wire new_AGEMA_signal_14333 ;
    wire new_AGEMA_signal_14334 ;
    wire new_AGEMA_signal_14335 ;
    wire new_AGEMA_signal_14336 ;
    wire new_AGEMA_signal_14337 ;
    wire new_AGEMA_signal_14338 ;
    wire new_AGEMA_signal_14339 ;
    wire new_AGEMA_signal_14340 ;
    wire new_AGEMA_signal_14341 ;
    wire new_AGEMA_signal_14342 ;
    wire new_AGEMA_signal_14343 ;
    wire new_AGEMA_signal_14344 ;
    wire new_AGEMA_signal_14345 ;
    wire new_AGEMA_signal_14346 ;
    wire new_AGEMA_signal_14347 ;
    wire new_AGEMA_signal_14348 ;
    wire new_AGEMA_signal_14349 ;
    wire new_AGEMA_signal_14350 ;
    wire new_AGEMA_signal_14351 ;
    wire new_AGEMA_signal_14352 ;
    wire new_AGEMA_signal_14353 ;
    wire new_AGEMA_signal_14354 ;
    wire new_AGEMA_signal_14355 ;
    wire new_AGEMA_signal_14356 ;
    wire new_AGEMA_signal_14357 ;
    wire new_AGEMA_signal_14358 ;
    wire new_AGEMA_signal_14359 ;
    wire new_AGEMA_signal_14360 ;
    wire new_AGEMA_signal_14361 ;
    wire new_AGEMA_signal_14362 ;
    wire new_AGEMA_signal_14363 ;
    wire new_AGEMA_signal_14364 ;
    wire new_AGEMA_signal_14365 ;
    wire new_AGEMA_signal_14366 ;
    wire new_AGEMA_signal_14367 ;
    wire new_AGEMA_signal_14368 ;
    wire new_AGEMA_signal_14369 ;
    wire new_AGEMA_signal_14370 ;
    wire new_AGEMA_signal_14371 ;
    wire new_AGEMA_signal_14372 ;
    wire new_AGEMA_signal_14373 ;
    wire new_AGEMA_signal_14374 ;
    wire new_AGEMA_signal_14375 ;
    wire new_AGEMA_signal_14376 ;
    wire new_AGEMA_signal_14377 ;
    wire new_AGEMA_signal_14378 ;
    wire new_AGEMA_signal_14379 ;
    wire new_AGEMA_signal_14380 ;
    wire new_AGEMA_signal_14381 ;
    wire new_AGEMA_signal_14382 ;
    wire new_AGEMA_signal_14383 ;
    wire new_AGEMA_signal_14384 ;
    wire new_AGEMA_signal_14385 ;
    wire new_AGEMA_signal_14386 ;
    wire new_AGEMA_signal_14387 ;
    wire new_AGEMA_signal_14388 ;
    wire new_AGEMA_signal_14389 ;
    wire new_AGEMA_signal_14390 ;
    wire new_AGEMA_signal_14391 ;
    wire new_AGEMA_signal_14392 ;
    wire new_AGEMA_signal_14393 ;
    wire new_AGEMA_signal_14394 ;
    wire new_AGEMA_signal_14395 ;
    wire new_AGEMA_signal_14396 ;
    wire new_AGEMA_signal_14397 ;
    wire new_AGEMA_signal_14398 ;
    wire new_AGEMA_signal_14399 ;
    wire new_AGEMA_signal_14400 ;
    wire new_AGEMA_signal_14401 ;
    wire new_AGEMA_signal_14402 ;
    wire new_AGEMA_signal_14403 ;
    wire new_AGEMA_signal_14404 ;
    wire new_AGEMA_signal_14405 ;
    wire new_AGEMA_signal_14406 ;
    wire new_AGEMA_signal_14407 ;
    wire new_AGEMA_signal_14408 ;
    wire new_AGEMA_signal_14409 ;
    wire new_AGEMA_signal_14410 ;
    wire new_AGEMA_signal_14411 ;
    wire new_AGEMA_signal_14412 ;
    wire new_AGEMA_signal_14413 ;
    wire new_AGEMA_signal_14414 ;
    wire new_AGEMA_signal_14415 ;
    wire new_AGEMA_signal_14416 ;
    wire new_AGEMA_signal_14417 ;
    wire new_AGEMA_signal_14418 ;
    wire new_AGEMA_signal_14419 ;
    wire new_AGEMA_signal_14420 ;
    wire new_AGEMA_signal_14421 ;
    wire new_AGEMA_signal_14422 ;
    wire new_AGEMA_signal_14423 ;
    wire new_AGEMA_signal_14424 ;
    wire new_AGEMA_signal_14425 ;
    wire new_AGEMA_signal_14426 ;
    wire new_AGEMA_signal_14427 ;
    wire new_AGEMA_signal_14428 ;
    wire new_AGEMA_signal_14429 ;
    wire new_AGEMA_signal_14430 ;
    wire new_AGEMA_signal_14431 ;
    wire new_AGEMA_signal_14432 ;
    wire new_AGEMA_signal_14433 ;
    wire new_AGEMA_signal_14434 ;
    wire new_AGEMA_signal_14435 ;
    wire new_AGEMA_signal_14436 ;
    wire new_AGEMA_signal_14437 ;
    wire new_AGEMA_signal_14438 ;
    wire new_AGEMA_signal_14439 ;
    wire new_AGEMA_signal_14440 ;
    wire new_AGEMA_signal_14441 ;
    wire new_AGEMA_signal_14442 ;
    wire new_AGEMA_signal_14443 ;
    wire new_AGEMA_signal_14444 ;
    wire new_AGEMA_signal_14445 ;
    wire new_AGEMA_signal_14446 ;
    wire new_AGEMA_signal_14447 ;
    wire new_AGEMA_signal_14448 ;
    wire new_AGEMA_signal_14449 ;
    wire new_AGEMA_signal_14450 ;
    wire new_AGEMA_signal_14451 ;
    wire new_AGEMA_signal_14452 ;
    wire new_AGEMA_signal_14453 ;
    wire new_AGEMA_signal_14454 ;
    wire new_AGEMA_signal_14455 ;
    wire new_AGEMA_signal_14456 ;
    wire new_AGEMA_signal_14457 ;
    wire new_AGEMA_signal_14458 ;
    wire new_AGEMA_signal_14459 ;
    wire new_AGEMA_signal_14460 ;
    wire new_AGEMA_signal_14461 ;
    wire new_AGEMA_signal_14462 ;
    wire new_AGEMA_signal_14463 ;
    wire new_AGEMA_signal_14464 ;
    wire new_AGEMA_signal_14465 ;
    wire new_AGEMA_signal_14466 ;
    wire new_AGEMA_signal_14467 ;
    wire new_AGEMA_signal_14468 ;
    wire new_AGEMA_signal_14469 ;
    wire new_AGEMA_signal_14470 ;
    wire new_AGEMA_signal_14471 ;
    wire new_AGEMA_signal_14472 ;
    wire new_AGEMA_signal_14473 ;
    wire new_AGEMA_signal_14474 ;
    wire new_AGEMA_signal_14475 ;
    wire new_AGEMA_signal_14476 ;
    wire new_AGEMA_signal_14477 ;
    wire new_AGEMA_signal_14478 ;
    wire new_AGEMA_signal_14479 ;
    wire new_AGEMA_signal_14480 ;
    wire new_AGEMA_signal_14481 ;
    wire new_AGEMA_signal_14482 ;
    wire new_AGEMA_signal_14483 ;
    wire new_AGEMA_signal_14484 ;
    wire new_AGEMA_signal_14485 ;
    wire new_AGEMA_signal_14486 ;
    wire new_AGEMA_signal_14487 ;
    wire new_AGEMA_signal_14488 ;
    wire new_AGEMA_signal_14489 ;
    wire new_AGEMA_signal_14490 ;
    wire new_AGEMA_signal_14491 ;
    wire new_AGEMA_signal_14492 ;
    wire new_AGEMA_signal_14493 ;
    wire new_AGEMA_signal_14494 ;
    wire new_AGEMA_signal_14495 ;
    wire new_AGEMA_signal_14496 ;
    wire new_AGEMA_signal_14497 ;
    wire new_AGEMA_signal_14498 ;
    wire new_AGEMA_signal_14499 ;
    wire new_AGEMA_signal_14500 ;
    wire new_AGEMA_signal_14501 ;
    wire new_AGEMA_signal_14502 ;
    wire new_AGEMA_signal_14503 ;
    wire new_AGEMA_signal_14504 ;
    wire new_AGEMA_signal_14505 ;
    wire new_AGEMA_signal_14506 ;
    wire new_AGEMA_signal_14507 ;
    wire new_AGEMA_signal_14508 ;
    wire new_AGEMA_signal_14509 ;
    wire new_AGEMA_signal_14510 ;
    wire new_AGEMA_signal_14511 ;
    wire new_AGEMA_signal_14512 ;
    wire new_AGEMA_signal_14513 ;
    wire new_AGEMA_signal_14514 ;
    wire new_AGEMA_signal_14515 ;
    wire new_AGEMA_signal_14516 ;
    wire new_AGEMA_signal_14517 ;
    wire new_AGEMA_signal_14518 ;
    wire new_AGEMA_signal_14519 ;
    wire new_AGEMA_signal_14520 ;
    wire new_AGEMA_signal_14524 ;
    wire new_AGEMA_signal_14525 ;
    wire new_AGEMA_signal_14526 ;
    wire new_AGEMA_signal_14530 ;
    wire new_AGEMA_signal_14531 ;
    wire new_AGEMA_signal_14532 ;
    wire new_AGEMA_signal_14536 ;
    wire new_AGEMA_signal_14537 ;
    wire new_AGEMA_signal_14538 ;
    wire new_AGEMA_signal_14542 ;
    wire new_AGEMA_signal_14543 ;
    wire new_AGEMA_signal_14544 ;
    wire new_AGEMA_signal_14548 ;
    wire new_AGEMA_signal_14549 ;
    wire new_AGEMA_signal_14550 ;
    wire new_AGEMA_signal_14554 ;
    wire new_AGEMA_signal_14555 ;
    wire new_AGEMA_signal_14556 ;
    wire new_AGEMA_signal_14560 ;
    wire new_AGEMA_signal_14561 ;
    wire new_AGEMA_signal_14562 ;
    wire new_AGEMA_signal_14566 ;
    wire new_AGEMA_signal_14567 ;
    wire new_AGEMA_signal_14568 ;
    wire new_AGEMA_signal_14572 ;
    wire new_AGEMA_signal_14573 ;
    wire new_AGEMA_signal_14574 ;
    wire new_AGEMA_signal_14578 ;
    wire new_AGEMA_signal_14579 ;
    wire new_AGEMA_signal_14580 ;
    wire new_AGEMA_signal_14584 ;
    wire new_AGEMA_signal_14585 ;
    wire new_AGEMA_signal_14586 ;
    wire new_AGEMA_signal_14590 ;
    wire new_AGEMA_signal_14591 ;
    wire new_AGEMA_signal_14592 ;
    wire new_AGEMA_signal_14596 ;
    wire new_AGEMA_signal_14597 ;
    wire new_AGEMA_signal_14598 ;
    wire new_AGEMA_signal_14602 ;
    wire new_AGEMA_signal_14603 ;
    wire new_AGEMA_signal_14604 ;
    wire new_AGEMA_signal_14608 ;
    wire new_AGEMA_signal_14609 ;
    wire new_AGEMA_signal_14610 ;
    wire new_AGEMA_signal_14614 ;
    wire new_AGEMA_signal_14615 ;
    wire new_AGEMA_signal_14616 ;
    wire new_AGEMA_signal_14620 ;
    wire new_AGEMA_signal_14621 ;
    wire new_AGEMA_signal_14622 ;
    wire new_AGEMA_signal_14626 ;
    wire new_AGEMA_signal_14627 ;
    wire new_AGEMA_signal_14628 ;
    wire new_AGEMA_signal_14632 ;
    wire new_AGEMA_signal_14633 ;
    wire new_AGEMA_signal_14634 ;
    wire new_AGEMA_signal_14638 ;
    wire new_AGEMA_signal_14639 ;
    wire new_AGEMA_signal_14640 ;
    wire new_AGEMA_signal_14644 ;
    wire new_AGEMA_signal_14645 ;
    wire new_AGEMA_signal_14646 ;
    wire new_AGEMA_signal_14650 ;
    wire new_AGEMA_signal_14651 ;
    wire new_AGEMA_signal_14652 ;
    wire new_AGEMA_signal_14656 ;
    wire new_AGEMA_signal_14657 ;
    wire new_AGEMA_signal_14658 ;
    wire new_AGEMA_signal_14662 ;
    wire new_AGEMA_signal_14663 ;
    wire new_AGEMA_signal_14664 ;
    wire new_AGEMA_signal_14668 ;
    wire new_AGEMA_signal_14669 ;
    wire new_AGEMA_signal_14670 ;
    wire new_AGEMA_signal_14674 ;
    wire new_AGEMA_signal_14675 ;
    wire new_AGEMA_signal_14676 ;
    wire new_AGEMA_signal_14680 ;
    wire new_AGEMA_signal_14681 ;
    wire new_AGEMA_signal_14682 ;
    wire new_AGEMA_signal_14686 ;
    wire new_AGEMA_signal_14687 ;
    wire new_AGEMA_signal_14688 ;
    wire new_AGEMA_signal_14692 ;
    wire new_AGEMA_signal_14693 ;
    wire new_AGEMA_signal_14694 ;
    wire new_AGEMA_signal_14698 ;
    wire new_AGEMA_signal_14699 ;
    wire new_AGEMA_signal_14700 ;
    wire new_AGEMA_signal_14704 ;
    wire new_AGEMA_signal_14705 ;
    wire new_AGEMA_signal_14706 ;
    wire new_AGEMA_signal_14710 ;
    wire new_AGEMA_signal_14711 ;
    wire new_AGEMA_signal_14712 ;
    wire new_AGEMA_signal_14713 ;
    wire new_AGEMA_signal_14714 ;
    wire new_AGEMA_signal_14715 ;
    wire new_AGEMA_signal_14716 ;
    wire new_AGEMA_signal_14717 ;
    wire new_AGEMA_signal_14718 ;
    wire new_AGEMA_signal_14719 ;
    wire new_AGEMA_signal_14720 ;
    wire new_AGEMA_signal_14721 ;
    wire new_AGEMA_signal_14722 ;
    wire new_AGEMA_signal_14723 ;
    wire new_AGEMA_signal_14724 ;
    wire new_AGEMA_signal_14725 ;
    wire new_AGEMA_signal_14726 ;
    wire new_AGEMA_signal_14727 ;
    wire new_AGEMA_signal_14728 ;
    wire new_AGEMA_signal_14729 ;
    wire new_AGEMA_signal_14730 ;
    wire new_AGEMA_signal_14731 ;
    wire new_AGEMA_signal_14732 ;
    wire new_AGEMA_signal_14733 ;
    wire new_AGEMA_signal_14734 ;
    wire new_AGEMA_signal_14735 ;
    wire new_AGEMA_signal_14736 ;
    wire new_AGEMA_signal_14737 ;
    wire new_AGEMA_signal_14738 ;
    wire new_AGEMA_signal_14739 ;
    wire new_AGEMA_signal_14740 ;
    wire new_AGEMA_signal_14741 ;
    wire new_AGEMA_signal_14742 ;
    wire new_AGEMA_signal_14743 ;
    wire new_AGEMA_signal_14744 ;
    wire new_AGEMA_signal_14745 ;
    wire new_AGEMA_signal_14746 ;
    wire new_AGEMA_signal_14747 ;
    wire new_AGEMA_signal_14748 ;
    wire new_AGEMA_signal_14749 ;
    wire new_AGEMA_signal_14750 ;
    wire new_AGEMA_signal_14751 ;
    wire new_AGEMA_signal_14752 ;
    wire new_AGEMA_signal_14753 ;
    wire new_AGEMA_signal_14754 ;
    wire new_AGEMA_signal_14755 ;
    wire new_AGEMA_signal_14756 ;
    wire new_AGEMA_signal_14757 ;
    wire new_AGEMA_signal_14758 ;
    wire new_AGEMA_signal_14759 ;
    wire new_AGEMA_signal_14760 ;
    wire new_AGEMA_signal_14761 ;
    wire new_AGEMA_signal_14762 ;
    wire new_AGEMA_signal_14763 ;
    wire new_AGEMA_signal_14764 ;
    wire new_AGEMA_signal_14765 ;
    wire new_AGEMA_signal_14766 ;
    wire new_AGEMA_signal_14767 ;
    wire new_AGEMA_signal_14768 ;
    wire new_AGEMA_signal_14769 ;
    wire new_AGEMA_signal_14770 ;
    wire new_AGEMA_signal_14771 ;
    wire new_AGEMA_signal_14772 ;
    wire new_AGEMA_signal_14773 ;
    wire new_AGEMA_signal_14774 ;
    wire new_AGEMA_signal_14775 ;
    wire new_AGEMA_signal_14776 ;
    wire new_AGEMA_signal_14777 ;
    wire new_AGEMA_signal_14778 ;
    wire new_AGEMA_signal_14779 ;
    wire new_AGEMA_signal_14780 ;
    wire new_AGEMA_signal_14781 ;
    wire new_AGEMA_signal_14782 ;
    wire new_AGEMA_signal_14783 ;
    wire new_AGEMA_signal_14784 ;
    wire new_AGEMA_signal_14785 ;
    wire new_AGEMA_signal_14786 ;
    wire new_AGEMA_signal_14787 ;
    wire new_AGEMA_signal_14788 ;
    wire new_AGEMA_signal_14789 ;
    wire new_AGEMA_signal_14790 ;
    wire new_AGEMA_signal_14791 ;
    wire new_AGEMA_signal_14792 ;
    wire new_AGEMA_signal_14793 ;
    wire new_AGEMA_signal_14794 ;
    wire new_AGEMA_signal_14795 ;
    wire new_AGEMA_signal_14796 ;
    wire new_AGEMA_signal_14797 ;
    wire new_AGEMA_signal_14798 ;
    wire new_AGEMA_signal_14799 ;
    wire new_AGEMA_signal_14800 ;
    wire new_AGEMA_signal_14801 ;
    wire new_AGEMA_signal_14802 ;
    wire new_AGEMA_signal_14803 ;
    wire new_AGEMA_signal_14804 ;
    wire new_AGEMA_signal_14805 ;
    wire new_AGEMA_signal_14806 ;
    wire new_AGEMA_signal_14807 ;
    wire new_AGEMA_signal_14808 ;
    wire new_AGEMA_signal_14809 ;
    wire new_AGEMA_signal_14810 ;
    wire new_AGEMA_signal_14811 ;
    wire new_AGEMA_signal_14812 ;
    wire new_AGEMA_signal_14813 ;
    wire new_AGEMA_signal_14814 ;
    wire new_AGEMA_signal_14815 ;
    wire new_AGEMA_signal_14816 ;
    wire new_AGEMA_signal_14817 ;
    wire new_AGEMA_signal_14818 ;
    wire new_AGEMA_signal_14819 ;
    wire new_AGEMA_signal_14820 ;
    wire new_AGEMA_signal_14821 ;
    wire new_AGEMA_signal_14822 ;
    wire new_AGEMA_signal_14823 ;
    wire new_AGEMA_signal_14824 ;
    wire new_AGEMA_signal_14825 ;
    wire new_AGEMA_signal_14826 ;
    wire new_AGEMA_signal_14827 ;
    wire new_AGEMA_signal_14828 ;
    wire new_AGEMA_signal_14829 ;
    wire new_AGEMA_signal_14830 ;
    wire new_AGEMA_signal_14831 ;
    wire new_AGEMA_signal_14832 ;
    wire new_AGEMA_signal_14833 ;
    wire new_AGEMA_signal_14834 ;
    wire new_AGEMA_signal_14835 ;
    wire new_AGEMA_signal_14836 ;
    wire new_AGEMA_signal_14837 ;
    wire new_AGEMA_signal_14838 ;
    wire new_AGEMA_signal_14839 ;
    wire new_AGEMA_signal_14840 ;
    wire new_AGEMA_signal_14841 ;
    wire new_AGEMA_signal_14842 ;
    wire new_AGEMA_signal_14843 ;
    wire new_AGEMA_signal_14844 ;
    wire new_AGEMA_signal_14845 ;
    wire new_AGEMA_signal_14846 ;
    wire new_AGEMA_signal_14847 ;
    wire new_AGEMA_signal_14848 ;
    wire new_AGEMA_signal_14849 ;
    wire new_AGEMA_signal_14850 ;
    wire new_AGEMA_signal_14851 ;
    wire new_AGEMA_signal_14852 ;
    wire new_AGEMA_signal_14853 ;
    wire new_AGEMA_signal_14854 ;
    wire new_AGEMA_signal_14855 ;
    wire new_AGEMA_signal_14856 ;
    wire new_AGEMA_signal_14857 ;
    wire new_AGEMA_signal_14858 ;
    wire new_AGEMA_signal_14859 ;
    wire new_AGEMA_signal_14860 ;
    wire new_AGEMA_signal_14861 ;
    wire new_AGEMA_signal_14862 ;
    wire new_AGEMA_signal_14863 ;
    wire new_AGEMA_signal_14864 ;
    wire new_AGEMA_signal_14865 ;
    wire new_AGEMA_signal_14866 ;
    wire new_AGEMA_signal_14867 ;
    wire new_AGEMA_signal_14868 ;
    wire new_AGEMA_signal_14869 ;
    wire new_AGEMA_signal_14870 ;
    wire new_AGEMA_signal_14871 ;
    wire new_AGEMA_signal_14872 ;
    wire new_AGEMA_signal_14873 ;
    wire new_AGEMA_signal_14874 ;
    wire new_AGEMA_signal_14875 ;
    wire new_AGEMA_signal_14876 ;
    wire new_AGEMA_signal_14877 ;
    wire new_AGEMA_signal_14878 ;
    wire new_AGEMA_signal_14879 ;
    wire new_AGEMA_signal_14880 ;
    wire new_AGEMA_signal_14881 ;
    wire new_AGEMA_signal_14882 ;
    wire new_AGEMA_signal_14883 ;
    wire new_AGEMA_signal_14884 ;
    wire new_AGEMA_signal_14885 ;
    wire new_AGEMA_signal_14886 ;
    wire new_AGEMA_signal_14887 ;
    wire new_AGEMA_signal_14888 ;
    wire new_AGEMA_signal_14889 ;
    wire new_AGEMA_signal_14890 ;
    wire new_AGEMA_signal_14891 ;
    wire new_AGEMA_signal_14892 ;
    wire new_AGEMA_signal_14893 ;
    wire new_AGEMA_signal_14894 ;
    wire new_AGEMA_signal_14895 ;
    wire new_AGEMA_signal_14896 ;
    wire new_AGEMA_signal_14897 ;
    wire new_AGEMA_signal_14898 ;
    wire new_AGEMA_signal_14899 ;
    wire new_AGEMA_signal_14900 ;
    wire new_AGEMA_signal_14901 ;
    wire new_AGEMA_signal_14902 ;
    wire new_AGEMA_signal_14903 ;
    wire new_AGEMA_signal_14904 ;
    wire new_AGEMA_signal_14905 ;
    wire new_AGEMA_signal_14906 ;
    wire new_AGEMA_signal_14907 ;
    wire new_AGEMA_signal_14908 ;
    wire new_AGEMA_signal_14909 ;
    wire new_AGEMA_signal_14910 ;
    wire new_AGEMA_signal_14911 ;
    wire new_AGEMA_signal_14912 ;
    wire new_AGEMA_signal_14913 ;
    wire new_AGEMA_signal_14914 ;
    wire new_AGEMA_signal_14915 ;
    wire new_AGEMA_signal_14916 ;
    wire new_AGEMA_signal_14917 ;
    wire new_AGEMA_signal_14918 ;
    wire new_AGEMA_signal_14919 ;
    wire new_AGEMA_signal_14920 ;
    wire new_AGEMA_signal_14921 ;
    wire new_AGEMA_signal_14922 ;
    wire new_AGEMA_signal_14923 ;
    wire new_AGEMA_signal_14924 ;
    wire new_AGEMA_signal_14925 ;
    wire new_AGEMA_signal_14926 ;
    wire new_AGEMA_signal_14927 ;
    wire new_AGEMA_signal_14928 ;
    wire new_AGEMA_signal_14929 ;
    wire new_AGEMA_signal_14930 ;
    wire new_AGEMA_signal_14931 ;
    wire new_AGEMA_signal_14932 ;
    wire new_AGEMA_signal_14933 ;
    wire new_AGEMA_signal_14934 ;
    wire new_AGEMA_signal_14935 ;
    wire new_AGEMA_signal_14936 ;
    wire new_AGEMA_signal_14937 ;
    wire new_AGEMA_signal_14938 ;
    wire new_AGEMA_signal_14939 ;
    wire new_AGEMA_signal_14940 ;
    wire new_AGEMA_signal_14941 ;
    wire new_AGEMA_signal_14942 ;
    wire new_AGEMA_signal_14943 ;
    wire new_AGEMA_signal_14944 ;
    wire new_AGEMA_signal_14945 ;
    wire new_AGEMA_signal_14946 ;
    wire new_AGEMA_signal_14947 ;
    wire new_AGEMA_signal_14948 ;
    wire new_AGEMA_signal_14949 ;
    wire new_AGEMA_signal_14950 ;
    wire new_AGEMA_signal_14951 ;
    wire new_AGEMA_signal_14952 ;
    wire new_AGEMA_signal_14953 ;
    wire new_AGEMA_signal_14954 ;
    wire new_AGEMA_signal_14955 ;
    wire new_AGEMA_signal_14956 ;
    wire new_AGEMA_signal_14957 ;
    wire new_AGEMA_signal_14958 ;
    wire new_AGEMA_signal_14959 ;
    wire new_AGEMA_signal_14960 ;
    wire new_AGEMA_signal_14961 ;
    wire new_AGEMA_signal_14962 ;
    wire new_AGEMA_signal_14963 ;
    wire new_AGEMA_signal_14964 ;
    wire new_AGEMA_signal_14965 ;
    wire new_AGEMA_signal_14966 ;
    wire new_AGEMA_signal_14967 ;
    wire new_AGEMA_signal_14968 ;
    wire new_AGEMA_signal_14969 ;
    wire new_AGEMA_signal_14970 ;
    wire new_AGEMA_signal_14971 ;
    wire new_AGEMA_signal_14972 ;
    wire new_AGEMA_signal_14973 ;
    wire new_AGEMA_signal_14974 ;
    wire new_AGEMA_signal_14975 ;
    wire new_AGEMA_signal_14976 ;
    wire new_AGEMA_signal_14977 ;
    wire new_AGEMA_signal_14978 ;
    wire new_AGEMA_signal_14979 ;
    wire new_AGEMA_signal_14980 ;
    wire new_AGEMA_signal_14981 ;
    wire new_AGEMA_signal_14982 ;
    wire new_AGEMA_signal_14983 ;
    wire new_AGEMA_signal_14984 ;
    wire new_AGEMA_signal_14985 ;
    wire new_AGEMA_signal_14986 ;
    wire new_AGEMA_signal_14987 ;
    wire new_AGEMA_signal_14988 ;
    wire new_AGEMA_signal_14989 ;
    wire new_AGEMA_signal_14990 ;
    wire new_AGEMA_signal_14991 ;
    wire new_AGEMA_signal_14992 ;
    wire new_AGEMA_signal_14993 ;
    wire new_AGEMA_signal_14994 ;
    wire new_AGEMA_signal_14995 ;
    wire new_AGEMA_signal_14996 ;
    wire new_AGEMA_signal_14997 ;
    wire new_AGEMA_signal_14998 ;
    wire new_AGEMA_signal_14999 ;
    wire new_AGEMA_signal_15000 ;
    wire new_AGEMA_signal_15001 ;
    wire new_AGEMA_signal_15002 ;
    wire new_AGEMA_signal_15003 ;
    wire new_AGEMA_signal_15004 ;
    wire new_AGEMA_signal_15005 ;
    wire new_AGEMA_signal_15006 ;
    wire new_AGEMA_signal_15007 ;
    wire new_AGEMA_signal_15008 ;
    wire new_AGEMA_signal_15009 ;
    wire new_AGEMA_signal_15010 ;
    wire new_AGEMA_signal_15011 ;
    wire new_AGEMA_signal_15012 ;
    wire new_AGEMA_signal_15013 ;
    wire new_AGEMA_signal_15014 ;
    wire new_AGEMA_signal_15015 ;
    wire new_AGEMA_signal_15016 ;
    wire new_AGEMA_signal_15017 ;
    wire new_AGEMA_signal_15018 ;
    wire new_AGEMA_signal_15019 ;
    wire new_AGEMA_signal_15020 ;
    wire new_AGEMA_signal_15021 ;
    wire new_AGEMA_signal_15022 ;
    wire new_AGEMA_signal_15023 ;
    wire new_AGEMA_signal_15024 ;
    wire new_AGEMA_signal_15025 ;
    wire new_AGEMA_signal_15026 ;
    wire new_AGEMA_signal_15027 ;
    wire new_AGEMA_signal_15028 ;
    wire new_AGEMA_signal_15029 ;
    wire new_AGEMA_signal_15030 ;
    wire new_AGEMA_signal_15031 ;
    wire new_AGEMA_signal_15032 ;
    wire new_AGEMA_signal_15033 ;
    wire new_AGEMA_signal_15034 ;
    wire new_AGEMA_signal_15035 ;
    wire new_AGEMA_signal_15036 ;
    wire new_AGEMA_signal_15037 ;
    wire new_AGEMA_signal_15038 ;
    wire new_AGEMA_signal_15039 ;
    wire new_AGEMA_signal_15040 ;
    wire new_AGEMA_signal_15041 ;
    wire new_AGEMA_signal_15042 ;
    wire new_AGEMA_signal_15043 ;
    wire new_AGEMA_signal_15044 ;
    wire new_AGEMA_signal_15045 ;
    wire new_AGEMA_signal_15046 ;
    wire new_AGEMA_signal_15047 ;
    wire new_AGEMA_signal_15048 ;
    wire new_AGEMA_signal_15049 ;
    wire new_AGEMA_signal_15050 ;
    wire new_AGEMA_signal_15051 ;
    wire new_AGEMA_signal_15052 ;
    wire new_AGEMA_signal_15053 ;
    wire new_AGEMA_signal_15054 ;
    wire new_AGEMA_signal_15055 ;
    wire new_AGEMA_signal_15056 ;
    wire new_AGEMA_signal_15057 ;
    wire new_AGEMA_signal_15058 ;
    wire new_AGEMA_signal_15059 ;
    wire new_AGEMA_signal_15060 ;
    wire new_AGEMA_signal_15061 ;
    wire new_AGEMA_signal_15062 ;
    wire new_AGEMA_signal_15063 ;
    wire new_AGEMA_signal_15064 ;
    wire new_AGEMA_signal_15065 ;
    wire new_AGEMA_signal_15066 ;
    wire new_AGEMA_signal_15067 ;
    wire new_AGEMA_signal_15068 ;
    wire new_AGEMA_signal_15069 ;
    wire new_AGEMA_signal_15070 ;
    wire new_AGEMA_signal_15071 ;
    wire new_AGEMA_signal_15072 ;
    wire new_AGEMA_signal_15073 ;
    wire new_AGEMA_signal_15074 ;
    wire new_AGEMA_signal_15075 ;
    wire new_AGEMA_signal_15076 ;
    wire new_AGEMA_signal_15077 ;
    wire new_AGEMA_signal_15078 ;
    wire new_AGEMA_signal_15079 ;
    wire new_AGEMA_signal_15080 ;
    wire new_AGEMA_signal_15081 ;
    wire new_AGEMA_signal_15082 ;
    wire new_AGEMA_signal_15083 ;
    wire new_AGEMA_signal_15084 ;
    wire new_AGEMA_signal_15085 ;
    wire new_AGEMA_signal_15086 ;
    wire new_AGEMA_signal_15087 ;
    wire new_AGEMA_signal_15088 ;
    wire new_AGEMA_signal_15089 ;
    wire new_AGEMA_signal_15090 ;
    wire new_AGEMA_signal_15091 ;
    wire new_AGEMA_signal_15092 ;
    wire new_AGEMA_signal_15093 ;
    wire new_AGEMA_signal_15094 ;
    wire new_AGEMA_signal_15095 ;
    wire new_AGEMA_signal_15096 ;
    wire new_AGEMA_signal_15097 ;
    wire new_AGEMA_signal_15098 ;
    wire new_AGEMA_signal_15099 ;
    wire new_AGEMA_signal_15100 ;
    wire new_AGEMA_signal_15101 ;
    wire new_AGEMA_signal_15102 ;
    wire new_AGEMA_signal_15103 ;
    wire new_AGEMA_signal_15104 ;
    wire new_AGEMA_signal_15105 ;
    wire new_AGEMA_signal_15106 ;
    wire new_AGEMA_signal_15107 ;
    wire new_AGEMA_signal_15108 ;
    wire new_AGEMA_signal_15109 ;
    wire new_AGEMA_signal_15110 ;
    wire new_AGEMA_signal_15111 ;
    wire new_AGEMA_signal_15112 ;
    wire new_AGEMA_signal_15113 ;
    wire new_AGEMA_signal_15114 ;
    wire new_AGEMA_signal_15115 ;
    wire new_AGEMA_signal_15116 ;
    wire new_AGEMA_signal_15117 ;
    wire new_AGEMA_signal_15118 ;
    wire new_AGEMA_signal_15119 ;
    wire new_AGEMA_signal_15120 ;
    wire new_AGEMA_signal_15121 ;
    wire new_AGEMA_signal_15122 ;
    wire new_AGEMA_signal_15123 ;
    wire new_AGEMA_signal_15124 ;
    wire new_AGEMA_signal_15125 ;
    wire new_AGEMA_signal_15126 ;
    wire new_AGEMA_signal_15127 ;
    wire new_AGEMA_signal_15128 ;
    wire new_AGEMA_signal_15129 ;
    wire new_AGEMA_signal_15130 ;
    wire new_AGEMA_signal_15131 ;
    wire new_AGEMA_signal_15132 ;
    wire new_AGEMA_signal_15133 ;
    wire new_AGEMA_signal_15134 ;
    wire new_AGEMA_signal_15135 ;
    wire new_AGEMA_signal_15136 ;
    wire new_AGEMA_signal_15137 ;
    wire new_AGEMA_signal_15138 ;
    wire new_AGEMA_signal_15139 ;
    wire new_AGEMA_signal_15140 ;
    wire new_AGEMA_signal_15141 ;
    wire new_AGEMA_signal_15142 ;
    wire new_AGEMA_signal_15143 ;
    wire new_AGEMA_signal_15144 ;
    wire new_AGEMA_signal_15145 ;
    wire new_AGEMA_signal_15146 ;
    wire new_AGEMA_signal_15147 ;
    wire new_AGEMA_signal_15148 ;
    wire new_AGEMA_signal_15149 ;
    wire new_AGEMA_signal_15150 ;
    wire new_AGEMA_signal_15151 ;
    wire new_AGEMA_signal_15152 ;
    wire new_AGEMA_signal_15153 ;
    wire new_AGEMA_signal_15154 ;
    wire new_AGEMA_signal_15155 ;
    wire new_AGEMA_signal_15156 ;
    wire new_AGEMA_signal_15157 ;
    wire new_AGEMA_signal_15158 ;
    wire new_AGEMA_signal_15159 ;
    wire new_AGEMA_signal_15160 ;
    wire new_AGEMA_signal_15161 ;
    wire new_AGEMA_signal_15162 ;
    wire new_AGEMA_signal_15163 ;
    wire new_AGEMA_signal_15164 ;
    wire new_AGEMA_signal_15165 ;
    wire new_AGEMA_signal_15166 ;
    wire new_AGEMA_signal_15167 ;
    wire new_AGEMA_signal_15168 ;
    wire new_AGEMA_signal_15169 ;
    wire new_AGEMA_signal_15170 ;
    wire new_AGEMA_signal_15171 ;
    wire new_AGEMA_signal_15172 ;
    wire new_AGEMA_signal_15173 ;
    wire new_AGEMA_signal_15174 ;
    wire new_AGEMA_signal_15175 ;
    wire new_AGEMA_signal_15176 ;
    wire new_AGEMA_signal_15177 ;
    wire new_AGEMA_signal_15178 ;
    wire new_AGEMA_signal_15179 ;
    wire new_AGEMA_signal_15180 ;
    wire new_AGEMA_signal_15181 ;
    wire new_AGEMA_signal_15182 ;
    wire new_AGEMA_signal_15183 ;
    wire new_AGEMA_signal_15184 ;
    wire new_AGEMA_signal_15185 ;
    wire new_AGEMA_signal_15186 ;
    wire new_AGEMA_signal_15187 ;
    wire new_AGEMA_signal_15188 ;
    wire new_AGEMA_signal_15189 ;
    wire new_AGEMA_signal_15190 ;
    wire new_AGEMA_signal_15191 ;
    wire new_AGEMA_signal_15192 ;
    wire new_AGEMA_signal_15196 ;
    wire new_AGEMA_signal_15197 ;
    wire new_AGEMA_signal_15198 ;
    wire new_AGEMA_signal_15202 ;
    wire new_AGEMA_signal_15203 ;
    wire new_AGEMA_signal_15204 ;
    wire new_AGEMA_signal_15208 ;
    wire new_AGEMA_signal_15209 ;
    wire new_AGEMA_signal_15210 ;
    wire new_AGEMA_signal_15214 ;
    wire new_AGEMA_signal_15215 ;
    wire new_AGEMA_signal_15216 ;
    wire new_AGEMA_signal_15220 ;
    wire new_AGEMA_signal_15221 ;
    wire new_AGEMA_signal_15222 ;
    wire new_AGEMA_signal_15226 ;
    wire new_AGEMA_signal_15227 ;
    wire new_AGEMA_signal_15228 ;
    wire new_AGEMA_signal_15232 ;
    wire new_AGEMA_signal_15233 ;
    wire new_AGEMA_signal_15234 ;
    wire new_AGEMA_signal_15238 ;
    wire new_AGEMA_signal_15239 ;
    wire new_AGEMA_signal_15240 ;
    wire new_AGEMA_signal_15244 ;
    wire new_AGEMA_signal_15245 ;
    wire new_AGEMA_signal_15246 ;
    wire new_AGEMA_signal_15250 ;
    wire new_AGEMA_signal_15251 ;
    wire new_AGEMA_signal_15252 ;
    wire new_AGEMA_signal_15256 ;
    wire new_AGEMA_signal_15257 ;
    wire new_AGEMA_signal_15258 ;
    wire new_AGEMA_signal_15262 ;
    wire new_AGEMA_signal_15263 ;
    wire new_AGEMA_signal_15264 ;
    wire new_AGEMA_signal_15268 ;
    wire new_AGEMA_signal_15269 ;
    wire new_AGEMA_signal_15270 ;
    wire new_AGEMA_signal_15274 ;
    wire new_AGEMA_signal_15275 ;
    wire new_AGEMA_signal_15276 ;
    wire new_AGEMA_signal_15280 ;
    wire new_AGEMA_signal_15281 ;
    wire new_AGEMA_signal_15282 ;
    wire new_AGEMA_signal_15286 ;
    wire new_AGEMA_signal_15287 ;
    wire new_AGEMA_signal_15288 ;
    wire new_AGEMA_signal_15292 ;
    wire new_AGEMA_signal_15293 ;
    wire new_AGEMA_signal_15294 ;
    wire new_AGEMA_signal_15298 ;
    wire new_AGEMA_signal_15299 ;
    wire new_AGEMA_signal_15300 ;
    wire new_AGEMA_signal_15304 ;
    wire new_AGEMA_signal_15305 ;
    wire new_AGEMA_signal_15306 ;
    wire new_AGEMA_signal_15310 ;
    wire new_AGEMA_signal_15311 ;
    wire new_AGEMA_signal_15312 ;
    wire new_AGEMA_signal_15316 ;
    wire new_AGEMA_signal_15317 ;
    wire new_AGEMA_signal_15318 ;
    wire new_AGEMA_signal_15322 ;
    wire new_AGEMA_signal_15323 ;
    wire new_AGEMA_signal_15324 ;
    wire new_AGEMA_signal_15328 ;
    wire new_AGEMA_signal_15329 ;
    wire new_AGEMA_signal_15330 ;
    wire new_AGEMA_signal_15334 ;
    wire new_AGEMA_signal_15335 ;
    wire new_AGEMA_signal_15336 ;
    wire new_AGEMA_signal_15340 ;
    wire new_AGEMA_signal_15341 ;
    wire new_AGEMA_signal_15342 ;
    wire new_AGEMA_signal_15346 ;
    wire new_AGEMA_signal_15347 ;
    wire new_AGEMA_signal_15348 ;
    wire new_AGEMA_signal_15352 ;
    wire new_AGEMA_signal_15353 ;
    wire new_AGEMA_signal_15354 ;
    wire new_AGEMA_signal_15358 ;
    wire new_AGEMA_signal_15359 ;
    wire new_AGEMA_signal_15360 ;
    wire new_AGEMA_signal_15364 ;
    wire new_AGEMA_signal_15365 ;
    wire new_AGEMA_signal_15366 ;
    wire new_AGEMA_signal_15370 ;
    wire new_AGEMA_signal_15371 ;
    wire new_AGEMA_signal_15372 ;
    wire new_AGEMA_signal_15376 ;
    wire new_AGEMA_signal_15377 ;
    wire new_AGEMA_signal_15378 ;
    wire new_AGEMA_signal_15382 ;
    wire new_AGEMA_signal_15383 ;
    wire new_AGEMA_signal_15384 ;
    wire new_AGEMA_signal_15385 ;
    wire new_AGEMA_signal_15386 ;
    wire new_AGEMA_signal_15387 ;
    wire new_AGEMA_signal_15388 ;
    wire new_AGEMA_signal_15389 ;
    wire new_AGEMA_signal_15390 ;
    wire new_AGEMA_signal_15391 ;
    wire new_AGEMA_signal_15392 ;
    wire new_AGEMA_signal_15393 ;
    wire new_AGEMA_signal_15394 ;
    wire new_AGEMA_signal_15395 ;
    wire new_AGEMA_signal_15396 ;
    wire new_AGEMA_signal_15397 ;
    wire new_AGEMA_signal_15398 ;
    wire new_AGEMA_signal_15399 ;
    wire new_AGEMA_signal_15400 ;
    wire new_AGEMA_signal_15401 ;
    wire new_AGEMA_signal_15402 ;
    wire new_AGEMA_signal_15403 ;
    wire new_AGEMA_signal_15404 ;
    wire new_AGEMA_signal_15405 ;
    wire new_AGEMA_signal_15406 ;
    wire new_AGEMA_signal_15407 ;
    wire new_AGEMA_signal_15408 ;
    wire new_AGEMA_signal_15409 ;
    wire new_AGEMA_signal_15410 ;
    wire new_AGEMA_signal_15411 ;
    wire new_AGEMA_signal_15412 ;
    wire new_AGEMA_signal_15413 ;
    wire new_AGEMA_signal_15414 ;
    wire new_AGEMA_signal_15415 ;
    wire new_AGEMA_signal_15416 ;
    wire new_AGEMA_signal_15417 ;
    wire new_AGEMA_signal_15418 ;
    wire new_AGEMA_signal_15419 ;
    wire new_AGEMA_signal_15420 ;
    wire new_AGEMA_signal_15421 ;
    wire new_AGEMA_signal_15422 ;
    wire new_AGEMA_signal_15423 ;
    wire new_AGEMA_signal_15424 ;
    wire new_AGEMA_signal_15425 ;
    wire new_AGEMA_signal_15426 ;
    wire new_AGEMA_signal_15427 ;
    wire new_AGEMA_signal_15428 ;
    wire new_AGEMA_signal_15429 ;
    wire new_AGEMA_signal_15430 ;
    wire new_AGEMA_signal_15431 ;
    wire new_AGEMA_signal_15432 ;
    wire new_AGEMA_signal_15433 ;
    wire new_AGEMA_signal_15434 ;
    wire new_AGEMA_signal_15435 ;
    wire new_AGEMA_signal_15436 ;
    wire new_AGEMA_signal_15437 ;
    wire new_AGEMA_signal_15438 ;
    wire new_AGEMA_signal_15439 ;
    wire new_AGEMA_signal_15440 ;
    wire new_AGEMA_signal_15441 ;
    wire new_AGEMA_signal_15442 ;
    wire new_AGEMA_signal_15443 ;
    wire new_AGEMA_signal_15444 ;
    wire new_AGEMA_signal_15445 ;
    wire new_AGEMA_signal_15446 ;
    wire new_AGEMA_signal_15447 ;
    wire new_AGEMA_signal_15448 ;
    wire new_AGEMA_signal_15449 ;
    wire new_AGEMA_signal_15450 ;
    wire new_AGEMA_signal_15451 ;
    wire new_AGEMA_signal_15452 ;
    wire new_AGEMA_signal_15453 ;
    wire new_AGEMA_signal_15454 ;
    wire new_AGEMA_signal_15455 ;
    wire new_AGEMA_signal_15456 ;
    wire new_AGEMA_signal_15457 ;
    wire new_AGEMA_signal_15458 ;
    wire new_AGEMA_signal_15459 ;
    wire new_AGEMA_signal_15460 ;
    wire new_AGEMA_signal_15461 ;
    wire new_AGEMA_signal_15462 ;
    wire new_AGEMA_signal_15463 ;
    wire new_AGEMA_signal_15464 ;
    wire new_AGEMA_signal_15465 ;
    wire new_AGEMA_signal_15466 ;
    wire new_AGEMA_signal_15467 ;
    wire new_AGEMA_signal_15468 ;
    wire new_AGEMA_signal_15469 ;
    wire new_AGEMA_signal_15470 ;
    wire new_AGEMA_signal_15471 ;
    wire new_AGEMA_signal_15472 ;
    wire new_AGEMA_signal_15473 ;
    wire new_AGEMA_signal_15474 ;
    wire new_AGEMA_signal_15475 ;
    wire new_AGEMA_signal_15476 ;
    wire new_AGEMA_signal_15477 ;
    wire new_AGEMA_signal_15478 ;
    wire new_AGEMA_signal_15479 ;
    wire new_AGEMA_signal_15480 ;
    wire new_AGEMA_signal_15481 ;
    wire new_AGEMA_signal_15482 ;
    wire new_AGEMA_signal_15483 ;
    wire new_AGEMA_signal_15484 ;
    wire new_AGEMA_signal_15485 ;
    wire new_AGEMA_signal_15486 ;
    wire new_AGEMA_signal_15487 ;
    wire new_AGEMA_signal_15488 ;
    wire new_AGEMA_signal_15489 ;
    wire new_AGEMA_signal_15490 ;
    wire new_AGEMA_signal_15491 ;
    wire new_AGEMA_signal_15492 ;
    wire new_AGEMA_signal_15493 ;
    wire new_AGEMA_signal_15494 ;
    wire new_AGEMA_signal_15495 ;
    wire new_AGEMA_signal_15496 ;
    wire new_AGEMA_signal_15497 ;
    wire new_AGEMA_signal_15498 ;
    wire new_AGEMA_signal_15499 ;
    wire new_AGEMA_signal_15500 ;
    wire new_AGEMA_signal_15501 ;
    wire new_AGEMA_signal_15502 ;
    wire new_AGEMA_signal_15503 ;
    wire new_AGEMA_signal_15504 ;
    wire new_AGEMA_signal_15505 ;
    wire new_AGEMA_signal_15506 ;
    wire new_AGEMA_signal_15507 ;
    wire new_AGEMA_signal_15508 ;
    wire new_AGEMA_signal_15509 ;
    wire new_AGEMA_signal_15510 ;
    wire new_AGEMA_signal_15511 ;
    wire new_AGEMA_signal_15512 ;
    wire new_AGEMA_signal_15513 ;
    wire new_AGEMA_signal_15514 ;
    wire new_AGEMA_signal_15515 ;
    wire new_AGEMA_signal_15516 ;
    wire new_AGEMA_signal_15517 ;
    wire new_AGEMA_signal_15518 ;
    wire new_AGEMA_signal_15519 ;
    wire new_AGEMA_signal_15520 ;
    wire new_AGEMA_signal_15521 ;
    wire new_AGEMA_signal_15522 ;
    wire new_AGEMA_signal_15523 ;
    wire new_AGEMA_signal_15524 ;
    wire new_AGEMA_signal_15525 ;
    wire new_AGEMA_signal_15526 ;
    wire new_AGEMA_signal_15527 ;
    wire new_AGEMA_signal_15528 ;
    wire new_AGEMA_signal_15529 ;
    wire new_AGEMA_signal_15530 ;
    wire new_AGEMA_signal_15531 ;
    wire new_AGEMA_signal_15532 ;
    wire new_AGEMA_signal_15533 ;
    wire new_AGEMA_signal_15534 ;
    wire new_AGEMA_signal_15535 ;
    wire new_AGEMA_signal_15536 ;
    wire new_AGEMA_signal_15537 ;
    wire new_AGEMA_signal_15538 ;
    wire new_AGEMA_signal_15539 ;
    wire new_AGEMA_signal_15540 ;
    wire new_AGEMA_signal_15541 ;
    wire new_AGEMA_signal_15542 ;
    wire new_AGEMA_signal_15543 ;
    wire new_AGEMA_signal_15544 ;
    wire new_AGEMA_signal_15545 ;
    wire new_AGEMA_signal_15546 ;
    wire new_AGEMA_signal_15547 ;
    wire new_AGEMA_signal_15548 ;
    wire new_AGEMA_signal_15549 ;
    wire new_AGEMA_signal_15550 ;
    wire new_AGEMA_signal_15551 ;
    wire new_AGEMA_signal_15552 ;
    wire new_AGEMA_signal_15553 ;
    wire new_AGEMA_signal_15554 ;
    wire new_AGEMA_signal_15555 ;
    wire new_AGEMA_signal_15556 ;
    wire new_AGEMA_signal_15557 ;
    wire new_AGEMA_signal_15558 ;
    wire new_AGEMA_signal_15559 ;
    wire new_AGEMA_signal_15560 ;
    wire new_AGEMA_signal_15561 ;
    wire new_AGEMA_signal_15562 ;
    wire new_AGEMA_signal_15563 ;
    wire new_AGEMA_signal_15564 ;
    wire new_AGEMA_signal_15565 ;
    wire new_AGEMA_signal_15566 ;
    wire new_AGEMA_signal_15567 ;
    wire new_AGEMA_signal_15568 ;
    wire new_AGEMA_signal_15569 ;
    wire new_AGEMA_signal_15570 ;
    wire new_AGEMA_signal_15571 ;
    wire new_AGEMA_signal_15572 ;
    wire new_AGEMA_signal_15573 ;
    wire new_AGEMA_signal_15574 ;
    wire new_AGEMA_signal_15575 ;
    wire new_AGEMA_signal_15576 ;
    wire new_AGEMA_signal_15577 ;
    wire new_AGEMA_signal_15578 ;
    wire new_AGEMA_signal_15579 ;
    wire new_AGEMA_signal_15580 ;
    wire new_AGEMA_signal_15581 ;
    wire new_AGEMA_signal_15582 ;
    wire new_AGEMA_signal_15583 ;
    wire new_AGEMA_signal_15584 ;
    wire new_AGEMA_signal_15585 ;
    wire new_AGEMA_signal_15586 ;
    wire new_AGEMA_signal_15587 ;
    wire new_AGEMA_signal_15588 ;
    wire new_AGEMA_signal_15589 ;
    wire new_AGEMA_signal_15590 ;
    wire new_AGEMA_signal_15591 ;
    wire new_AGEMA_signal_15592 ;
    wire new_AGEMA_signal_15593 ;
    wire new_AGEMA_signal_15594 ;
    wire new_AGEMA_signal_15595 ;
    wire new_AGEMA_signal_15596 ;
    wire new_AGEMA_signal_15597 ;
    wire new_AGEMA_signal_15598 ;
    wire new_AGEMA_signal_15599 ;
    wire new_AGEMA_signal_15600 ;
    wire new_AGEMA_signal_15601 ;
    wire new_AGEMA_signal_15602 ;
    wire new_AGEMA_signal_15603 ;
    wire new_AGEMA_signal_15604 ;
    wire new_AGEMA_signal_15605 ;
    wire new_AGEMA_signal_15606 ;
    wire new_AGEMA_signal_15607 ;
    wire new_AGEMA_signal_15608 ;
    wire new_AGEMA_signal_15609 ;
    wire new_AGEMA_signal_15610 ;
    wire new_AGEMA_signal_15611 ;
    wire new_AGEMA_signal_15612 ;
    wire new_AGEMA_signal_15613 ;
    wire new_AGEMA_signal_15614 ;
    wire new_AGEMA_signal_15615 ;
    wire new_AGEMA_signal_15616 ;
    wire new_AGEMA_signal_15617 ;
    wire new_AGEMA_signal_15618 ;
    wire new_AGEMA_signal_15619 ;
    wire new_AGEMA_signal_15620 ;
    wire new_AGEMA_signal_15621 ;
    wire new_AGEMA_signal_15622 ;
    wire new_AGEMA_signal_15623 ;
    wire new_AGEMA_signal_15624 ;
    wire new_AGEMA_signal_15625 ;
    wire new_AGEMA_signal_15626 ;
    wire new_AGEMA_signal_15627 ;
    wire new_AGEMA_signal_15628 ;
    wire new_AGEMA_signal_15629 ;
    wire new_AGEMA_signal_15630 ;
    wire new_AGEMA_signal_15631 ;
    wire new_AGEMA_signal_15632 ;
    wire new_AGEMA_signal_15633 ;
    wire new_AGEMA_signal_15634 ;
    wire new_AGEMA_signal_15635 ;
    wire new_AGEMA_signal_15636 ;
    wire new_AGEMA_signal_15637 ;
    wire new_AGEMA_signal_15638 ;
    wire new_AGEMA_signal_15639 ;
    wire new_AGEMA_signal_15640 ;
    wire new_AGEMA_signal_15641 ;
    wire new_AGEMA_signal_15642 ;
    wire new_AGEMA_signal_15643 ;
    wire new_AGEMA_signal_15644 ;
    wire new_AGEMA_signal_15645 ;
    wire new_AGEMA_signal_15646 ;
    wire new_AGEMA_signal_15647 ;
    wire new_AGEMA_signal_15648 ;
    wire new_AGEMA_signal_15649 ;
    wire new_AGEMA_signal_15650 ;
    wire new_AGEMA_signal_15651 ;
    wire new_AGEMA_signal_15652 ;
    wire new_AGEMA_signal_15653 ;
    wire new_AGEMA_signal_15654 ;
    wire new_AGEMA_signal_15655 ;
    wire new_AGEMA_signal_15656 ;
    wire new_AGEMA_signal_15657 ;
    wire new_AGEMA_signal_15658 ;
    wire new_AGEMA_signal_15659 ;
    wire new_AGEMA_signal_15660 ;
    wire new_AGEMA_signal_15661 ;
    wire new_AGEMA_signal_15662 ;
    wire new_AGEMA_signal_15663 ;
    wire new_AGEMA_signal_15664 ;
    wire new_AGEMA_signal_15665 ;
    wire new_AGEMA_signal_15666 ;
    wire new_AGEMA_signal_15667 ;
    wire new_AGEMA_signal_15668 ;
    wire new_AGEMA_signal_15669 ;
    wire new_AGEMA_signal_15670 ;
    wire new_AGEMA_signal_15671 ;
    wire new_AGEMA_signal_15672 ;
    wire new_AGEMA_signal_15673 ;
    wire new_AGEMA_signal_15674 ;
    wire new_AGEMA_signal_15675 ;
    wire new_AGEMA_signal_15676 ;
    wire new_AGEMA_signal_15677 ;
    wire new_AGEMA_signal_15678 ;
    wire new_AGEMA_signal_15679 ;
    wire new_AGEMA_signal_15680 ;
    wire new_AGEMA_signal_15681 ;
    wire new_AGEMA_signal_15682 ;
    wire new_AGEMA_signal_15683 ;
    wire new_AGEMA_signal_15684 ;
    wire new_AGEMA_signal_15685 ;
    wire new_AGEMA_signal_15686 ;
    wire new_AGEMA_signal_15687 ;
    wire new_AGEMA_signal_15688 ;
    wire new_AGEMA_signal_15689 ;
    wire new_AGEMA_signal_15690 ;
    wire new_AGEMA_signal_15691 ;
    wire new_AGEMA_signal_15692 ;
    wire new_AGEMA_signal_15693 ;
    wire new_AGEMA_signal_15694 ;
    wire new_AGEMA_signal_15695 ;
    wire new_AGEMA_signal_15696 ;
    wire new_AGEMA_signal_15697 ;
    wire new_AGEMA_signal_15698 ;
    wire new_AGEMA_signal_15699 ;
    wire new_AGEMA_signal_15700 ;
    wire new_AGEMA_signal_15701 ;
    wire new_AGEMA_signal_15702 ;
    wire new_AGEMA_signal_15703 ;
    wire new_AGEMA_signal_15704 ;
    wire new_AGEMA_signal_15705 ;
    wire new_AGEMA_signal_15706 ;
    wire new_AGEMA_signal_15707 ;
    wire new_AGEMA_signal_15708 ;
    wire new_AGEMA_signal_15709 ;
    wire new_AGEMA_signal_15710 ;
    wire new_AGEMA_signal_15711 ;
    wire new_AGEMA_signal_15712 ;
    wire new_AGEMA_signal_15713 ;
    wire new_AGEMA_signal_15714 ;
    wire new_AGEMA_signal_15715 ;
    wire new_AGEMA_signal_15716 ;
    wire new_AGEMA_signal_15717 ;
    wire new_AGEMA_signal_15718 ;
    wire new_AGEMA_signal_15719 ;
    wire new_AGEMA_signal_15720 ;
    wire new_AGEMA_signal_15721 ;
    wire new_AGEMA_signal_15722 ;
    wire new_AGEMA_signal_15723 ;
    wire new_AGEMA_signal_15724 ;
    wire new_AGEMA_signal_15725 ;
    wire new_AGEMA_signal_15726 ;
    wire new_AGEMA_signal_15727 ;
    wire new_AGEMA_signal_15728 ;
    wire new_AGEMA_signal_15729 ;
    wire new_AGEMA_signal_15730 ;
    wire new_AGEMA_signal_15731 ;
    wire new_AGEMA_signal_15732 ;
    wire new_AGEMA_signal_15733 ;
    wire new_AGEMA_signal_15734 ;
    wire new_AGEMA_signal_15735 ;
    wire new_AGEMA_signal_15736 ;
    wire new_AGEMA_signal_15737 ;
    wire new_AGEMA_signal_15738 ;
    wire new_AGEMA_signal_15739 ;
    wire new_AGEMA_signal_15740 ;
    wire new_AGEMA_signal_15741 ;
    wire new_AGEMA_signal_15742 ;
    wire new_AGEMA_signal_15743 ;
    wire new_AGEMA_signal_15744 ;
    wire new_AGEMA_signal_15745 ;
    wire new_AGEMA_signal_15746 ;
    wire new_AGEMA_signal_15747 ;
    wire new_AGEMA_signal_15748 ;
    wire new_AGEMA_signal_15749 ;
    wire new_AGEMA_signal_15750 ;
    wire new_AGEMA_signal_15751 ;
    wire new_AGEMA_signal_15752 ;
    wire new_AGEMA_signal_15753 ;
    wire new_AGEMA_signal_15754 ;
    wire new_AGEMA_signal_15755 ;
    wire new_AGEMA_signal_15756 ;
    wire new_AGEMA_signal_15757 ;
    wire new_AGEMA_signal_15758 ;
    wire new_AGEMA_signal_15759 ;
    wire new_AGEMA_signal_15760 ;
    wire new_AGEMA_signal_15761 ;
    wire new_AGEMA_signal_15762 ;
    wire new_AGEMA_signal_15763 ;
    wire new_AGEMA_signal_15764 ;
    wire new_AGEMA_signal_15765 ;
    wire new_AGEMA_signal_15766 ;
    wire new_AGEMA_signal_15767 ;
    wire new_AGEMA_signal_15768 ;
    wire new_AGEMA_signal_15769 ;
    wire new_AGEMA_signal_15770 ;
    wire new_AGEMA_signal_15771 ;
    wire new_AGEMA_signal_15772 ;
    wire new_AGEMA_signal_15773 ;
    wire new_AGEMA_signal_15774 ;
    wire new_AGEMA_signal_15775 ;
    wire new_AGEMA_signal_15776 ;
    wire new_AGEMA_signal_15777 ;
    wire new_AGEMA_signal_15778 ;
    wire new_AGEMA_signal_15779 ;
    wire new_AGEMA_signal_15780 ;
    wire new_AGEMA_signal_15781 ;
    wire new_AGEMA_signal_15782 ;
    wire new_AGEMA_signal_15783 ;
    wire new_AGEMA_signal_15784 ;
    wire new_AGEMA_signal_15785 ;
    wire new_AGEMA_signal_15786 ;
    wire new_AGEMA_signal_15787 ;
    wire new_AGEMA_signal_15788 ;
    wire new_AGEMA_signal_15789 ;
    wire new_AGEMA_signal_15790 ;
    wire new_AGEMA_signal_15791 ;
    wire new_AGEMA_signal_15792 ;
    wire new_AGEMA_signal_15793 ;
    wire new_AGEMA_signal_15794 ;
    wire new_AGEMA_signal_15795 ;
    wire new_AGEMA_signal_15796 ;
    wire new_AGEMA_signal_15797 ;
    wire new_AGEMA_signal_15798 ;
    wire new_AGEMA_signal_15799 ;
    wire new_AGEMA_signal_15800 ;
    wire new_AGEMA_signal_15801 ;
    wire new_AGEMA_signal_15802 ;
    wire new_AGEMA_signal_15803 ;
    wire new_AGEMA_signal_15804 ;
    wire new_AGEMA_signal_15805 ;
    wire new_AGEMA_signal_15806 ;
    wire new_AGEMA_signal_15807 ;
    wire new_AGEMA_signal_15808 ;
    wire new_AGEMA_signal_15809 ;
    wire new_AGEMA_signal_15810 ;
    wire new_AGEMA_signal_15811 ;
    wire new_AGEMA_signal_15812 ;
    wire new_AGEMA_signal_15813 ;
    wire new_AGEMA_signal_15814 ;
    wire new_AGEMA_signal_15815 ;
    wire new_AGEMA_signal_15816 ;
    wire new_AGEMA_signal_15817 ;
    wire new_AGEMA_signal_15818 ;
    wire new_AGEMA_signal_15819 ;
    wire new_AGEMA_signal_15820 ;
    wire new_AGEMA_signal_15821 ;
    wire new_AGEMA_signal_15822 ;
    wire new_AGEMA_signal_15823 ;
    wire new_AGEMA_signal_15824 ;
    wire new_AGEMA_signal_15825 ;
    wire new_AGEMA_signal_15826 ;
    wire new_AGEMA_signal_15827 ;
    wire new_AGEMA_signal_15828 ;
    wire new_AGEMA_signal_15829 ;
    wire new_AGEMA_signal_15830 ;
    wire new_AGEMA_signal_15831 ;
    wire new_AGEMA_signal_15832 ;
    wire new_AGEMA_signal_15833 ;
    wire new_AGEMA_signal_15834 ;
    wire new_AGEMA_signal_15835 ;
    wire new_AGEMA_signal_15836 ;
    wire new_AGEMA_signal_15837 ;
    wire new_AGEMA_signal_15838 ;
    wire new_AGEMA_signal_15839 ;
    wire new_AGEMA_signal_15840 ;
    wire new_AGEMA_signal_15841 ;
    wire new_AGEMA_signal_15842 ;
    wire new_AGEMA_signal_15843 ;
    wire new_AGEMA_signal_15844 ;
    wire new_AGEMA_signal_15845 ;
    wire new_AGEMA_signal_15846 ;
    wire new_AGEMA_signal_15847 ;
    wire new_AGEMA_signal_15848 ;
    wire new_AGEMA_signal_15849 ;
    wire new_AGEMA_signal_15850 ;
    wire new_AGEMA_signal_15851 ;
    wire new_AGEMA_signal_15852 ;
    wire new_AGEMA_signal_15853 ;
    wire new_AGEMA_signal_15854 ;
    wire new_AGEMA_signal_15855 ;
    wire new_AGEMA_signal_15859 ;
    wire new_AGEMA_signal_15860 ;
    wire new_AGEMA_signal_15861 ;
    wire new_AGEMA_signal_15865 ;
    wire new_AGEMA_signal_15866 ;
    wire new_AGEMA_signal_15867 ;
    wire new_AGEMA_signal_15871 ;
    wire new_AGEMA_signal_15872 ;
    wire new_AGEMA_signal_15873 ;
    wire new_AGEMA_signal_15877 ;
    wire new_AGEMA_signal_15878 ;
    wire new_AGEMA_signal_15879 ;
    wire new_AGEMA_signal_15883 ;
    wire new_AGEMA_signal_15884 ;
    wire new_AGEMA_signal_15885 ;
    wire new_AGEMA_signal_15889 ;
    wire new_AGEMA_signal_15890 ;
    wire new_AGEMA_signal_15891 ;
    wire new_AGEMA_signal_15895 ;
    wire new_AGEMA_signal_15896 ;
    wire new_AGEMA_signal_15897 ;
    wire new_AGEMA_signal_15901 ;
    wire new_AGEMA_signal_15902 ;
    wire new_AGEMA_signal_15903 ;
    wire new_AGEMA_signal_15907 ;
    wire new_AGEMA_signal_15908 ;
    wire new_AGEMA_signal_15909 ;
    wire new_AGEMA_signal_15913 ;
    wire new_AGEMA_signal_15914 ;
    wire new_AGEMA_signal_15915 ;
    wire new_AGEMA_signal_15919 ;
    wire new_AGEMA_signal_15920 ;
    wire new_AGEMA_signal_15921 ;
    wire new_AGEMA_signal_15925 ;
    wire new_AGEMA_signal_15926 ;
    wire new_AGEMA_signal_15927 ;
    wire new_AGEMA_signal_15931 ;
    wire new_AGEMA_signal_15932 ;
    wire new_AGEMA_signal_15933 ;
    wire new_AGEMA_signal_15937 ;
    wire new_AGEMA_signal_15938 ;
    wire new_AGEMA_signal_15939 ;
    wire new_AGEMA_signal_15943 ;
    wire new_AGEMA_signal_15944 ;
    wire new_AGEMA_signal_15945 ;
    wire new_AGEMA_signal_15949 ;
    wire new_AGEMA_signal_15950 ;
    wire new_AGEMA_signal_15951 ;
    wire new_AGEMA_signal_15955 ;
    wire new_AGEMA_signal_15956 ;
    wire new_AGEMA_signal_15957 ;
    wire new_AGEMA_signal_15961 ;
    wire new_AGEMA_signal_15962 ;
    wire new_AGEMA_signal_15963 ;
    wire new_AGEMA_signal_15967 ;
    wire new_AGEMA_signal_15968 ;
    wire new_AGEMA_signal_15969 ;
    wire new_AGEMA_signal_15973 ;
    wire new_AGEMA_signal_15974 ;
    wire new_AGEMA_signal_15975 ;
    wire new_AGEMA_signal_15979 ;
    wire new_AGEMA_signal_15980 ;
    wire new_AGEMA_signal_15981 ;
    wire new_AGEMA_signal_15985 ;
    wire new_AGEMA_signal_15986 ;
    wire new_AGEMA_signal_15987 ;
    wire new_AGEMA_signal_15991 ;
    wire new_AGEMA_signal_15992 ;
    wire new_AGEMA_signal_15993 ;
    wire new_AGEMA_signal_15997 ;
    wire new_AGEMA_signal_15998 ;
    wire new_AGEMA_signal_15999 ;
    wire new_AGEMA_signal_16003 ;
    wire new_AGEMA_signal_16004 ;
    wire new_AGEMA_signal_16005 ;
    wire new_AGEMA_signal_16009 ;
    wire new_AGEMA_signal_16010 ;
    wire new_AGEMA_signal_16011 ;
    wire new_AGEMA_signal_16015 ;
    wire new_AGEMA_signal_16016 ;
    wire new_AGEMA_signal_16017 ;
    wire new_AGEMA_signal_16021 ;
    wire new_AGEMA_signal_16022 ;
    wire new_AGEMA_signal_16023 ;
    wire new_AGEMA_signal_16027 ;
    wire new_AGEMA_signal_16028 ;
    wire new_AGEMA_signal_16029 ;
    wire new_AGEMA_signal_16030 ;
    wire new_AGEMA_signal_16031 ;
    wire new_AGEMA_signal_16032 ;
    wire new_AGEMA_signal_16033 ;
    wire new_AGEMA_signal_16034 ;
    wire new_AGEMA_signal_16035 ;
    wire new_AGEMA_signal_16036 ;
    wire new_AGEMA_signal_16037 ;
    wire new_AGEMA_signal_16038 ;
    wire new_AGEMA_signal_16039 ;
    wire new_AGEMA_signal_16040 ;
    wire new_AGEMA_signal_16041 ;
    wire new_AGEMA_signal_16042 ;
    wire new_AGEMA_signal_16043 ;
    wire new_AGEMA_signal_16044 ;
    wire new_AGEMA_signal_16045 ;
    wire new_AGEMA_signal_16046 ;
    wire new_AGEMA_signal_16047 ;
    wire new_AGEMA_signal_16048 ;
    wire new_AGEMA_signal_16049 ;
    wire new_AGEMA_signal_16050 ;
    wire new_AGEMA_signal_16051 ;
    wire new_AGEMA_signal_16052 ;
    wire new_AGEMA_signal_16053 ;
    wire new_AGEMA_signal_16054 ;
    wire new_AGEMA_signal_16055 ;
    wire new_AGEMA_signal_16056 ;
    wire new_AGEMA_signal_16057 ;
    wire new_AGEMA_signal_16058 ;
    wire new_AGEMA_signal_16059 ;
    wire new_AGEMA_signal_16060 ;
    wire new_AGEMA_signal_16061 ;
    wire new_AGEMA_signal_16062 ;
    wire new_AGEMA_signal_16063 ;
    wire new_AGEMA_signal_16064 ;
    wire new_AGEMA_signal_16065 ;
    wire new_AGEMA_signal_16066 ;
    wire new_AGEMA_signal_16067 ;
    wire new_AGEMA_signal_16068 ;
    wire new_AGEMA_signal_16069 ;
    wire new_AGEMA_signal_16070 ;
    wire new_AGEMA_signal_16071 ;
    wire new_AGEMA_signal_16072 ;
    wire new_AGEMA_signal_16073 ;
    wire new_AGEMA_signal_16074 ;
    wire new_AGEMA_signal_16075 ;
    wire new_AGEMA_signal_16076 ;
    wire new_AGEMA_signal_16077 ;
    wire new_AGEMA_signal_16078 ;
    wire new_AGEMA_signal_16079 ;
    wire new_AGEMA_signal_16080 ;
    wire new_AGEMA_signal_16081 ;
    wire new_AGEMA_signal_16082 ;
    wire new_AGEMA_signal_16083 ;
    wire new_AGEMA_signal_16084 ;
    wire new_AGEMA_signal_16085 ;
    wire new_AGEMA_signal_16086 ;
    wire new_AGEMA_signal_16087 ;
    wire new_AGEMA_signal_16088 ;
    wire new_AGEMA_signal_16089 ;
    wire new_AGEMA_signal_16090 ;
    wire new_AGEMA_signal_16091 ;
    wire new_AGEMA_signal_16092 ;
    wire new_AGEMA_signal_16093 ;
    wire new_AGEMA_signal_16094 ;
    wire new_AGEMA_signal_16095 ;
    wire new_AGEMA_signal_16096 ;
    wire new_AGEMA_signal_16097 ;
    wire new_AGEMA_signal_16098 ;
    wire new_AGEMA_signal_16099 ;
    wire new_AGEMA_signal_16100 ;
    wire new_AGEMA_signal_16101 ;
    wire new_AGEMA_signal_16102 ;
    wire new_AGEMA_signal_16103 ;
    wire new_AGEMA_signal_16104 ;
    wire new_AGEMA_signal_16105 ;
    wire new_AGEMA_signal_16106 ;
    wire new_AGEMA_signal_16107 ;
    wire new_AGEMA_signal_16108 ;
    wire new_AGEMA_signal_16109 ;
    wire new_AGEMA_signal_16110 ;
    wire new_AGEMA_signal_16111 ;
    wire new_AGEMA_signal_16112 ;
    wire new_AGEMA_signal_16113 ;
    wire new_AGEMA_signal_16114 ;
    wire new_AGEMA_signal_16115 ;
    wire new_AGEMA_signal_16116 ;
    wire new_AGEMA_signal_16117 ;
    wire new_AGEMA_signal_16118 ;
    wire new_AGEMA_signal_16119 ;
    wire new_AGEMA_signal_16120 ;
    wire new_AGEMA_signal_16121 ;
    wire new_AGEMA_signal_16122 ;
    wire new_AGEMA_signal_16123 ;
    wire new_AGEMA_signal_16124 ;
    wire new_AGEMA_signal_16125 ;
    wire new_AGEMA_signal_16126 ;
    wire new_AGEMA_signal_16127 ;
    wire new_AGEMA_signal_16128 ;
    wire new_AGEMA_signal_16129 ;
    wire new_AGEMA_signal_16130 ;
    wire new_AGEMA_signal_16131 ;
    wire new_AGEMA_signal_16132 ;
    wire new_AGEMA_signal_16133 ;
    wire new_AGEMA_signal_16134 ;
    wire new_AGEMA_signal_16135 ;
    wire new_AGEMA_signal_16136 ;
    wire new_AGEMA_signal_16137 ;
    wire new_AGEMA_signal_16138 ;
    wire new_AGEMA_signal_16139 ;
    wire new_AGEMA_signal_16140 ;
    wire new_AGEMA_signal_16141 ;
    wire new_AGEMA_signal_16142 ;
    wire new_AGEMA_signal_16143 ;
    wire new_AGEMA_signal_16144 ;
    wire new_AGEMA_signal_16145 ;
    wire new_AGEMA_signal_16146 ;
    wire new_AGEMA_signal_16147 ;
    wire new_AGEMA_signal_16148 ;
    wire new_AGEMA_signal_16149 ;
    wire new_AGEMA_signal_16150 ;
    wire new_AGEMA_signal_16151 ;
    wire new_AGEMA_signal_16152 ;
    wire new_AGEMA_signal_16153 ;
    wire new_AGEMA_signal_16154 ;
    wire new_AGEMA_signal_16155 ;
    wire new_AGEMA_signal_16156 ;
    wire new_AGEMA_signal_16157 ;
    wire new_AGEMA_signal_16158 ;
    wire new_AGEMA_signal_16159 ;
    wire new_AGEMA_signal_16160 ;
    wire new_AGEMA_signal_16161 ;
    wire new_AGEMA_signal_16162 ;
    wire new_AGEMA_signal_16163 ;
    wire new_AGEMA_signal_16164 ;
    wire new_AGEMA_signal_16165 ;
    wire new_AGEMA_signal_16166 ;
    wire new_AGEMA_signal_16167 ;
    wire new_AGEMA_signal_16168 ;
    wire new_AGEMA_signal_16169 ;
    wire new_AGEMA_signal_16170 ;
    wire new_AGEMA_signal_16171 ;
    wire new_AGEMA_signal_16172 ;
    wire new_AGEMA_signal_16173 ;
    wire new_AGEMA_signal_16174 ;
    wire new_AGEMA_signal_16175 ;
    wire new_AGEMA_signal_16176 ;
    wire new_AGEMA_signal_16177 ;
    wire new_AGEMA_signal_16178 ;
    wire new_AGEMA_signal_16179 ;
    wire new_AGEMA_signal_16180 ;
    wire new_AGEMA_signal_16181 ;
    wire new_AGEMA_signal_16182 ;
    wire new_AGEMA_signal_16183 ;
    wire new_AGEMA_signal_16184 ;
    wire new_AGEMA_signal_16185 ;
    wire new_AGEMA_signal_16186 ;
    wire new_AGEMA_signal_16187 ;
    wire new_AGEMA_signal_16188 ;
    wire new_AGEMA_signal_16189 ;
    wire new_AGEMA_signal_16190 ;
    wire new_AGEMA_signal_16191 ;
    wire new_AGEMA_signal_16192 ;
    wire new_AGEMA_signal_16193 ;
    wire new_AGEMA_signal_16194 ;
    wire new_AGEMA_signal_16198 ;
    wire new_AGEMA_signal_16199 ;
    wire new_AGEMA_signal_16200 ;
    wire new_AGEMA_signal_16204 ;
    wire new_AGEMA_signal_16205 ;
    wire new_AGEMA_signal_16206 ;
    wire new_AGEMA_signal_16210 ;
    wire new_AGEMA_signal_16211 ;
    wire new_AGEMA_signal_16212 ;
    wire new_AGEMA_signal_16216 ;
    wire new_AGEMA_signal_16217 ;
    wire new_AGEMA_signal_16218 ;
    wire new_AGEMA_signal_16222 ;
    wire new_AGEMA_signal_16223 ;
    wire new_AGEMA_signal_16224 ;
    wire new_AGEMA_signal_16228 ;
    wire new_AGEMA_signal_16229 ;
    wire new_AGEMA_signal_16230 ;
    wire new_AGEMA_signal_16234 ;
    wire new_AGEMA_signal_16235 ;
    wire new_AGEMA_signal_16236 ;
    wire new_AGEMA_signal_16240 ;
    wire new_AGEMA_signal_16241 ;
    wire new_AGEMA_signal_16242 ;
    wire new_AGEMA_signal_16246 ;
    wire new_AGEMA_signal_16247 ;
    wire new_AGEMA_signal_16248 ;
    wire new_AGEMA_signal_16252 ;
    wire new_AGEMA_signal_16253 ;
    wire new_AGEMA_signal_16254 ;
    wire new_AGEMA_signal_16258 ;
    wire new_AGEMA_signal_16259 ;
    wire new_AGEMA_signal_16260 ;
    wire new_AGEMA_signal_16264 ;
    wire new_AGEMA_signal_16265 ;
    wire new_AGEMA_signal_16266 ;
    wire new_AGEMA_signal_16270 ;
    wire new_AGEMA_signal_16271 ;
    wire new_AGEMA_signal_16272 ;
    wire new_AGEMA_signal_16276 ;
    wire new_AGEMA_signal_16277 ;
    wire new_AGEMA_signal_16278 ;
    wire new_AGEMA_signal_16282 ;
    wire new_AGEMA_signal_16283 ;
    wire new_AGEMA_signal_16284 ;
    wire new_AGEMA_signal_16288 ;
    wire new_AGEMA_signal_16289 ;
    wire new_AGEMA_signal_16290 ;
    wire new_AGEMA_signal_16294 ;
    wire new_AGEMA_signal_16295 ;
    wire new_AGEMA_signal_16296 ;
    wire new_AGEMA_signal_16300 ;
    wire new_AGEMA_signal_16301 ;
    wire new_AGEMA_signal_16302 ;
    wire new_AGEMA_signal_16306 ;
    wire new_AGEMA_signal_16307 ;
    wire new_AGEMA_signal_16308 ;
    wire new_AGEMA_signal_16312 ;
    wire new_AGEMA_signal_16313 ;
    wire new_AGEMA_signal_16314 ;
    wire new_AGEMA_signal_16318 ;
    wire new_AGEMA_signal_16319 ;
    wire new_AGEMA_signal_16320 ;
    wire new_AGEMA_signal_16324 ;
    wire new_AGEMA_signal_16325 ;
    wire new_AGEMA_signal_16326 ;
    wire new_AGEMA_signal_16330 ;
    wire new_AGEMA_signal_16331 ;
    wire new_AGEMA_signal_16332 ;
    wire new_AGEMA_signal_16336 ;
    wire new_AGEMA_signal_16337 ;
    wire new_AGEMA_signal_16338 ;
    wire new_AGEMA_signal_16342 ;
    wire new_AGEMA_signal_16343 ;
    wire new_AGEMA_signal_16344 ;
    wire new_AGEMA_signal_16348 ;
    wire new_AGEMA_signal_16349 ;
    wire new_AGEMA_signal_16350 ;
    wire new_AGEMA_signal_16354 ;
    wire new_AGEMA_signal_16355 ;
    wire new_AGEMA_signal_16356 ;
    wire new_AGEMA_signal_16360 ;
    wire new_AGEMA_signal_16361 ;
    wire new_AGEMA_signal_16362 ;
    wire new_AGEMA_signal_16366 ;
    wire new_AGEMA_signal_16367 ;
    wire new_AGEMA_signal_16368 ;
    wire new_AGEMA_signal_16372 ;
    wire new_AGEMA_signal_16373 ;
    wire new_AGEMA_signal_16374 ;
    wire new_AGEMA_signal_16378 ;
    wire new_AGEMA_signal_16379 ;
    wire new_AGEMA_signal_16380 ;
    wire new_AGEMA_signal_16384 ;
    wire new_AGEMA_signal_16385 ;
    wire new_AGEMA_signal_16386 ;
    wire new_AGEMA_signal_16390 ;
    wire new_AGEMA_signal_16391 ;
    wire new_AGEMA_signal_16392 ;
    wire new_AGEMA_signal_16396 ;
    wire new_AGEMA_signal_16397 ;
    wire new_AGEMA_signal_16398 ;
    wire new_AGEMA_signal_16402 ;
    wire new_AGEMA_signal_16403 ;
    wire new_AGEMA_signal_16404 ;
    wire new_AGEMA_signal_16408 ;
    wire new_AGEMA_signal_16409 ;
    wire new_AGEMA_signal_16410 ;
    wire new_AGEMA_signal_16414 ;
    wire new_AGEMA_signal_16415 ;
    wire new_AGEMA_signal_16416 ;
    wire new_AGEMA_signal_16420 ;
    wire new_AGEMA_signal_16421 ;
    wire new_AGEMA_signal_16422 ;
    wire new_AGEMA_signal_16426 ;
    wire new_AGEMA_signal_16427 ;
    wire new_AGEMA_signal_16428 ;
    wire new_AGEMA_signal_16432 ;
    wire new_AGEMA_signal_16433 ;
    wire new_AGEMA_signal_16434 ;
    wire new_AGEMA_signal_16438 ;
    wire new_AGEMA_signal_16439 ;
    wire new_AGEMA_signal_16440 ;
    wire new_AGEMA_signal_16444 ;
    wire new_AGEMA_signal_16445 ;
    wire new_AGEMA_signal_16446 ;
    wire new_AGEMA_signal_16450 ;
    wire new_AGEMA_signal_16451 ;
    wire new_AGEMA_signal_16452 ;
    wire new_AGEMA_signal_16456 ;
    wire new_AGEMA_signal_16457 ;
    wire new_AGEMA_signal_16458 ;
    wire new_AGEMA_signal_16462 ;
    wire new_AGEMA_signal_16463 ;
    wire new_AGEMA_signal_16464 ;
    wire new_AGEMA_signal_16468 ;
    wire new_AGEMA_signal_16469 ;
    wire new_AGEMA_signal_16470 ;
    wire new_AGEMA_signal_16474 ;
    wire new_AGEMA_signal_16475 ;
    wire new_AGEMA_signal_16476 ;
    wire new_AGEMA_signal_16480 ;
    wire new_AGEMA_signal_16481 ;
    wire new_AGEMA_signal_16482 ;
    wire new_AGEMA_signal_16486 ;
    wire new_AGEMA_signal_16487 ;
    wire new_AGEMA_signal_16488 ;
    wire new_AGEMA_signal_16492 ;
    wire new_AGEMA_signal_16493 ;
    wire new_AGEMA_signal_16494 ;
    wire new_AGEMA_signal_16498 ;
    wire new_AGEMA_signal_16499 ;
    wire new_AGEMA_signal_16500 ;
    wire new_AGEMA_signal_16504 ;
    wire new_AGEMA_signal_16505 ;
    wire new_AGEMA_signal_16506 ;
    wire new_AGEMA_signal_16510 ;
    wire new_AGEMA_signal_16511 ;
    wire new_AGEMA_signal_16512 ;
    wire new_AGEMA_signal_16516 ;
    wire new_AGEMA_signal_16517 ;
    wire new_AGEMA_signal_16518 ;
    wire new_AGEMA_signal_16522 ;
    wire new_AGEMA_signal_16523 ;
    wire new_AGEMA_signal_16524 ;
    wire new_AGEMA_signal_16528 ;
    wire new_AGEMA_signal_16529 ;
    wire new_AGEMA_signal_16530 ;
    wire new_AGEMA_signal_16534 ;
    wire new_AGEMA_signal_16535 ;
    wire new_AGEMA_signal_16536 ;
    wire new_AGEMA_signal_16540 ;
    wire new_AGEMA_signal_16541 ;
    wire new_AGEMA_signal_16542 ;
    wire new_AGEMA_signal_16546 ;
    wire new_AGEMA_signal_16547 ;
    wire new_AGEMA_signal_16548 ;
    wire new_AGEMA_signal_16552 ;
    wire new_AGEMA_signal_16553 ;
    wire new_AGEMA_signal_16554 ;
    wire new_AGEMA_signal_16558 ;
    wire new_AGEMA_signal_16559 ;
    wire new_AGEMA_signal_16560 ;
    wire new_AGEMA_signal_16564 ;
    wire new_AGEMA_signal_16565 ;
    wire new_AGEMA_signal_16566 ;
    wire new_AGEMA_signal_16570 ;
    wire new_AGEMA_signal_16571 ;
    wire new_AGEMA_signal_16572 ;
    wire new_AGEMA_signal_16576 ;
    wire new_AGEMA_signal_16577 ;
    wire new_AGEMA_signal_16578 ;
    wire new_AGEMA_signal_16582 ;
    wire new_AGEMA_signal_16583 ;
    wire new_AGEMA_signal_16584 ;
    wire new_AGEMA_signal_16588 ;
    wire new_AGEMA_signal_16589 ;
    wire new_AGEMA_signal_16590 ;
    wire new_AGEMA_signal_16594 ;
    wire new_AGEMA_signal_16595 ;
    wire new_AGEMA_signal_16596 ;
    wire new_AGEMA_signal_16600 ;
    wire new_AGEMA_signal_16601 ;
    wire new_AGEMA_signal_16602 ;
    wire new_AGEMA_signal_16606 ;
    wire new_AGEMA_signal_16607 ;
    wire new_AGEMA_signal_16608 ;
    wire new_AGEMA_signal_16612 ;
    wire new_AGEMA_signal_16613 ;
    wire new_AGEMA_signal_16614 ;
    wire new_AGEMA_signal_16618 ;
    wire new_AGEMA_signal_16619 ;
    wire new_AGEMA_signal_16620 ;
    wire new_AGEMA_signal_16624 ;
    wire new_AGEMA_signal_16625 ;
    wire new_AGEMA_signal_16626 ;
    wire new_AGEMA_signal_16630 ;
    wire new_AGEMA_signal_16631 ;
    wire new_AGEMA_signal_16632 ;
    wire new_AGEMA_signal_16636 ;
    wire new_AGEMA_signal_16637 ;
    wire new_AGEMA_signal_16638 ;
    wire new_AGEMA_signal_16642 ;
    wire new_AGEMA_signal_16643 ;
    wire new_AGEMA_signal_16644 ;
    wire new_AGEMA_signal_16648 ;
    wire new_AGEMA_signal_16649 ;
    wire new_AGEMA_signal_16650 ;
    wire new_AGEMA_signal_16654 ;
    wire new_AGEMA_signal_16655 ;
    wire new_AGEMA_signal_16656 ;
    wire new_AGEMA_signal_16660 ;
    wire new_AGEMA_signal_16661 ;
    wire new_AGEMA_signal_16662 ;
    wire new_AGEMA_signal_16666 ;
    wire new_AGEMA_signal_16667 ;
    wire new_AGEMA_signal_16668 ;
    wire new_AGEMA_signal_16672 ;
    wire new_AGEMA_signal_16673 ;
    wire new_AGEMA_signal_16674 ;
    wire new_AGEMA_signal_16678 ;
    wire new_AGEMA_signal_16679 ;
    wire new_AGEMA_signal_16680 ;
    wire new_AGEMA_signal_16684 ;
    wire new_AGEMA_signal_16685 ;
    wire new_AGEMA_signal_16686 ;
    wire new_AGEMA_signal_16690 ;
    wire new_AGEMA_signal_16691 ;
    wire new_AGEMA_signal_16692 ;
    wire new_AGEMA_signal_16696 ;
    wire new_AGEMA_signal_16697 ;
    wire new_AGEMA_signal_16698 ;
    wire new_AGEMA_signal_16702 ;
    wire new_AGEMA_signal_16703 ;
    wire new_AGEMA_signal_16704 ;
    wire new_AGEMA_signal_16708 ;
    wire new_AGEMA_signal_16709 ;
    wire new_AGEMA_signal_16710 ;
    wire new_AGEMA_signal_16714 ;
    wire new_AGEMA_signal_16715 ;
    wire new_AGEMA_signal_16716 ;
    wire new_AGEMA_signal_16720 ;
    wire new_AGEMA_signal_16721 ;
    wire new_AGEMA_signal_16722 ;
    wire new_AGEMA_signal_16726 ;
    wire new_AGEMA_signal_16727 ;
    wire new_AGEMA_signal_16728 ;
    wire new_AGEMA_signal_16732 ;
    wire new_AGEMA_signal_16733 ;
    wire new_AGEMA_signal_16734 ;
    wire new_AGEMA_signal_16738 ;
    wire new_AGEMA_signal_16739 ;
    wire new_AGEMA_signal_16740 ;
    wire new_AGEMA_signal_16744 ;
    wire new_AGEMA_signal_16745 ;
    wire new_AGEMA_signal_16746 ;
    wire new_AGEMA_signal_16750 ;
    wire new_AGEMA_signal_16751 ;
    wire new_AGEMA_signal_16752 ;
    wire new_AGEMA_signal_16756 ;
    wire new_AGEMA_signal_16757 ;
    wire new_AGEMA_signal_16758 ;
    wire new_AGEMA_signal_16762 ;
    wire new_AGEMA_signal_16763 ;
    wire new_AGEMA_signal_16764 ;
    wire new_AGEMA_signal_16768 ;
    wire new_AGEMA_signal_16769 ;
    wire new_AGEMA_signal_16770 ;
    wire new_AGEMA_signal_16774 ;
    wire new_AGEMA_signal_16775 ;
    wire new_AGEMA_signal_16776 ;
    wire new_AGEMA_signal_16780 ;
    wire new_AGEMA_signal_16781 ;
    wire new_AGEMA_signal_16782 ;
    wire new_AGEMA_signal_16786 ;
    wire new_AGEMA_signal_16787 ;
    wire new_AGEMA_signal_16788 ;
    wire new_AGEMA_signal_16792 ;
    wire new_AGEMA_signal_16793 ;
    wire new_AGEMA_signal_16794 ;
    wire new_AGEMA_signal_16798 ;
    wire new_AGEMA_signal_16799 ;
    wire new_AGEMA_signal_16800 ;
    wire new_AGEMA_signal_16804 ;
    wire new_AGEMA_signal_16805 ;
    wire new_AGEMA_signal_16806 ;
    wire new_AGEMA_signal_16810 ;
    wire new_AGEMA_signal_16811 ;
    wire new_AGEMA_signal_16812 ;
    wire new_AGEMA_signal_16816 ;
    wire new_AGEMA_signal_16817 ;
    wire new_AGEMA_signal_16818 ;
    wire new_AGEMA_signal_16822 ;
    wire new_AGEMA_signal_16823 ;
    wire new_AGEMA_signal_16824 ;
    wire new_AGEMA_signal_16828 ;
    wire new_AGEMA_signal_16829 ;
    wire new_AGEMA_signal_16830 ;
    wire new_AGEMA_signal_16834 ;
    wire new_AGEMA_signal_16835 ;
    wire new_AGEMA_signal_16836 ;
    wire new_AGEMA_signal_16840 ;
    wire new_AGEMA_signal_16841 ;
    wire new_AGEMA_signal_16842 ;
    wire new_AGEMA_signal_16846 ;
    wire new_AGEMA_signal_16847 ;
    wire new_AGEMA_signal_16848 ;
    wire new_AGEMA_signal_16852 ;
    wire new_AGEMA_signal_16853 ;
    wire new_AGEMA_signal_16854 ;
    wire new_AGEMA_signal_16858 ;
    wire new_AGEMA_signal_16859 ;
    wire new_AGEMA_signal_16860 ;
    wire new_AGEMA_signal_16864 ;
    wire new_AGEMA_signal_16865 ;
    wire new_AGEMA_signal_16866 ;
    wire new_AGEMA_signal_16870 ;
    wire new_AGEMA_signal_16871 ;
    wire new_AGEMA_signal_16872 ;
    wire new_AGEMA_signal_16876 ;
    wire new_AGEMA_signal_16877 ;
    wire new_AGEMA_signal_16878 ;
    wire new_AGEMA_signal_16882 ;
    wire new_AGEMA_signal_16883 ;
    wire new_AGEMA_signal_16884 ;
    wire new_AGEMA_signal_16888 ;
    wire new_AGEMA_signal_16889 ;
    wire new_AGEMA_signal_16890 ;
    wire new_AGEMA_signal_16894 ;
    wire new_AGEMA_signal_16895 ;
    wire new_AGEMA_signal_16896 ;
    wire new_AGEMA_signal_16900 ;
    wire new_AGEMA_signal_16901 ;
    wire new_AGEMA_signal_16902 ;
    wire new_AGEMA_signal_16906 ;
    wire new_AGEMA_signal_16907 ;
    wire new_AGEMA_signal_16908 ;
    wire new_AGEMA_signal_16912 ;
    wire new_AGEMA_signal_16913 ;
    wire new_AGEMA_signal_16914 ;
    wire new_AGEMA_signal_16918 ;
    wire new_AGEMA_signal_16919 ;
    wire new_AGEMA_signal_16920 ;
    wire new_AGEMA_signal_16924 ;
    wire new_AGEMA_signal_16925 ;
    wire new_AGEMA_signal_16926 ;
    wire new_AGEMA_signal_16930 ;
    wire new_AGEMA_signal_16931 ;
    wire new_AGEMA_signal_16932 ;
    wire new_AGEMA_signal_16936 ;
    wire new_AGEMA_signal_16937 ;
    wire new_AGEMA_signal_16938 ;
    wire new_AGEMA_signal_16942 ;
    wire new_AGEMA_signal_16943 ;
    wire new_AGEMA_signal_16944 ;
    wire new_AGEMA_signal_16948 ;
    wire new_AGEMA_signal_16949 ;
    wire new_AGEMA_signal_16950 ;
    wire new_AGEMA_signal_16954 ;
    wire new_AGEMA_signal_16955 ;
    wire new_AGEMA_signal_16956 ;
    wire new_AGEMA_signal_16960 ;
    wire new_AGEMA_signal_16961 ;
    wire new_AGEMA_signal_16962 ;
    wire new_AGEMA_signal_16966 ;
    wire new_AGEMA_signal_16967 ;
    wire new_AGEMA_signal_16968 ;
    wire new_AGEMA_signal_16972 ;
    wire new_AGEMA_signal_16973 ;
    wire new_AGEMA_signal_16974 ;
    wire new_AGEMA_signal_16978 ;
    wire new_AGEMA_signal_16979 ;
    wire new_AGEMA_signal_16980 ;
    wire new_AGEMA_signal_16984 ;
    wire new_AGEMA_signal_16985 ;
    wire new_AGEMA_signal_16986 ;
    wire new_AGEMA_signal_16990 ;
    wire new_AGEMA_signal_16991 ;
    wire new_AGEMA_signal_16992 ;
    wire new_AGEMA_signal_16996 ;
    wire new_AGEMA_signal_16997 ;
    wire new_AGEMA_signal_16998 ;
    wire new_AGEMA_signal_17002 ;
    wire new_AGEMA_signal_17003 ;
    wire new_AGEMA_signal_17004 ;
    wire clk_gated ;

    /* cells in depth 0 */
    INV_X1 U830 ( .A (n314), .ZN (n319) ) ;
    INV_X1 U831 ( .A (n314), .ZN (n320) ) ;
    INV_X1 U832 ( .A (n314), .ZN (n317) ) ;
    INV_X1 U833 ( .A (n314), .ZN (n315) ) ;
    INV_X1 U834 ( .A (n314), .ZN (n316) ) ;
    INV_X1 U835 ( .A (n314), .ZN (n318) ) ;
    NOR2_X1 U836 ( .A1 (n325), .A2 (n330), .ZN (n314) ) ;
    INV_X1 U837 ( .A (RoundCounter[0]), .ZN (n325) ) ;
    INV_X1 U838 ( .A (n314), .ZN (n321) ) ;
    NOR2_X1 U839 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n323) ) ;
    INV_X1 U840 ( .A (n323), .ZN (n322) ) ;
    NOR2_X1 U841 ( .A1 (RoundCounter[0]), .A2 (n322), .ZN (Rcon[0]) ) ;
    NOR2_X1 U842 ( .A1 (RoundCounter[0]), .A2 (RoundCounter[3]), .ZN (n337) ) ;
    NOR2_X1 U843 ( .A1 (n337), .A2 (n322), .ZN (Rcon[1]) ) ;
    NAND2_X1 U844 ( .A1 (RoundCounter[3]), .A2 (n323), .ZN (n330) ) ;
    INV_X1 U845 ( .A (RoundCounter[2]), .ZN (n328) ) ;
    AND2_X1 U846 ( .A1 (n328), .A2 (RoundCounter[1]), .ZN (n333) ) ;
    NAND2_X1 U847 ( .A1 (n337), .A2 (n333), .ZN (n324) ) ;
    NAND2_X1 U848 ( .A1 (n321), .A2 (n324), .ZN (Rcon[2]) ) ;
    NOR2_X1 U849 ( .A1 (RoundCounter[3]), .A2 (n325), .ZN (n335) ) ;
    NAND2_X1 U850 ( .A1 (n333), .A2 (n335), .ZN (n327) ) ;
    NAND2_X1 U851 ( .A1 (RoundCounter[3]), .A2 (Rcon[0]), .ZN (n326) ) ;
    NAND2_X1 U852 ( .A1 (n327), .A2 (n326), .ZN (Rcon[3]) ) ;
    NOR2_X1 U853 ( .A1 (RoundCounter[1]), .A2 (n328), .ZN (n331) ) ;
    NAND2_X1 U854 ( .A1 (n337), .A2 (n331), .ZN (n329) ) ;
    NAND2_X1 U855 ( .A1 (n330), .A2 (n329), .ZN (Rcon[4]) ) ;
    NAND2_X1 U856 ( .A1 (n335), .A2 (n331), .ZN (n332) ) ;
    NAND2_X1 U857 ( .A1 (n321), .A2 (n332), .ZN (Rcon[5]) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U986 ( .a ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .c ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U987 ( .a ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, RoundInput[100]}), .b ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundKey[100]}), .c ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U988 ( .a ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[101]}), .b ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, RoundKey[101]}), .c ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U989 ( .a ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, RoundInput[102]}), .b ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundKey[102]}), .c ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U990 ( .a ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[103]}), .b ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, RoundKey[103]}), .c ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U991 ( .a ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, RoundInput[104]}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundKey[104]}), .c ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U992 ( .a ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[105]}), .b ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, RoundKey[105]}), .c ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U993 ( .a ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, RoundInput[106]}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundKey[106]}), .c ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U994 ( .a ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[107]}), .b ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, RoundKey[107]}), .c ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U995 ( .a ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, RoundInput[108]}), .b ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundKey[108]}), .c ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U996 ( .a ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[109]}), .b ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, RoundKey[109]}), .c ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U997 ( .a ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, RoundInput[10]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U998 ( .a ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[110]}), .b ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, RoundKey[110]}), .c ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U999 ( .a ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, RoundInput[111]}), .b ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundKey[111]}), .c ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1000 ( .a ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[112]}), .b ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, RoundKey[112]}), .c ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1001 ( .a ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, RoundInput[113]}), .b ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundKey[113]}), .c ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1002 ( .a ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[114]}), .b ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, RoundKey[114]}), .c ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1003 ( .a ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, RoundInput[115]}), .b ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundKey[115]}), .c ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1004 ( .a ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[116]}), .b ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, RoundKey[116]}), .c ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1005 ( .a ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, RoundInput[117]}), .b ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundKey[117]}), .c ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1006 ( .a ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[118]}), .b ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, RoundKey[118]}), .c ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1007 ( .a ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, RoundInput[119]}), .b ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundKey[119]}), .c ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1008 ( .a ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[11]}), .b ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}), .c ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1009 ( .a ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, RoundInput[120]}), .b ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundKey[120]}), .c ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1010 ( .a ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[121]}), .b ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, RoundKey[121]}), .c ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1011 ( .a ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, RoundInput[122]}), .b ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundKey[122]}), .c ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1012 ( .a ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[123]}), .b ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, RoundKey[123]}), .c ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1013 ( .a ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, RoundInput[124]}), .b ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundKey[124]}), .c ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1014 ( .a ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[125]}), .b ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, RoundKey[125]}), .c ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1015 ( .a ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, RoundInput[126]}), .b ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundKey[126]}), .c ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1016 ( .a ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[127]}), .b ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, RoundKey[127]}), .c ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1017 ( .a ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, RoundInput[12]}), .b ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .c ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1018 ( .a ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[13]}), .b ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .c ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1019 ( .a ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, RoundInput[14]}), .b ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .c ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1020 ( .a ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[15]}), .b ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .c ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1021 ( .a ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, RoundInput[16]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .c ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1022 ( .a ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[17]}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .c ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1023 ( .a ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, RoundInput[18]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1024 ( .a ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[19]}), .b ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}), .c ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1025 ( .a ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, RoundInput[1]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .c ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1026 ( .a ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[20]}), .b ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .c ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1027 ( .a ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, RoundInput[21]}), .b ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .c ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1028 ( .a ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[22]}), .b ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .c ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1029 ( .a ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, RoundInput[23]}), .b ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .c ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1030 ( .a ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[24]}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .c ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1031 ( .a ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, RoundInput[25]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .c ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1032 ( .a ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[26]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1033 ( .a ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, RoundInput[27]}), .b ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}), .c ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1034 ( .a ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[28]}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .c ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1035 ( .a ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, RoundInput[29]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .c ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1036 ( .a ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[2]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1037 ( .a ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, RoundInput[30]}), .b ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .c ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1038 ( .a ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[31]}), .b ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .c ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1039 ( .a ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, RoundInput[32]}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundKey[32]}), .c ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1040 ( .a ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[33]}), .b ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, RoundKey[33]}), .c ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1041 ( .a ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, RoundInput[34]}), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundKey[34]}), .c ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1042 ( .a ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[35]}), .b ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKey[35]}), .c ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1043 ( .a ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundInput[36]}), .b ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundKey[36]}), .c ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1044 ( .a ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[37]}), .b ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKey[37]}), .c ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1045 ( .a ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundInput[38]}), .b ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundKey[38]}), .c ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1046 ( .a ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[39]}), .b ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKey[39]}), .c ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1047 ( .a ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundInput[3]}), .b ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}), .c ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1048 ( .a ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[40]}), .b ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, RoundKey[40]}), .c ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1049 ( .a ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, RoundInput[41]}), .b ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundKey[41]}), .c ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1050 ( .a ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[42]}), .b ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, RoundKey[42]}), .c ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1051 ( .a ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, RoundInput[43]}), .b ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundKey[43]}), .c ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1052 ( .a ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[44]}), .b ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, RoundKey[44]}), .c ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1053 ( .a ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, RoundInput[45]}), .b ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundKey[45]}), .c ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1054 ( .a ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[46]}), .b ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, RoundKey[46]}), .c ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1055 ( .a ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, RoundInput[47]}), .b ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundKey[47]}), .c ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1056 ( .a ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[48]}), .b ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, RoundKey[48]}), .c ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1057 ( .a ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, RoundInput[49]}), .b ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundKey[49]}), .c ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1058 ( .a ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[4]}), .b ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .c ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1059 ( .a ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, RoundInput[50]}), .b ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundKey[50]}), .c ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1060 ( .a ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[51]}), .b ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, RoundKey[51]}), .c ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1061 ( .a ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, RoundInput[52]}), .b ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundKey[52]}), .c ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1062 ( .a ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[53]}), .b ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, RoundKey[53]}), .c ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1063 ( .a ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, RoundInput[54]}), .b ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundKey[54]}), .c ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1064 ( .a ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[55]}), .b ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, RoundKey[55]}), .c ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1065 ( .a ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, RoundInput[56]}), .b ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundKey[56]}), .c ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1066 ( .a ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[57]}), .b ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, RoundKey[57]}), .c ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1067 ( .a ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, RoundInput[58]}), .b ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundKey[58]}), .c ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1068 ( .a ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[59]}), .b ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, RoundKey[59]}), .c ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1069 ( .a ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, RoundInput[5]}), .b ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .c ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1070 ( .a ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[60]}), .b ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, RoundKey[60]}), .c ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1071 ( .a ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, RoundInput[61]}), .b ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, RoundKey[61]}), .c ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1072 ( .a ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, new_AGEMA_signal_5323, RoundInput[62]}), .b ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, RoundKey[62]}), .c ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1073 ( .a ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundInput[63]}), .b ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, RoundKey[63]}), .c ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1074 ( .a ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, RoundInput[64]}), .b ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKey[64]}), .c ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1075 ( .a ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundInput[65]}), .b ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, RoundKey[65]}), .c ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1076 ( .a ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, new_AGEMA_signal_5359, RoundInput[66]}), .b ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKey[66]}), .c ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1077 ( .a ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundInput[67]}), .b ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, RoundKey[67]}), .c ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1078 ( .a ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, RoundInput[68]}), .b ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKey[68]}), .c ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1079 ( .a ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundInput[69]}), .b ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, RoundKey[69]}), .c ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1080 ( .a ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, new_AGEMA_signal_5395, RoundInput[6]}), .b ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .c ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1081 ( .a ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, new_AGEMA_signal_5404, RoundInput[70]}), .b ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, RoundKey[70]}), .c ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1082 ( .a ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, RoundInput[71]}), .b ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, RoundKey[71]}), .c ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1083 ( .a ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, new_AGEMA_signal_5422, RoundInput[72]}), .b ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, RoundKey[72]}), .c ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1084 ( .a ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, new_AGEMA_signal_5431, RoundInput[73]}), .b ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, RoundKey[73]}), .c ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1085 ( .a ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, new_AGEMA_signal_5440, RoundInput[74]}), .b ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, RoundKey[74]}), .c ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1086 ( .a ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, RoundInput[75]}), .b ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, RoundKey[75]}), .c ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1087 ( .a ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, new_AGEMA_signal_5458, RoundInput[76]}), .b ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, RoundKey[76]}), .c ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1088 ( .a ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, new_AGEMA_signal_5467, RoundInput[77]}), .b ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, RoundKey[77]}), .c ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1089 ( .a ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, new_AGEMA_signal_5476, RoundInput[78]}), .b ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, RoundKey[78]}), .c ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1090 ( .a ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, RoundInput[79]}), .b ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, RoundKey[79]}), .c ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1091 ( .a ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, new_AGEMA_signal_5494, RoundInput[7]}), .b ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .c ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1092 ( .a ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, new_AGEMA_signal_5503, RoundInput[80]}), .b ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, RoundKey[80]}), .c ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1093 ( .a ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, new_AGEMA_signal_5512, RoundInput[81]}), .b ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, RoundKey[81]}), .c ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1094 ( .a ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, RoundInput[82]}), .b ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, RoundKey[82]}), .c ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1095 ( .a ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, new_AGEMA_signal_5530, RoundInput[83]}), .b ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, RoundKey[83]}), .c ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1096 ( .a ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5539, RoundInput[84]}), .b ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, RoundKey[84]}), .c ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1097 ( .a ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, RoundInput[85]}), .b ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, RoundKey[85]}), .c ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1098 ( .a ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5557, RoundInput[86]}), .b ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, RoundKey[86]}), .c ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1099 ( .a ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, new_AGEMA_signal_5566, RoundInput[87]}), .b ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, RoundKey[87]}), .c ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1100 ( .a ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, RoundInput[88]}), .b ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, RoundKey[88]}), .c ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1101 ( .a ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, RoundInput[89]}), .b ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, RoundKey[89]}), .c ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1102 ( .a ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, new_AGEMA_signal_5593, RoundInput[8]}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .c ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1103 ( .a ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, RoundInput[90]}), .b ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, RoundKey[90]}), .c ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1104 ( .a ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, RoundInput[91]}), .b ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, RoundKey[91]}), .c ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1105 ( .a ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, new_AGEMA_signal_5620, RoundInput[92]}), .b ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, RoundKey[92]}), .c ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1106 ( .a ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, new_AGEMA_signal_5629, RoundInput[93]}), .b ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, RoundKey[93]}), .c ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1107 ( .a ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, RoundInput[94]}), .b ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, RoundKey[94]}), .c ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1108 ( .a ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, new_AGEMA_signal_5647, RoundInput[95]}), .b ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKey[95]}), .c ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1109 ( .a ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundInput[96]}), .b ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, RoundKey[96]}), .c ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1110 ( .a ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, RoundInput[97]}), .b ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKey[97]}), .c ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1111 ( .a ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundInput[98]}), .b ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, RoundKey[98]}), .c ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1112 ( .a ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, new_AGEMA_signal_5683, RoundInput[99]}), .b ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKey[99]}), .c ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) U1113 ( .a ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundInput[9]}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .c ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    NAND2_X1 U1114 ( .A1 (RoundCounter[3]), .A2 (n333), .ZN (n334) ) ;
    NOR2_X1 U1115 ( .A1 (RoundCounter[0]), .A2 (n334), .ZN (done) ) ;
    INV_X1 U1116 ( .A (n335), .ZN (n336) ) ;
    NAND2_X1 U1117 ( .A1 (RoundCounter[2]), .A2 (RoundCounter[1]), .ZN (n338) ) ;
    NOR2_X1 U1118 ( .A1 (n336), .A2 (n338), .ZN (n283) ) ;
    INV_X1 U1119 ( .A (n337), .ZN (n339) ) ;
    NOR2_X1 U1120 ( .A1 (n339), .A2 (n338), .ZN (n285) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T1_U1 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T2_U1 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T3_U1 ( .a ({ciphertext_s3[7], ciphertext_s2[7], ciphertext_s1[7], ciphertext_s0[7]}), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T4_U1 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T5_U1 ( .a ({ciphertext_s3[3], ciphertext_s2[3], ciphertext_s1[3], ciphertext_s0[3]}), .b ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T7_U1 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T8_U1 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T9_U1 ( .a ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T11_U1 ( .a ({ciphertext_s3[6], ciphertext_s2[6], ciphertext_s1[6], ciphertext_s0[6]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T12_U1 ( .a ({ciphertext_s3[5], ciphertext_s2[5], ciphertext_s1[5], ciphertext_s0[5]}), .b ({ciphertext_s3[2], ciphertext_s2[2], ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5841, new_AGEMA_signal_5840, new_AGEMA_signal_5839, SubBytesIns_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5835, new_AGEMA_signal_5834, new_AGEMA_signal_5833, SubBytesIns_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T18_U1 ( .a ({ciphertext_s3[4], ciphertext_s2[4], ciphertext_s1[4], ciphertext_s0[4]}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5847, new_AGEMA_signal_5846, new_AGEMA_signal_5845, SubBytesIns_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T21_U1 ( .a ({ciphertext_s3[1], ciphertext_s2[1], ciphertext_s1[1], ciphertext_s0[1]}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, new_AGEMA_signal_5848, SubBytesIns_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5838, new_AGEMA_signal_5837, new_AGEMA_signal_5836, SubBytesIns_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5850, new_AGEMA_signal_5849, new_AGEMA_signal_5848, SubBytesIns_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_7671, new_AGEMA_signal_7670, new_AGEMA_signal_7669, SubBytesIns_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, new_AGEMA_signal_7672, SubBytesIns_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, new_AGEMA_signal_6955, SubBytesIns_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5844, new_AGEMA_signal_5843, new_AGEMA_signal_5842, SubBytesIns_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T1_U1 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T2_U1 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T3_U1 ( .a ({ciphertext_s3[15], ciphertext_s2[15], ciphertext_s1[15], ciphertext_s0[15]}), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T4_U1 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T5_U1 ( .a ({ciphertext_s3[11], ciphertext_s2[11], ciphertext_s1[11], ciphertext_s0[11]}), .b ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T7_U1 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T8_U1 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, SubBytesIns_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T9_U1 ( .a ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T11_U1 ( .a ({ciphertext_s3[14], ciphertext_s2[14], ciphertext_s1[14], ciphertext_s0[14]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T12_U1 ( .a ({ciphertext_s3[13], ciphertext_s2[13], ciphertext_s1[13], ciphertext_s0[13]}), .b ({ciphertext_s3[10], ciphertext_s2[10], ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, new_AGEMA_signal_6982, SubBytesIns_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5871, new_AGEMA_signal_5870, new_AGEMA_signal_5869, SubBytesIns_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5865, new_AGEMA_signal_5864, new_AGEMA_signal_5863, SubBytesIns_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T18_U1 ( .a ({ciphertext_s3[12], ciphertext_s2[12], ciphertext_s1[12], ciphertext_s0[12]}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5877, new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5877, new_AGEMA_signal_5876, new_AGEMA_signal_5875, SubBytesIns_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T21_U1 ( .a ({ciphertext_s3[9], ciphertext_s2[9], ciphertext_s1[9], ciphertext_s0[9]}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5868, new_AGEMA_signal_5867, new_AGEMA_signal_5866, SubBytesIns_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5880, new_AGEMA_signal_5879, new_AGEMA_signal_5878, SubBytesIns_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, new_AGEMA_signal_7696, SubBytesIns_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5874, new_AGEMA_signal_5873, new_AGEMA_signal_5872, SubBytesIns_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T1_U1 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T2_U1 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T3_U1 ( .a ({ciphertext_s3[23], ciphertext_s2[23], ciphertext_s1[23], ciphertext_s0[23]}), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T4_U1 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T5_U1 ( .a ({ciphertext_s3[19], ciphertext_s2[19], ciphertext_s1[19], ciphertext_s0[19]}), .b ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T7_U1 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T8_U1 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T9_U1 ( .a ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .b ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T11_U1 ( .a ({ciphertext_s3[22], ciphertext_s2[22], ciphertext_s1[22], ciphertext_s0[22]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T12_U1 ( .a ({ciphertext_s3[21], ciphertext_s2[21], ciphertext_s1[21], ciphertext_s0[21]}), .b ({ciphertext_s3[18], ciphertext_s2[18], ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5901, new_AGEMA_signal_5900, new_AGEMA_signal_5899, SubBytesIns_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5895, new_AGEMA_signal_5894, new_AGEMA_signal_5893, SubBytesIns_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T18_U1 ( .a ({ciphertext_s3[20], ciphertext_s2[20], ciphertext_s1[20], ciphertext_s0[20]}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5907, new_AGEMA_signal_5906, new_AGEMA_signal_5905, SubBytesIns_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T21_U1 ( .a ({ciphertext_s3[17], ciphertext_s2[17], ciphertext_s1[17], ciphertext_s0[17]}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5898, new_AGEMA_signal_5897, new_AGEMA_signal_5896, SubBytesIns_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5910, new_AGEMA_signal_5909, new_AGEMA_signal_5908, SubBytesIns_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, new_AGEMA_signal_7726, SubBytesIns_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5904, new_AGEMA_signal_5903, new_AGEMA_signal_5902, SubBytesIns_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T1_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T2_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T3_U1 ( .a ({ciphertext_s3[31], ciphertext_s2[31], ciphertext_s1[31], ciphertext_s0[31]}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T4_U1 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T5_U1 ( .a ({ciphertext_s3[27], ciphertext_s2[27], ciphertext_s1[27], ciphertext_s0[27]}), .b ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T7_U1 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T8_U1 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T9_U1 ( .a ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T11_U1 ( .a ({ciphertext_s3[30], ciphertext_s2[30], ciphertext_s1[30], ciphertext_s0[30]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T12_U1 ( .a ({ciphertext_s3[29], ciphertext_s2[29], ciphertext_s1[29], ciphertext_s0[29]}), .b ({ciphertext_s3[26], ciphertext_s2[26], ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5931, new_AGEMA_signal_5930, new_AGEMA_signal_5929, SubBytesIns_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5925, new_AGEMA_signal_5924, new_AGEMA_signal_5923, SubBytesIns_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T18_U1 ( .a ({ciphertext_s3[28], ciphertext_s2[28], ciphertext_s1[28], ciphertext_s0[28]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5937, new_AGEMA_signal_5936, new_AGEMA_signal_5935, SubBytesIns_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T21_U1 ( .a ({ciphertext_s3[25], ciphertext_s2[25], ciphertext_s1[25], ciphertext_s0[25]}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5928, new_AGEMA_signal_5927, new_AGEMA_signal_5926, SubBytesIns_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5940, new_AGEMA_signal_5939, new_AGEMA_signal_5938, SubBytesIns_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, new_AGEMA_signal_7750, SubBytesIns_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5934, new_AGEMA_signal_5933, new_AGEMA_signal_5932, SubBytesIns_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_3_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T1_U1 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T2_U1 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T3_U1 ( .a ({ciphertext_s3[39], ciphertext_s2[39], ciphertext_s1[39], ciphertext_s0[39]}), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T4_U1 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T5_U1 ( .a ({ciphertext_s3[35], ciphertext_s2[35], ciphertext_s1[35], ciphertext_s0[35]}), .b ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T6_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}), .c ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T7_U1 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T8_U1 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .c ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_4_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T9_U1 ( .a ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T10_U1 ( .a ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .c ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T11_U1 ( .a ({ciphertext_s3[38], ciphertext_s2[38], ciphertext_s1[38], ciphertext_s0[38]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_4_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T12_U1 ( .a ({ciphertext_s3[37], ciphertext_s2[37], ciphertext_s1[37], ciphertext_s0[37]}), .b ({ciphertext_s3[34], ciphertext_s2[34], ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_4_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T13_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}), .c ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_4_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T14_U1 ( .a ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_4_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T15_U1 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5961, new_AGEMA_signal_5960, new_AGEMA_signal_5959, SubBytesIns_Inst_Sbox_4_T11}), .c ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_4_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T16_U1 ( .a ({new_AGEMA_signal_5955, new_AGEMA_signal_5954, new_AGEMA_signal_5953, SubBytesIns_Inst_Sbox_4_T5}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T17_U1 ( .a ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T18_U1 ( .a ({ciphertext_s3[36], ciphertext_s2[36], ciphertext_s1[36], ciphertext_s0[36]}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_4_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T19_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5967, new_AGEMA_signal_5966, new_AGEMA_signal_5965, SubBytesIns_Inst_Sbox_4_T18}), .c ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T20_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}), .c ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T21_U1 ( .a ({ciphertext_s3[33], ciphertext_s2[33], ciphertext_s1[33], ciphertext_s0[33]}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_4_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T22_U1 ( .a ({new_AGEMA_signal_5958, new_AGEMA_signal_5957, new_AGEMA_signal_5956, SubBytesIns_Inst_Sbox_4_T7}), .b ({new_AGEMA_signal_5970, new_AGEMA_signal_5969, new_AGEMA_signal_5968, SubBytesIns_Inst_Sbox_4_T21}), .c ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T23_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}), .c ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_4_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T24_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}), .c ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_4_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T25_U1 ( .a ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}), .c ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, new_AGEMA_signal_7780, SubBytesIns_Inst_Sbox_4_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T26_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .c ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_4_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_T27_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_5964, new_AGEMA_signal_5963, new_AGEMA_signal_5962, SubBytesIns_Inst_Sbox_4_T12}), .c ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, SubBytesIns_Inst_Sbox_4_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T1_U1 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T2_U1 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T3_U1 ( .a ({ciphertext_s3[47], ciphertext_s2[47], ciphertext_s1[47], ciphertext_s0[47]}), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T4_U1 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T5_U1 ( .a ({ciphertext_s3[43], ciphertext_s2[43], ciphertext_s1[43], ciphertext_s0[43]}), .b ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T6_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}), .c ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T7_U1 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T8_U1 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .c ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_5_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T9_U1 ( .a ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T10_U1 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .c ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T11_U1 ( .a ({ciphertext_s3[46], ciphertext_s2[46], ciphertext_s1[46], ciphertext_s0[46]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_5_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T12_U1 ( .a ({ciphertext_s3[45], ciphertext_s2[45], ciphertext_s1[45], ciphertext_s0[45]}), .b ({ciphertext_s3[42], ciphertext_s2[42], ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_5_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T13_U1 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}), .c ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_5_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T14_U1 ( .a ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .b ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, new_AGEMA_signal_7138, SubBytesIns_Inst_Sbox_5_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T15_U1 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5991, new_AGEMA_signal_5990, new_AGEMA_signal_5989, SubBytesIns_Inst_Sbox_5_T11}), .c ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, SubBytesIns_Inst_Sbox_5_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T16_U1 ( .a ({new_AGEMA_signal_5985, new_AGEMA_signal_5984, new_AGEMA_signal_5983, SubBytesIns_Inst_Sbox_5_T5}), .b ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T17_U1 ( .a ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T18_U1 ( .a ({ciphertext_s3[44], ciphertext_s2[44], ciphertext_s1[44], ciphertext_s0[44]}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_5997, new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_5_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T19_U1 ( .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_5997, new_AGEMA_signal_5996, new_AGEMA_signal_5995, SubBytesIns_Inst_Sbox_5_T18}), .c ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T20_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}), .c ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T21_U1 ( .a ({ciphertext_s3[41], ciphertext_s2[41], ciphertext_s1[41], ciphertext_s0[41]}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, SubBytesIns_Inst_Sbox_5_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T22_U1 ( .a ({new_AGEMA_signal_5988, new_AGEMA_signal_5987, new_AGEMA_signal_5986, SubBytesIns_Inst_Sbox_5_T7}), .b ({new_AGEMA_signal_6000, new_AGEMA_signal_5999, new_AGEMA_signal_5998, SubBytesIns_Inst_Sbox_5_T21}), .c ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T23_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}), .c ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, SubBytesIns_Inst_Sbox_5_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T24_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}), .c ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, new_AGEMA_signal_7804, SubBytesIns_Inst_Sbox_5_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T25_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}), .c ({new_AGEMA_signal_7809, new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_5_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T26_U1 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .c ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, new_AGEMA_signal_7150, SubBytesIns_Inst_Sbox_5_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_T27_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_5994, new_AGEMA_signal_5993, new_AGEMA_signal_5992, SubBytesIns_Inst_Sbox_5_T12}), .c ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, SubBytesIns_Inst_Sbox_5_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T1_U1 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T2_U1 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T3_U1 ( .a ({ciphertext_s3[55], ciphertext_s2[55], ciphertext_s1[55], ciphertext_s0[55]}), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T4_U1 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T5_U1 ( .a ({ciphertext_s3[51], ciphertext_s2[51], ciphertext_s1[51], ciphertext_s0[51]}), .b ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T6_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}), .c ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T7_U1 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T8_U1 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .c ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_6_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T9_U1 ( .a ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T10_U1 ( .a ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .c ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T11_U1 ( .a ({ciphertext_s3[54], ciphertext_s2[54], ciphertext_s1[54], ciphertext_s0[54]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_6_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T12_U1 ( .a ({ciphertext_s3[53], ciphertext_s2[53], ciphertext_s1[53], ciphertext_s0[53]}), .b ({ciphertext_s3[50], ciphertext_s2[50], ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_6_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T13_U1 ( .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}), .c ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_6_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T14_U1 ( .a ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .b ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_6_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T15_U1 ( .a ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_6021, new_AGEMA_signal_6020, new_AGEMA_signal_6019, SubBytesIns_Inst_Sbox_6_T11}), .c ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, SubBytesIns_Inst_Sbox_6_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T16_U1 ( .a ({new_AGEMA_signal_6015, new_AGEMA_signal_6014, new_AGEMA_signal_6013, SubBytesIns_Inst_Sbox_6_T5}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T17_U1 ( .a ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T18_U1 ( .a ({ciphertext_s3[52], ciphertext_s2[52], ciphertext_s1[52], ciphertext_s0[52]}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_6_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T19_U1 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_6027, new_AGEMA_signal_6026, new_AGEMA_signal_6025, SubBytesIns_Inst_Sbox_6_T18}), .c ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T20_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}), .c ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T21_U1 ( .a ({ciphertext_s3[49], ciphertext_s2[49], ciphertext_s1[49], ciphertext_s0[49]}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_6_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T22_U1 ( .a ({new_AGEMA_signal_6018, new_AGEMA_signal_6017, new_AGEMA_signal_6016, SubBytesIns_Inst_Sbox_6_T7}), .b ({new_AGEMA_signal_6030, new_AGEMA_signal_6029, new_AGEMA_signal_6028, SubBytesIns_Inst_Sbox_6_T21}), .c ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T23_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}), .c ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_6_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T24_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}), .c ({new_AGEMA_signal_7833, new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_6_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T25_U1 ( .a ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}), .c ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, new_AGEMA_signal_7834, SubBytesIns_Inst_Sbox_6_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T26_U1 ( .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .c ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_6_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_T27_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6024, new_AGEMA_signal_6023, new_AGEMA_signal_6022, SubBytesIns_Inst_Sbox_6_T12}), .c ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_6_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T1_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T2_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T3_U1 ( .a ({ciphertext_s3[63], ciphertext_s2[63], ciphertext_s1[63], ciphertext_s0[63]}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T4_U1 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T5_U1 ( .a ({ciphertext_s3[59], ciphertext_s2[59], ciphertext_s1[59], ciphertext_s0[59]}), .b ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T6_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}), .c ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T7_U1 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T8_U1 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .c ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_7_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T9_U1 ( .a ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T10_U1 ( .a ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .c ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T11_U1 ( .a ({ciphertext_s3[62], ciphertext_s2[62], ciphertext_s1[62], ciphertext_s0[62]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T12_U1 ( .a ({ciphertext_s3[61], ciphertext_s2[61], ciphertext_s1[61], ciphertext_s0[61]}), .b ({ciphertext_s3[58], ciphertext_s2[58], ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T13_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}), .c ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_7_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T14_U1 ( .a ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .b ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_7_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T15_U1 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_6051, new_AGEMA_signal_6050, new_AGEMA_signal_6049, SubBytesIns_Inst_Sbox_7_T11}), .c ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_7_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T16_U1 ( .a ({new_AGEMA_signal_6045, new_AGEMA_signal_6044, new_AGEMA_signal_6043, SubBytesIns_Inst_Sbox_7_T5}), .b ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T17_U1 ( .a ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T18_U1 ( .a ({ciphertext_s3[60], ciphertext_s2[60], ciphertext_s1[60], ciphertext_s0[60]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_7_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T19_U1 ( .a ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_6057, new_AGEMA_signal_6056, new_AGEMA_signal_6055, SubBytesIns_Inst_Sbox_7_T18}), .c ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T20_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}), .c ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T21_U1 ( .a ({ciphertext_s3[57], ciphertext_s2[57], ciphertext_s1[57], ciphertext_s0[57]}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_7_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T22_U1 ( .a ({new_AGEMA_signal_6048, new_AGEMA_signal_6047, new_AGEMA_signal_6046, SubBytesIns_Inst_Sbox_7_T7}), .b ({new_AGEMA_signal_6060, new_AGEMA_signal_6059, new_AGEMA_signal_6058, SubBytesIns_Inst_Sbox_7_T21}), .c ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T23_U1 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}), .c ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_7_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T24_U1 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}), .c ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, new_AGEMA_signal_7858, SubBytesIns_Inst_Sbox_7_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T25_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}), .c ({new_AGEMA_signal_7863, new_AGEMA_signal_7862, new_AGEMA_signal_7861, SubBytesIns_Inst_Sbox_7_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T26_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .c ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_7_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_T27_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6054, new_AGEMA_signal_6053, new_AGEMA_signal_6052, SubBytesIns_Inst_Sbox_7_T12}), .c ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_7_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T1_U1 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T2_U1 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T3_U1 ( .a ({ciphertext_s3[71], ciphertext_s2[71], ciphertext_s1[71], ciphertext_s0[71]}), .b ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T4_U1 ( .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T5_U1 ( .a ({ciphertext_s3[67], ciphertext_s2[67], ciphertext_s1[67], ciphertext_s0[67]}), .b ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T6_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}), .c ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T7_U1 ( .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T8_U1 ( .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .c ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_8_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T9_U1 ( .a ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T10_U1 ( .a ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .c ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T11_U1 ( .a ({ciphertext_s3[70], ciphertext_s2[70], ciphertext_s1[70], ciphertext_s0[70]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_8_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T12_U1 ( .a ({ciphertext_s3[69], ciphertext_s2[69], ciphertext_s1[69], ciphertext_s0[69]}), .b ({ciphertext_s3[66], ciphertext_s2[66], ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_8_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T13_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}), .c ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_8_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T14_U1 ( .a ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_8_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T15_U1 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_6081, new_AGEMA_signal_6080, new_AGEMA_signal_6079, SubBytesIns_Inst_Sbox_8_T11}), .c ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_8_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T16_U1 ( .a ({new_AGEMA_signal_6075, new_AGEMA_signal_6074, new_AGEMA_signal_6073, SubBytesIns_Inst_Sbox_8_T5}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T17_U1 ( .a ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T18_U1 ( .a ({ciphertext_s3[68], ciphertext_s2[68], ciphertext_s1[68], ciphertext_s0[68]}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_8_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T19_U1 ( .a ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_6087, new_AGEMA_signal_6086, new_AGEMA_signal_6085, SubBytesIns_Inst_Sbox_8_T18}), .c ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T20_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}), .c ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T21_U1 ( .a ({ciphertext_s3[65], ciphertext_s2[65], ciphertext_s1[65], ciphertext_s0[65]}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_8_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T22_U1 ( .a ({new_AGEMA_signal_6078, new_AGEMA_signal_6077, new_AGEMA_signal_6076, SubBytesIns_Inst_Sbox_8_T7}), .b ({new_AGEMA_signal_6090, new_AGEMA_signal_6089, new_AGEMA_signal_6088, SubBytesIns_Inst_Sbox_8_T21}), .c ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T23_U1 ( .a ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}), .c ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, SubBytesIns_Inst_Sbox_8_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T24_U1 ( .a ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}), .c ({new_AGEMA_signal_7887, new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_8_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T25_U1 ( .a ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}), .c ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, new_AGEMA_signal_7888, SubBytesIns_Inst_Sbox_8_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T26_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .c ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_T27_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6084, new_AGEMA_signal_6083, new_AGEMA_signal_6082, SubBytesIns_Inst_Sbox_8_T12}), .c ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_8_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T1_U1 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T2_U1 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T3_U1 ( .a ({ciphertext_s3[79], ciphertext_s2[79], ciphertext_s1[79], ciphertext_s0[79]}), .b ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T4_U1 ( .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T5_U1 ( .a ({ciphertext_s3[75], ciphertext_s2[75], ciphertext_s1[75], ciphertext_s0[75]}), .b ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T6_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}), .c ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T7_U1 ( .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T8_U1 ( .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .c ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_9_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T9_U1 ( .a ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T10_U1 ( .a ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .c ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T11_U1 ( .a ({ciphertext_s3[78], ciphertext_s2[78], ciphertext_s1[78], ciphertext_s0[78]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, SubBytesIns_Inst_Sbox_9_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T12_U1 ( .a ({ciphertext_s3[77], ciphertext_s2[77], ciphertext_s1[77], ciphertext_s0[77]}), .b ({ciphertext_s3[74], ciphertext_s2[74], ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, SubBytesIns_Inst_Sbox_9_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T13_U1 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}), .c ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_9_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T14_U1 ( .a ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .b ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_9_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T15_U1 ( .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_6111, new_AGEMA_signal_6110, new_AGEMA_signal_6109, SubBytesIns_Inst_Sbox_9_T11}), .c ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_9_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T16_U1 ( .a ({new_AGEMA_signal_6105, new_AGEMA_signal_6104, new_AGEMA_signal_6103, SubBytesIns_Inst_Sbox_9_T5}), .b ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T17_U1 ( .a ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T18_U1 ( .a ({ciphertext_s3[76], ciphertext_s2[76], ciphertext_s1[76], ciphertext_s0[76]}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_9_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T19_U1 ( .a ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_6117, new_AGEMA_signal_6116, new_AGEMA_signal_6115, SubBytesIns_Inst_Sbox_9_T18}), .c ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T20_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}), .c ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T21_U1 ( .a ({ciphertext_s3[73], ciphertext_s2[73], ciphertext_s1[73], ciphertext_s0[73]}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_9_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T22_U1 ( .a ({new_AGEMA_signal_6108, new_AGEMA_signal_6107, new_AGEMA_signal_6106, SubBytesIns_Inst_Sbox_9_T7}), .b ({new_AGEMA_signal_6120, new_AGEMA_signal_6119, new_AGEMA_signal_6118, SubBytesIns_Inst_Sbox_9_T21}), .c ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T23_U1 ( .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}), .c ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_9_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T24_U1 ( .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}), .c ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, new_AGEMA_signal_7912, SubBytesIns_Inst_Sbox_9_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T25_U1 ( .a ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}), .c ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_9_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T26_U1 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .c ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_9_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_T27_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6114, new_AGEMA_signal_6113, new_AGEMA_signal_6112, SubBytesIns_Inst_Sbox_9_T12}), .c ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_9_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T1_U1 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T2_U1 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T3_U1 ( .a ({ciphertext_s3[87], ciphertext_s2[87], ciphertext_s1[87], ciphertext_s0[87]}), .b ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T4_U1 ( .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T5_U1 ( .a ({ciphertext_s3[83], ciphertext_s2[83], ciphertext_s1[83], ciphertext_s0[83]}), .b ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T6_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}), .c ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T7_U1 ( .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T8_U1 ( .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .c ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_10_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T9_U1 ( .a ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T10_U1 ( .a ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .c ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T11_U1 ( .a ({ciphertext_s3[86], ciphertext_s2[86], ciphertext_s1[86], ciphertext_s0[86]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_10_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T12_U1 ( .a ({ciphertext_s3[85], ciphertext_s2[85], ciphertext_s1[85], ciphertext_s0[85]}), .b ({ciphertext_s3[82], ciphertext_s2[82], ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_10_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T13_U1 ( .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}), .c ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_10_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T14_U1 ( .a ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .b ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_10_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T15_U1 ( .a ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_6141, new_AGEMA_signal_6140, new_AGEMA_signal_6139, SubBytesIns_Inst_Sbox_10_T11}), .c ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_10_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T16_U1 ( .a ({new_AGEMA_signal_6135, new_AGEMA_signal_6134, new_AGEMA_signal_6133, SubBytesIns_Inst_Sbox_10_T5}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T17_U1 ( .a ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T18_U1 ( .a ({ciphertext_s3[84], ciphertext_s2[84], ciphertext_s1[84], ciphertext_s0[84]}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_10_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T19_U1 ( .a ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_6147, new_AGEMA_signal_6146, new_AGEMA_signal_6145, SubBytesIns_Inst_Sbox_10_T18}), .c ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T20_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}), .c ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T21_U1 ( .a ({ciphertext_s3[81], ciphertext_s2[81], ciphertext_s1[81], ciphertext_s0[81]}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_10_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T22_U1 ( .a ({new_AGEMA_signal_6138, new_AGEMA_signal_6137, new_AGEMA_signal_6136, SubBytesIns_Inst_Sbox_10_T7}), .b ({new_AGEMA_signal_6150, new_AGEMA_signal_6149, new_AGEMA_signal_6148, SubBytesIns_Inst_Sbox_10_T21}), .c ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T23_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}), .c ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_10_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T24_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}), .c ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_10_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T25_U1 ( .a ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}), .c ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, new_AGEMA_signal_7942, SubBytesIns_Inst_Sbox_10_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T26_U1 ( .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .c ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_10_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_T27_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6144, new_AGEMA_signal_6143, new_AGEMA_signal_6142, SubBytesIns_Inst_Sbox_10_T12}), .c ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_10_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T1_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T2_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T3_U1 ( .a ({ciphertext_s3[95], ciphertext_s2[95], ciphertext_s1[95], ciphertext_s0[95]}), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T4_U1 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T5_U1 ( .a ({ciphertext_s3[91], ciphertext_s2[91], ciphertext_s1[91], ciphertext_s0[91]}), .b ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T6_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}), .c ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T7_U1 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T8_U1 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .c ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, SubBytesIns_Inst_Sbox_11_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T9_U1 ( .a ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T10_U1 ( .a ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .c ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T11_U1 ( .a ({ciphertext_s3[94], ciphertext_s2[94], ciphertext_s1[94], ciphertext_s0[94]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T12_U1 ( .a ({ciphertext_s3[93], ciphertext_s2[93], ciphertext_s1[93], ciphertext_s0[93]}), .b ({ciphertext_s3[90], ciphertext_s2[90], ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T13_U1 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}), .c ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_11_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T14_U1 ( .a ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .b ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, new_AGEMA_signal_7372, SubBytesIns_Inst_Sbox_11_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T15_U1 ( .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_6171, new_AGEMA_signal_6170, new_AGEMA_signal_6169, SubBytesIns_Inst_Sbox_11_T11}), .c ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_11_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T16_U1 ( .a ({new_AGEMA_signal_6165, new_AGEMA_signal_6164, new_AGEMA_signal_6163, SubBytesIns_Inst_Sbox_11_T5}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T17_U1 ( .a ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T18_U1 ( .a ({ciphertext_s3[92], ciphertext_s2[92], ciphertext_s1[92], ciphertext_s0[92]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_6177, new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_11_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T19_U1 ( .a ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_6177, new_AGEMA_signal_6176, new_AGEMA_signal_6175, SubBytesIns_Inst_Sbox_11_T18}), .c ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T20_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}), .c ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T21_U1 ( .a ({ciphertext_s3[89], ciphertext_s2[89], ciphertext_s1[89], ciphertext_s0[89]}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_11_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T22_U1 ( .a ({new_AGEMA_signal_6168, new_AGEMA_signal_6167, new_AGEMA_signal_6166, SubBytesIns_Inst_Sbox_11_T7}), .b ({new_AGEMA_signal_6180, new_AGEMA_signal_6179, new_AGEMA_signal_6178, SubBytesIns_Inst_Sbox_11_T21}), .c ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T23_U1 ( .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}), .c ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_11_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T24_U1 ( .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}), .c ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, new_AGEMA_signal_7966, SubBytesIns_Inst_Sbox_11_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T25_U1 ( .a ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}), .c ({new_AGEMA_signal_7971, new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_11_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T26_U1 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .c ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, new_AGEMA_signal_7384, SubBytesIns_Inst_Sbox_11_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_T27_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6174, new_AGEMA_signal_6173, new_AGEMA_signal_6172, SubBytesIns_Inst_Sbox_11_T12}), .c ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_11_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T1_U1 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T2_U1 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T3_U1 ( .a ({ciphertext_s3[103], ciphertext_s2[103], ciphertext_s1[103], ciphertext_s0[103]}), .b ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T4_U1 ( .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T5_U1 ( .a ({ciphertext_s3[99], ciphertext_s2[99], ciphertext_s1[99], ciphertext_s0[99]}), .b ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T6_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}), .c ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T7_U1 ( .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T8_U1 ( .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .c ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T9_U1 ( .a ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .b ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T10_U1 ( .a ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .c ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T11_U1 ( .a ({ciphertext_s3[102], ciphertext_s2[102], ciphertext_s1[102], ciphertext_s0[102]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_12_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T12_U1 ( .a ({ciphertext_s3[101], ciphertext_s2[101], ciphertext_s1[101], ciphertext_s0[101]}), .b ({ciphertext_s3[98], ciphertext_s2[98], ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, SubBytesIns_Inst_Sbox_12_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T13_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}), .c ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_12_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T14_U1 ( .a ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T15_U1 ( .a ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_6201, new_AGEMA_signal_6200, new_AGEMA_signal_6199, SubBytesIns_Inst_Sbox_12_T11}), .c ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_12_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T16_U1 ( .a ({new_AGEMA_signal_6195, new_AGEMA_signal_6194, new_AGEMA_signal_6193, SubBytesIns_Inst_Sbox_12_T5}), .b ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T17_U1 ( .a ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T18_U1 ( .a ({ciphertext_s3[100], ciphertext_s2[100], ciphertext_s1[100], ciphertext_s0[100]}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_6207, new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_12_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T19_U1 ( .a ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_6207, new_AGEMA_signal_6206, new_AGEMA_signal_6205, SubBytesIns_Inst_Sbox_12_T18}), .c ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T20_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}), .c ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T21_U1 ( .a ({ciphertext_s3[97], ciphertext_s2[97], ciphertext_s1[97], ciphertext_s0[97]}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, new_AGEMA_signal_6208, SubBytesIns_Inst_Sbox_12_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T22_U1 ( .a ({new_AGEMA_signal_6198, new_AGEMA_signal_6197, new_AGEMA_signal_6196, SubBytesIns_Inst_Sbox_12_T7}), .b ({new_AGEMA_signal_6210, new_AGEMA_signal_6209, new_AGEMA_signal_6208, SubBytesIns_Inst_Sbox_12_T21}), .c ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T23_U1 ( .a ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}), .c ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, SubBytesIns_Inst_Sbox_12_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T24_U1 ( .a ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}), .c ({new_AGEMA_signal_7995, new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_12_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T25_U1 ( .a ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}), .c ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, new_AGEMA_signal_7996, SubBytesIns_Inst_Sbox_12_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T26_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .c ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_12_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_T27_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6204, new_AGEMA_signal_6203, new_AGEMA_signal_6202, SubBytesIns_Inst_Sbox_12_T12}), .c ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T1_U1 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T2_U1 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T3_U1 ( .a ({ciphertext_s3[111], ciphertext_s2[111], ciphertext_s1[111], ciphertext_s0[111]}), .b ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T4_U1 ( .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T5_U1 ( .a ({ciphertext_s3[107], ciphertext_s2[107], ciphertext_s1[107], ciphertext_s0[107]}), .b ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T6_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}), .c ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T7_U1 ( .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T8_U1 ( .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .c ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, SubBytesIns_Inst_Sbox_13_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T9_U1 ( .a ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T10_U1 ( .a ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .c ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T11_U1 ( .a ({ciphertext_s3[110], ciphertext_s2[110], ciphertext_s1[110], ciphertext_s0[110]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_13_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T12_U1 ( .a ({ciphertext_s3[109], ciphertext_s2[109], ciphertext_s1[109], ciphertext_s0[109]}), .b ({ciphertext_s3[106], ciphertext_s2[106], ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_13_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T13_U1 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}), .c ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_13_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T14_U1 ( .a ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .b ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, new_AGEMA_signal_7450, SubBytesIns_Inst_Sbox_13_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T15_U1 ( .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_6231, new_AGEMA_signal_6230, new_AGEMA_signal_6229, SubBytesIns_Inst_Sbox_13_T11}), .c ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T16_U1 ( .a ({new_AGEMA_signal_6225, new_AGEMA_signal_6224, new_AGEMA_signal_6223, SubBytesIns_Inst_Sbox_13_T5}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T17_U1 ( .a ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T18_U1 ( .a ({ciphertext_s3[108], ciphertext_s2[108], ciphertext_s1[108], ciphertext_s0[108]}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_13_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T19_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_6237, new_AGEMA_signal_6236, new_AGEMA_signal_6235, SubBytesIns_Inst_Sbox_13_T18}), .c ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T20_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}), .c ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T21_U1 ( .a ({ciphertext_s3[105], ciphertext_s2[105], ciphertext_s1[105], ciphertext_s0[105]}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_13_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T22_U1 ( .a ({new_AGEMA_signal_6228, new_AGEMA_signal_6227, new_AGEMA_signal_6226, SubBytesIns_Inst_Sbox_13_T7}), .b ({new_AGEMA_signal_6240, new_AGEMA_signal_6239, new_AGEMA_signal_6238, SubBytesIns_Inst_Sbox_13_T21}), .c ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T23_U1 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}), .c ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, SubBytesIns_Inst_Sbox_13_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T24_U1 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}), .c ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, new_AGEMA_signal_8020, SubBytesIns_Inst_Sbox_13_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T25_U1 ( .a ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}), .c ({new_AGEMA_signal_8025, new_AGEMA_signal_8024, new_AGEMA_signal_8023, SubBytesIns_Inst_Sbox_13_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T26_U1 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .c ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, new_AGEMA_signal_7462, SubBytesIns_Inst_Sbox_13_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_T27_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6234, new_AGEMA_signal_6233, new_AGEMA_signal_6232, SubBytesIns_Inst_Sbox_13_T12}), .c ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_13_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T1_U1 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T2_U1 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T3_U1 ( .a ({ciphertext_s3[119], ciphertext_s2[119], ciphertext_s1[119], ciphertext_s0[119]}), .b ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T4_U1 ( .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T5_U1 ( .a ({ciphertext_s3[115], ciphertext_s2[115], ciphertext_s1[115], ciphertext_s0[115]}), .b ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T6_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}), .c ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T7_U1 ( .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T8_U1 ( .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .c ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_14_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T9_U1 ( .a ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .b ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T10_U1 ( .a ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .c ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T11_U1 ( .a ({ciphertext_s3[118], ciphertext_s2[118], ciphertext_s1[118], ciphertext_s0[118]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_14_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T12_U1 ( .a ({ciphertext_s3[117], ciphertext_s2[117], ciphertext_s1[117], ciphertext_s0[117]}), .b ({ciphertext_s3[114], ciphertext_s2[114], ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_14_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T13_U1 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}), .c ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T14_U1 ( .a ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_14_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T15_U1 ( .a ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_6261, new_AGEMA_signal_6260, new_AGEMA_signal_6259, SubBytesIns_Inst_Sbox_14_T11}), .c ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_14_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T16_U1 ( .a ({new_AGEMA_signal_6255, new_AGEMA_signal_6254, new_AGEMA_signal_6253, SubBytesIns_Inst_Sbox_14_T5}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T17_U1 ( .a ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T18_U1 ( .a ({ciphertext_s3[116], ciphertext_s2[116], ciphertext_s1[116], ciphertext_s0[116]}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_6267, new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T19_U1 ( .a ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_6267, new_AGEMA_signal_6266, new_AGEMA_signal_6265, SubBytesIns_Inst_Sbox_14_T18}), .c ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T20_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}), .c ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T21_U1 ( .a ({ciphertext_s3[113], ciphertext_s2[113], ciphertext_s1[113], ciphertext_s0[113]}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T22_U1 ( .a ({new_AGEMA_signal_6258, new_AGEMA_signal_6257, new_AGEMA_signal_6256, SubBytesIns_Inst_Sbox_14_T7}), .b ({new_AGEMA_signal_6270, new_AGEMA_signal_6269, new_AGEMA_signal_6268, SubBytesIns_Inst_Sbox_14_T21}), .c ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T23_U1 ( .a ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}), .c ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, SubBytesIns_Inst_Sbox_14_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T24_U1 ( .a ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}), .c ({new_AGEMA_signal_8049, new_AGEMA_signal_8048, new_AGEMA_signal_8047, SubBytesIns_Inst_Sbox_14_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T25_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}), .c ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, new_AGEMA_signal_8050, SubBytesIns_Inst_Sbox_14_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T26_U1 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .c ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_14_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_T27_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6264, new_AGEMA_signal_6263, new_AGEMA_signal_6262, SubBytesIns_Inst_Sbox_14_T12}), .c ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, SubBytesIns_Inst_Sbox_14_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T1_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T2_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T3_U1 ( .a ({ciphertext_s3[127], ciphertext_s2[127], ciphertext_s1[127], ciphertext_s0[127]}), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T4_U1 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T5_U1 ( .a ({ciphertext_s3[123], ciphertext_s2[123], ciphertext_s1[123], ciphertext_s0[123]}), .b ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T6_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}), .c ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T7_U1 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T8_U1 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .c ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, SubBytesIns_Inst_Sbox_15_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T9_U1 ( .a ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T10_U1 ( .a ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .c ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T11_U1 ( .a ({ciphertext_s3[126], ciphertext_s2[126], ciphertext_s1[126], ciphertext_s0[126]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_15_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T12_U1 ( .a ({ciphertext_s3[125], ciphertext_s2[125], ciphertext_s1[125], ciphertext_s0[125]}), .b ({ciphertext_s3[122], ciphertext_s2[122], ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, SubBytesIns_Inst_Sbox_15_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T13_U1 ( .a ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}), .c ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_15_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T14_U1 ( .a ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .b ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, new_AGEMA_signal_7528, SubBytesIns_Inst_Sbox_15_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T15_U1 ( .a ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_6291, new_AGEMA_signal_6290, new_AGEMA_signal_6289, SubBytesIns_Inst_Sbox_15_T11}), .c ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, SubBytesIns_Inst_Sbox_15_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T16_U1 ( .a ({new_AGEMA_signal_6285, new_AGEMA_signal_6284, new_AGEMA_signal_6283, SubBytesIns_Inst_Sbox_15_T5}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T17_U1 ( .a ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T18_U1 ( .a ({ciphertext_s3[124], ciphertext_s2[124], ciphertext_s1[124], ciphertext_s0[124]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_6297, new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_15_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T19_U1 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_6297, new_AGEMA_signal_6296, new_AGEMA_signal_6295, SubBytesIns_Inst_Sbox_15_T18}), .c ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T20_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}), .c ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T21_U1 ( .a ({ciphertext_s3[121], ciphertext_s2[121], ciphertext_s1[121], ciphertext_s0[121]}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, new_AGEMA_signal_6298, SubBytesIns_Inst_Sbox_15_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T22_U1 ( .a ({new_AGEMA_signal_6288, new_AGEMA_signal_6287, new_AGEMA_signal_6286, SubBytesIns_Inst_Sbox_15_T7}), .b ({new_AGEMA_signal_6300, new_AGEMA_signal_6299, new_AGEMA_signal_6298, SubBytesIns_Inst_Sbox_15_T21}), .c ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T23_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}), .c ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_15_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T24_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}), .c ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, new_AGEMA_signal_8074, SubBytesIns_Inst_Sbox_15_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T25_U1 ( .a ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}), .c ({new_AGEMA_signal_8079, new_AGEMA_signal_8078, new_AGEMA_signal_8077, SubBytesIns_Inst_Sbox_15_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T26_U1 ( .a ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .c ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, new_AGEMA_signal_7540, SubBytesIns_Inst_Sbox_15_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_T27_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6294, new_AGEMA_signal_6293, new_AGEMA_signal_6292, SubBytesIns_Inst_Sbox_15_T12}), .c ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, SubBytesIns_Inst_Sbox_15_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T1_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .c ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T2_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T3_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .c ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T4_U1 ( .a ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T5_U1 ( .a ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}), .b ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .c ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T6_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .c ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T7_U1 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .b ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .c ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T8_U1 ( .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .c ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T9_U1 ( .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T10_U1 ( .a ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .c ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T11_U1 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T12_U1 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .c ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T13_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .c ({new_AGEMA_signal_6309, new_AGEMA_signal_6308, new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T14_U1 ( .a ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T15_U1 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5721, new_AGEMA_signal_5720, new_AGEMA_signal_5719, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T11}), .c ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T16_U1 ( .a ({new_AGEMA_signal_5715, new_AGEMA_signal_5714, new_AGEMA_signal_5713, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T5}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T17_U1 ( .a ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T18_U1 ( .a ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .c ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T19_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5727, new_AGEMA_signal_5726, new_AGEMA_signal_5725, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T18}), .c ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T20_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .c ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T21_U1 ( .a ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .c ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T22_U1 ( .a ({new_AGEMA_signal_5718, new_AGEMA_signal_5717, new_AGEMA_signal_5716, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T7}), .b ({new_AGEMA_signal_5730, new_AGEMA_signal_5729, new_AGEMA_signal_5728, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T21}), .c ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T23_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .c ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T24_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .c ({new_AGEMA_signal_7563, new_AGEMA_signal_7562, new_AGEMA_signal_7561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T25_U1 ( .a ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .c ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, new_AGEMA_signal_7564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T26_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .c ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, new_AGEMA_signal_6799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_T27_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_5724, new_AGEMA_signal_5723, new_AGEMA_signal_5722, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T12}), .c ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T1_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .c ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T2_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T3_U1 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .c ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T4_U1 ( .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T5_U1 ( .a ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}), .b ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .c ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T6_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .c ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T7_U1 ( .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .b ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .c ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T8_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .c ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T9_U1 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T10_U1 ( .a ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .c ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T11_U1 ( .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T12_U1 ( .a ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .b ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .c ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T13_U1 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .c ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T14_U1 ( .a ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, new_AGEMA_signal_6826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T15_U1 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5751, new_AGEMA_signal_5750, new_AGEMA_signal_5749, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T11}), .c ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T16_U1 ( .a ({new_AGEMA_signal_5745, new_AGEMA_signal_5744, new_AGEMA_signal_5743, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T5}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T17_U1 ( .a ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T18_U1 ( .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .c ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T19_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5757, new_AGEMA_signal_5756, new_AGEMA_signal_5755, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T18}), .c ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T20_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .c ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T21_U1 ( .a ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .c ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T22_U1 ( .a ({new_AGEMA_signal_5748, new_AGEMA_signal_5747, new_AGEMA_signal_5746, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T7}), .b ({new_AGEMA_signal_5760, new_AGEMA_signal_5759, new_AGEMA_signal_5758, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T21}), .c ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T23_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .c ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T24_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .c ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, new_AGEMA_signal_7588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T25_U1 ( .a ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .c ({new_AGEMA_signal_7593, new_AGEMA_signal_7592, new_AGEMA_signal_7591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T26_U1 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .c ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, new_AGEMA_signal_6838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_T27_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_5754, new_AGEMA_signal_5753, new_AGEMA_signal_5752, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T12}), .c ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T1_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .c ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T2_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T3_U1 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .c ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T4_U1 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T5_U1 ( .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}), .b ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .c ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T6_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .c ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T7_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .b ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .c ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T8_U1 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .c ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T9_U1 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T10_U1 ( .a ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .c ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T11_U1 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T12_U1 ( .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .b ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .c ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T13_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .c ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T14_U1 ( .a ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, new_AGEMA_signal_6865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T15_U1 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5781, new_AGEMA_signal_5780, new_AGEMA_signal_5779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T11}), .c ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T16_U1 ( .a ({new_AGEMA_signal_5775, new_AGEMA_signal_5774, new_AGEMA_signal_5773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T5}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T17_U1 ( .a ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T18_U1 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .c ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, new_AGEMA_signal_5785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T19_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5787, new_AGEMA_signal_5786, new_AGEMA_signal_5785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T18}), .c ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T20_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .c ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T21_U1 ( .a ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .c ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, new_AGEMA_signal_5788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T22_U1 ( .a ({new_AGEMA_signal_5778, new_AGEMA_signal_5777, new_AGEMA_signal_5776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T7}), .b ({new_AGEMA_signal_5790, new_AGEMA_signal_5789, new_AGEMA_signal_5788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T21}), .c ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T23_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .c ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T24_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .c ({new_AGEMA_signal_7617, new_AGEMA_signal_7616, new_AGEMA_signal_7615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T25_U1 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .c ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, new_AGEMA_signal_7618, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T26_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .c ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, new_AGEMA_signal_6877, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_T27_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_5784, new_AGEMA_signal_5783, new_AGEMA_signal_5782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T12}), .c ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T1_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .c ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T2_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T3_U1 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .c ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T4_U1 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T5_U1 ( .a ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}), .b ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .c ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T6_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .c ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T7_U1 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .c ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T8_U1 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .c ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T9_U1 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T10_U1 ( .a ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .c ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T11_U1 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T12_U1 ( .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .b ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .c ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T13_U1 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .c ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T14_U1 ( .a ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .b ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, new_AGEMA_signal_6904, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T15_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5811, new_AGEMA_signal_5810, new_AGEMA_signal_5809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T11}), .c ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T16_U1 ( .a ({new_AGEMA_signal_5805, new_AGEMA_signal_5804, new_AGEMA_signal_5803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T5}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T17_U1 ( .a ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T18_U1 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .c ({new_AGEMA_signal_5817, new_AGEMA_signal_5816, new_AGEMA_signal_5815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T19_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5817, new_AGEMA_signal_5816, new_AGEMA_signal_5815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T18}), .c ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T20_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .c ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T21_U1 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .c ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T22_U1 ( .a ({new_AGEMA_signal_5808, new_AGEMA_signal_5807, new_AGEMA_signal_5806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T7}), .b ({new_AGEMA_signal_5820, new_AGEMA_signal_5819, new_AGEMA_signal_5818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T21}), .c ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T23_U1 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .c ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T24_U1 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .c ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, new_AGEMA_signal_7642, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T25_U1 ( .a ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .c ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, new_AGEMA_signal_7645, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T26_U1 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .c ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, new_AGEMA_signal_6916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_T27_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_5814, new_AGEMA_signal_5813, new_AGEMA_signal_5812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T12}), .c ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}) ) ;
    INV_X1 RoundCounterIns_U14 ( .A (RoundCounterIns_n13), .ZN (RoundCounterIns_n1) ) ;
    MUX2_X1 RoundCounterIns_U13 ( .S (RoundCounterIns_n5), .A (RoundCounterIns_n12), .B (RoundCounterIns_n11), .Z (RoundCounterIns_n13) ) ;
    NOR2_X1 RoundCounterIns_U12 ( .A1 (reset), .A2 (RoundCounterIns_n10), .ZN (RoundCounterIns_N8) ) ;
    XNOR2_X1 RoundCounterIns_U11 ( .A (RoundCounter[0]), .B (RoundCounter[1]), .ZN (RoundCounterIns_n10) ) ;
    MUX2_X1 RoundCounterIns_U10 ( .S (RoundCounter[3]), .A (RoundCounterIns_n9), .B (RoundCounterIns_n8), .Z (RoundCounterIns_N10) ) ;
    NAND2_X1 RoundCounterIns_U9 ( .A1 (RoundCounterIns_n12), .A2 (RoundCounterIns_n7), .ZN (RoundCounterIns_n8) ) ;
    NAND2_X1 RoundCounterIns_U8 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n2), .ZN (RoundCounterIns_n7) ) ;
    NOR2_X1 RoundCounterIns_U7 ( .A1 (RoundCounterIns_n4), .A2 (RoundCounterIns_N7), .ZN (RoundCounterIns_n12) ) ;
    NOR2_X1 RoundCounterIns_U6 ( .A1 (RoundCounter[1]), .A2 (reset), .ZN (RoundCounterIns_n4) ) ;
    NOR2_X1 RoundCounterIns_U5 ( .A1 (RoundCounterIns_n5), .A2 (RoundCounterIns_n11), .ZN (RoundCounterIns_n9) ) ;
    NAND2_X1 RoundCounterIns_U4 ( .A1 (RoundCounter[1]), .A2 (RoundCounterIns_n3), .ZN (RoundCounterIns_n11) ) ;
    NOR2_X1 RoundCounterIns_U3 ( .A1 (reset), .A2 (RoundCounterIns_n6), .ZN (RoundCounterIns_n3) ) ;
    NOR2_X1 RoundCounterIns_U2 ( .A1 (reset), .A2 (RoundCounter[0]), .ZN (RoundCounterIns_N7) ) ;
    INV_X1 RoundCounterIns_U1 ( .A (reset), .ZN (RoundCounterIns_n2) ) ;
    INV_X1 RoundCounterIns_count_reg_0__U1 ( .A (RoundCounter[0]), .ZN (RoundCounterIns_n6) ) ;
    INV_X1 RoundCounterIns_count_reg_2__U1 ( .A (RoundCounter[2]), .ZN (RoundCounterIns_n5) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk (clk), .rst (reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, SubBytesIns_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, new_AGEMA_signal_7675, SubBytesIns_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_6945, new_AGEMA_signal_6944, new_AGEMA_signal_6943, SubBytesIns_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, new_AGEMA_signal_7678, SubBytesIns_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6963, new_AGEMA_signal_6962, new_AGEMA_signal_6961, SubBytesIns_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6960, new_AGEMA_signal_6959, new_AGEMA_signal_6958, SubBytesIns_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, SubBytesIns_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_6957, new_AGEMA_signal_6956, new_AGEMA_signal_6955, SubBytesIns_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, new_AGEMA_signal_7684, SubBytesIns_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_7689, new_AGEMA_signal_7688, new_AGEMA_signal_7687, SubBytesIns_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6966, new_AGEMA_signal_6965, new_AGEMA_signal_6964, SubBytesIns_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, SubBytesIns_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6975, new_AGEMA_signal_6974, new_AGEMA_signal_6973, SubBytesIns_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, SubBytesIns_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_7695, new_AGEMA_signal_7694, new_AGEMA_signal_7693, SubBytesIns_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6972, new_AGEMA_signal_6971, new_AGEMA_signal_6970, SubBytesIns_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, new_AGEMA_signal_8164, SubBytesIns_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_7680, new_AGEMA_signal_7679, new_AGEMA_signal_7678, SubBytesIns_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_7677, new_AGEMA_signal_7676, new_AGEMA_signal_7675, SubBytesIns_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_7683, new_AGEMA_signal_7682, new_AGEMA_signal_7681, SubBytesIns_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_7671, new_AGEMA_signal_7670, new_AGEMA_signal_7669, SubBytesIns_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, new_AGEMA_signal_8170, SubBytesIns_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_7686, new_AGEMA_signal_7685, new_AGEMA_signal_7684, SubBytesIns_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6969, new_AGEMA_signal_6968, new_AGEMA_signal_6967, SubBytesIns_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_8163, new_AGEMA_signal_8162, new_AGEMA_signal_8161, SubBytesIns_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, new_AGEMA_signal_8164, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8451, new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_8169, new_AGEMA_signal_8168, new_AGEMA_signal_8167, SubBytesIns_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_8172, new_AGEMA_signal_8171, new_AGEMA_signal_8170, SubBytesIns_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_8166, new_AGEMA_signal_8165, new_AGEMA_signal_8164, SubBytesIns_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_8175, new_AGEMA_signal_8174, new_AGEMA_signal_8173, SubBytesIns_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_7692, new_AGEMA_signal_7691, new_AGEMA_signal_7690, SubBytesIns_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_8451, new_AGEMA_signal_8450, new_AGEMA_signal_8449, SubBytesIns_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_7674, new_AGEMA_signal_7673, new_AGEMA_signal_7672, SubBytesIns_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, new_AGEMA_signal_7702, SubBytesIns_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_6984, new_AGEMA_signal_6983, new_AGEMA_signal_6982, SubBytesIns_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_7002, new_AGEMA_signal_7001, new_AGEMA_signal_7000, SubBytesIns_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6999, new_AGEMA_signal_6998, new_AGEMA_signal_6997, SubBytesIns_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, new_AGEMA_signal_7708, SubBytesIns_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_6996, new_AGEMA_signal_6995, new_AGEMA_signal_6994, SubBytesIns_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, new_AGEMA_signal_7714, SubBytesIns_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_7716, new_AGEMA_signal_7715, new_AGEMA_signal_7714, SubBytesIns_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_7005, new_AGEMA_signal_7004, new_AGEMA_signal_7003, SubBytesIns_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, new_AGEMA_signal_8176, SubBytesIns_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_7014, new_AGEMA_signal_7013, new_AGEMA_signal_7012, SubBytesIns_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, new_AGEMA_signal_7720, SubBytesIns_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_7722, new_AGEMA_signal_7721, new_AGEMA_signal_7720, SubBytesIns_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_7011, new_AGEMA_signal_7010, new_AGEMA_signal_7009, SubBytesIns_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_7707, new_AGEMA_signal_7706, new_AGEMA_signal_7705, SubBytesIns_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_7704, new_AGEMA_signal_7703, new_AGEMA_signal_7702, SubBytesIns_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, new_AGEMA_signal_8182, SubBytesIns_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_7710, new_AGEMA_signal_7709, new_AGEMA_signal_7708, SubBytesIns_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_7698, new_AGEMA_signal_7697, new_AGEMA_signal_7696, SubBytesIns_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_7713, new_AGEMA_signal_7712, new_AGEMA_signal_7711, SubBytesIns_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_7008, new_AGEMA_signal_7007, new_AGEMA_signal_7006, SubBytesIns_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, new_AGEMA_signal_8188, SubBytesIns_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_8178, new_AGEMA_signal_8177, new_AGEMA_signal_8176, SubBytesIns_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8463, new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_8184, new_AGEMA_signal_8183, new_AGEMA_signal_8182, SubBytesIns_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_8187, new_AGEMA_signal_8186, new_AGEMA_signal_8185, SubBytesIns_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_8181, new_AGEMA_signal_8180, new_AGEMA_signal_8179, SubBytesIns_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_8190, new_AGEMA_signal_8189, new_AGEMA_signal_8188, SubBytesIns_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_7719, new_AGEMA_signal_7718, new_AGEMA_signal_7717, SubBytesIns_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_8463, new_AGEMA_signal_8462, new_AGEMA_signal_8461, SubBytesIns_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_7701, new_AGEMA_signal_7700, new_AGEMA_signal_7699, SubBytesIns_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, new_AGEMA_signal_8956, SubBytesIns_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_7023, new_AGEMA_signal_7022, new_AGEMA_signal_7021, SubBytesIns_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, new_AGEMA_signal_7732, SubBytesIns_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_7041, new_AGEMA_signal_7040, new_AGEMA_signal_7039, SubBytesIns_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_7038, new_AGEMA_signal_7037, new_AGEMA_signal_7036, SubBytesIns_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126]}), .c ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132]}), .c ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_7035, new_AGEMA_signal_7034, new_AGEMA_signal_7033, SubBytesIns_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, new_AGEMA_signal_7738, SubBytesIns_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138]}), .c ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_7743, new_AGEMA_signal_7742, new_AGEMA_signal_7741, SubBytesIns_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_7044, new_AGEMA_signal_7043, new_AGEMA_signal_7042, SubBytesIns_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .c ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150]}), .c ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_7053, new_AGEMA_signal_7052, new_AGEMA_signal_7051, SubBytesIns_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, SubBytesIns_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156]}), .c ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_7749, new_AGEMA_signal_7748, new_AGEMA_signal_7747, SubBytesIns_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_7050, new_AGEMA_signal_7049, new_AGEMA_signal_7048, SubBytesIns_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, new_AGEMA_signal_8194, SubBytesIns_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_7734, new_AGEMA_signal_7733, new_AGEMA_signal_7732, SubBytesIns_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_7731, new_AGEMA_signal_7730, new_AGEMA_signal_7729, SubBytesIns_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_7737, new_AGEMA_signal_7736, new_AGEMA_signal_7735, SubBytesIns_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_7725, new_AGEMA_signal_7724, new_AGEMA_signal_7723, SubBytesIns_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, new_AGEMA_signal_8200, SubBytesIns_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_7740, new_AGEMA_signal_7739, new_AGEMA_signal_7738, SubBytesIns_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_7047, new_AGEMA_signal_7046, new_AGEMA_signal_7045, SubBytesIns_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_8193, new_AGEMA_signal_8192, new_AGEMA_signal_8191, SubBytesIns_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, new_AGEMA_signal_8194, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8475, new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_8199, new_AGEMA_signal_8198, new_AGEMA_signal_8197, SubBytesIns_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_8202, new_AGEMA_signal_8201, new_AGEMA_signal_8200, SubBytesIns_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_8196, new_AGEMA_signal_8195, new_AGEMA_signal_8194, SubBytesIns_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_8205, new_AGEMA_signal_8204, new_AGEMA_signal_8203, SubBytesIns_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_7746, new_AGEMA_signal_7745, new_AGEMA_signal_7744, SubBytesIns_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_8475, new_AGEMA_signal_8474, new_AGEMA_signal_8473, SubBytesIns_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_7728, new_AGEMA_signal_7727, new_AGEMA_signal_7726, SubBytesIns_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, new_AGEMA_signal_8971, SubBytesIns_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162]}), .c ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168]}), .c ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, new_AGEMA_signal_7756, SubBytesIns_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_7062, new_AGEMA_signal_7061, new_AGEMA_signal_7060, SubBytesIns_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174]}), .c ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_7080, new_AGEMA_signal_7079, new_AGEMA_signal_7078, SubBytesIns_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_7077, new_AGEMA_signal_7076, new_AGEMA_signal_7075, SubBytesIns_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, new_AGEMA_signal_7762, SubBytesIns_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180]}), .c ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186]}), .c ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_7074, new_AGEMA_signal_7073, new_AGEMA_signal_7072, SubBytesIns_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .c ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, new_AGEMA_signal_7768, SubBytesIns_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_7770, new_AGEMA_signal_7769, new_AGEMA_signal_7768, SubBytesIns_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_7083, new_AGEMA_signal_7082, new_AGEMA_signal_7081, SubBytesIns_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, new_AGEMA_signal_8206, SubBytesIns_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198]}), .c ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204]}), .c ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_7092, new_AGEMA_signal_7091, new_AGEMA_signal_7090, SubBytesIns_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210]}), .c ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, new_AGEMA_signal_7774, SubBytesIns_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_7776, new_AGEMA_signal_7775, new_AGEMA_signal_7774, SubBytesIns_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_7089, new_AGEMA_signal_7088, new_AGEMA_signal_7087, SubBytesIns_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_7761, new_AGEMA_signal_7760, new_AGEMA_signal_7759, SubBytesIns_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_7758, new_AGEMA_signal_7757, new_AGEMA_signal_7756, SubBytesIns_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, new_AGEMA_signal_8212, SubBytesIns_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_7764, new_AGEMA_signal_7763, new_AGEMA_signal_7762, SubBytesIns_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_7752, new_AGEMA_signal_7751, new_AGEMA_signal_7750, SubBytesIns_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_7767, new_AGEMA_signal_7766, new_AGEMA_signal_7765, SubBytesIns_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_7086, new_AGEMA_signal_7085, new_AGEMA_signal_7084, SubBytesIns_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, new_AGEMA_signal_8218, SubBytesIns_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_8208, new_AGEMA_signal_8207, new_AGEMA_signal_8206, SubBytesIns_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8487, new_AGEMA_signal_8486, new_AGEMA_signal_8485, SubBytesIns_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_8214, new_AGEMA_signal_8213, new_AGEMA_signal_8212, SubBytesIns_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_8217, new_AGEMA_signal_8216, new_AGEMA_signal_8215, SubBytesIns_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_8211, new_AGEMA_signal_8210, new_AGEMA_signal_8209, SubBytesIns_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_8220, new_AGEMA_signal_8219, new_AGEMA_signal_8218, SubBytesIns_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_7773, new_AGEMA_signal_7772, new_AGEMA_signal_7771, SubBytesIns_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_8487, new_AGEMA_signal_8486, new_AGEMA_signal_8485, SubBytesIns_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_7755, new_AGEMA_signal_7754, new_AGEMA_signal_7753, SubBytesIns_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, new_AGEMA_signal_8986, SubBytesIns_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_3_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M1_U1 ( .a ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_4_T13}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216]}), .c ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_4_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M2_U1 ( .a ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_4_T23}), .b ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222]}), .c ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_4_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M3_U1 ( .a ({new_AGEMA_signal_7101, new_AGEMA_signal_7100, new_AGEMA_signal_7099, SubBytesIns_Inst_Sbox_4_T14}), .b ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, new_AGEMA_signal_7786, SubBytesIns_Inst_Sbox_4_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M4_U1 ( .a ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228]}), .c ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_4_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M5_U1 ( .a ({new_AGEMA_signal_7119, new_AGEMA_signal_7118, new_AGEMA_signal_7117, SubBytesIns_Inst_Sbox_4_M4}), .b ({new_AGEMA_signal_7116, new_AGEMA_signal_7115, new_AGEMA_signal_7114, SubBytesIns_Inst_Sbox_4_M1}), .c ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_4_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M6_U1 ( .a ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234]}), .c ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_4_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M7_U1 ( .a ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .c ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_4_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M8_U1 ( .a ({new_AGEMA_signal_7113, new_AGEMA_signal_7112, new_AGEMA_signal_7111, SubBytesIns_Inst_Sbox_4_T26}), .b ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, new_AGEMA_signal_7792, SubBytesIns_Inst_Sbox_4_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M9_U1 ( .a ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}), .b ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246]}), .c ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_4_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M10_U1 ( .a ({new_AGEMA_signal_7797, new_AGEMA_signal_7796, new_AGEMA_signal_7795, SubBytesIns_Inst_Sbox_4_M9}), .b ({new_AGEMA_signal_7122, new_AGEMA_signal_7121, new_AGEMA_signal_7120, SubBytesIns_Inst_Sbox_4_M6}), .c ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_4_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M11_U1 ( .a ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .b ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252]}), .c ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_4_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M12_U1 ( .a ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}), .b ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258]}), .c ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_4_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M13_U1 ( .a ({new_AGEMA_signal_7131, new_AGEMA_signal_7130, new_AGEMA_signal_7129, SubBytesIns_Inst_Sbox_4_M12}), .b ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, SubBytesIns_Inst_Sbox_4_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M14_U1 ( .a ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .b ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264]}), .c ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_4_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M15_U1 ( .a ({new_AGEMA_signal_7803, new_AGEMA_signal_7802, new_AGEMA_signal_7801, SubBytesIns_Inst_Sbox_4_M14}), .b ({new_AGEMA_signal_7128, new_AGEMA_signal_7127, new_AGEMA_signal_7126, SubBytesIns_Inst_Sbox_4_M11}), .c ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, new_AGEMA_signal_8224, SubBytesIns_Inst_Sbox_4_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M16_U1 ( .a ({new_AGEMA_signal_7788, new_AGEMA_signal_7787, new_AGEMA_signal_7786, SubBytesIns_Inst_Sbox_4_M3}), .b ({new_AGEMA_signal_7785, new_AGEMA_signal_7784, new_AGEMA_signal_7783, SubBytesIns_Inst_Sbox_4_M2}), .c ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_4_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M17_U1 ( .a ({new_AGEMA_signal_7791, new_AGEMA_signal_7790, new_AGEMA_signal_7789, SubBytesIns_Inst_Sbox_4_M5}), .b ({new_AGEMA_signal_7779, new_AGEMA_signal_7778, new_AGEMA_signal_7777, SubBytesIns_Inst_Sbox_4_T24}), .c ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, new_AGEMA_signal_8230, SubBytesIns_Inst_Sbox_4_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M18_U1 ( .a ({new_AGEMA_signal_7794, new_AGEMA_signal_7793, new_AGEMA_signal_7792, SubBytesIns_Inst_Sbox_4_M8}), .b ({new_AGEMA_signal_7125, new_AGEMA_signal_7124, new_AGEMA_signal_7123, SubBytesIns_Inst_Sbox_4_M7}), .c ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_4_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M19_U1 ( .a ({new_AGEMA_signal_8223, new_AGEMA_signal_8222, new_AGEMA_signal_8221, SubBytesIns_Inst_Sbox_4_M10}), .b ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, new_AGEMA_signal_8224, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, new_AGEMA_signal_8497, SubBytesIns_Inst_Sbox_4_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M20_U1 ( .a ({new_AGEMA_signal_8229, new_AGEMA_signal_8228, new_AGEMA_signal_8227, SubBytesIns_Inst_Sbox_4_M16}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M21_U1 ( .a ({new_AGEMA_signal_8232, new_AGEMA_signal_8231, new_AGEMA_signal_8230, SubBytesIns_Inst_Sbox_4_M17}), .b ({new_AGEMA_signal_8226, new_AGEMA_signal_8225, new_AGEMA_signal_8224, SubBytesIns_Inst_Sbox_4_M15}), .c ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M22_U1 ( .a ({new_AGEMA_signal_8235, new_AGEMA_signal_8234, new_AGEMA_signal_8233, SubBytesIns_Inst_Sbox_4_M18}), .b ({new_AGEMA_signal_7800, new_AGEMA_signal_7799, new_AGEMA_signal_7798, SubBytesIns_Inst_Sbox_4_M13}), .c ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M23_U1 ( .a ({new_AGEMA_signal_8499, new_AGEMA_signal_8498, new_AGEMA_signal_8497, SubBytesIns_Inst_Sbox_4_M19}), .b ({new_AGEMA_signal_7782, new_AGEMA_signal_7781, new_AGEMA_signal_7780, SubBytesIns_Inst_Sbox_4_T25}), .c ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M24_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}), .c ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, new_AGEMA_signal_9001, SubBytesIns_Inst_Sbox_4_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M27_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}), .c ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_4_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M1_U1 ( .a ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_5_T13}), .b ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270]}), .c ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_5_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M2_U1 ( .a ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, SubBytesIns_Inst_Sbox_5_T23}), .b ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276]}), .c ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, new_AGEMA_signal_7810, SubBytesIns_Inst_Sbox_5_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M3_U1 ( .a ({new_AGEMA_signal_7140, new_AGEMA_signal_7139, new_AGEMA_signal_7138, SubBytesIns_Inst_Sbox_5_T14}), .b ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_7815, new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_5_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M4_U1 ( .a ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282]}), .c ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, new_AGEMA_signal_7156, SubBytesIns_Inst_Sbox_5_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M5_U1 ( .a ({new_AGEMA_signal_7158, new_AGEMA_signal_7157, new_AGEMA_signal_7156, SubBytesIns_Inst_Sbox_5_M4}), .b ({new_AGEMA_signal_7155, new_AGEMA_signal_7154, new_AGEMA_signal_7153, SubBytesIns_Inst_Sbox_5_M1}), .c ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, new_AGEMA_signal_7816, SubBytesIns_Inst_Sbox_5_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M6_U1 ( .a ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .c ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_5_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M7_U1 ( .a ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}), .b ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294]}), .c ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, new_AGEMA_signal_7162, SubBytesIns_Inst_Sbox_5_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M8_U1 ( .a ({new_AGEMA_signal_7152, new_AGEMA_signal_7151, new_AGEMA_signal_7150, SubBytesIns_Inst_Sbox_5_T26}), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_5_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M9_U1 ( .a ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}), .b ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300]}), .c ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, new_AGEMA_signal_7822, SubBytesIns_Inst_Sbox_5_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M10_U1 ( .a ({new_AGEMA_signal_7824, new_AGEMA_signal_7823, new_AGEMA_signal_7822, SubBytesIns_Inst_Sbox_5_M9}), .b ({new_AGEMA_signal_7161, new_AGEMA_signal_7160, new_AGEMA_signal_7159, SubBytesIns_Inst_Sbox_5_M6}), .c ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, new_AGEMA_signal_8236, SubBytesIns_Inst_Sbox_5_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M11_U1 ( .a ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306]}), .c ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_5_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M12_U1 ( .a ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}), .b ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312]}), .c ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, new_AGEMA_signal_7168, SubBytesIns_Inst_Sbox_5_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M13_U1 ( .a ({new_AGEMA_signal_7170, new_AGEMA_signal_7169, new_AGEMA_signal_7168, SubBytesIns_Inst_Sbox_5_M12}), .b ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_5_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M14_U1 ( .a ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318]}), .c ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, new_AGEMA_signal_7828, SubBytesIns_Inst_Sbox_5_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M15_U1 ( .a ({new_AGEMA_signal_7830, new_AGEMA_signal_7829, new_AGEMA_signal_7828, SubBytesIns_Inst_Sbox_5_M14}), .b ({new_AGEMA_signal_7167, new_AGEMA_signal_7166, new_AGEMA_signal_7165, SubBytesIns_Inst_Sbox_5_M11}), .c ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_5_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M16_U1 ( .a ({new_AGEMA_signal_7815, new_AGEMA_signal_7814, new_AGEMA_signal_7813, SubBytesIns_Inst_Sbox_5_M3}), .b ({new_AGEMA_signal_7812, new_AGEMA_signal_7811, new_AGEMA_signal_7810, SubBytesIns_Inst_Sbox_5_M2}), .c ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, new_AGEMA_signal_8242, SubBytesIns_Inst_Sbox_5_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M17_U1 ( .a ({new_AGEMA_signal_7818, new_AGEMA_signal_7817, new_AGEMA_signal_7816, SubBytesIns_Inst_Sbox_5_M5}), .b ({new_AGEMA_signal_7806, new_AGEMA_signal_7805, new_AGEMA_signal_7804, SubBytesIns_Inst_Sbox_5_T24}), .c ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_5_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M18_U1 ( .a ({new_AGEMA_signal_7821, new_AGEMA_signal_7820, new_AGEMA_signal_7819, SubBytesIns_Inst_Sbox_5_M8}), .b ({new_AGEMA_signal_7164, new_AGEMA_signal_7163, new_AGEMA_signal_7162, SubBytesIns_Inst_Sbox_5_M7}), .c ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, new_AGEMA_signal_8248, SubBytesIns_Inst_Sbox_5_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M19_U1 ( .a ({new_AGEMA_signal_8238, new_AGEMA_signal_8237, new_AGEMA_signal_8236, SubBytesIns_Inst_Sbox_5_M10}), .b ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, new_AGEMA_signal_8509, SubBytesIns_Inst_Sbox_5_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M20_U1 ( .a ({new_AGEMA_signal_8244, new_AGEMA_signal_8243, new_AGEMA_signal_8242, SubBytesIns_Inst_Sbox_5_M16}), .b ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M21_U1 ( .a ({new_AGEMA_signal_8247, new_AGEMA_signal_8246, new_AGEMA_signal_8245, SubBytesIns_Inst_Sbox_5_M17}), .b ({new_AGEMA_signal_8241, new_AGEMA_signal_8240, new_AGEMA_signal_8239, SubBytesIns_Inst_Sbox_5_M15}), .c ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M22_U1 ( .a ({new_AGEMA_signal_8250, new_AGEMA_signal_8249, new_AGEMA_signal_8248, SubBytesIns_Inst_Sbox_5_M18}), .b ({new_AGEMA_signal_7827, new_AGEMA_signal_7826, new_AGEMA_signal_7825, SubBytesIns_Inst_Sbox_5_M13}), .c ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M23_U1 ( .a ({new_AGEMA_signal_8511, new_AGEMA_signal_8510, new_AGEMA_signal_8509, SubBytesIns_Inst_Sbox_5_M19}), .b ({new_AGEMA_signal_7809, new_AGEMA_signal_7808, new_AGEMA_signal_7807, SubBytesIns_Inst_Sbox_5_T25}), .c ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M24_U1 ( .a ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}), .c ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, new_AGEMA_signal_9016, SubBytesIns_Inst_Sbox_5_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M27_U1 ( .a ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}), .c ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_5_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M1_U1 ( .a ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_6_T13}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324]}), .c ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_6_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M2_U1 ( .a ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_6_T23}), .b ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330]}), .c ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, new_AGEMA_signal_7837, SubBytesIns_Inst_Sbox_6_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M3_U1 ( .a ({new_AGEMA_signal_7179, new_AGEMA_signal_7178, new_AGEMA_signal_7177, SubBytesIns_Inst_Sbox_6_T14}), .b ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, new_AGEMA_signal_7840, SubBytesIns_Inst_Sbox_6_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M4_U1 ( .a ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .c ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_6_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M5_U1 ( .a ({new_AGEMA_signal_7197, new_AGEMA_signal_7196, new_AGEMA_signal_7195, SubBytesIns_Inst_Sbox_6_M4}), .b ({new_AGEMA_signal_7194, new_AGEMA_signal_7193, new_AGEMA_signal_7192, SubBytesIns_Inst_Sbox_6_M1}), .c ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, new_AGEMA_signal_7843, SubBytesIns_Inst_Sbox_6_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M6_U1 ( .a ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342]}), .c ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, new_AGEMA_signal_7198, SubBytesIns_Inst_Sbox_6_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M7_U1 ( .a ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348]}), .c ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M8_U1 ( .a ({new_AGEMA_signal_7191, new_AGEMA_signal_7190, new_AGEMA_signal_7189, SubBytesIns_Inst_Sbox_6_T26}), .b ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, new_AGEMA_signal_7198, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, new_AGEMA_signal_7846, SubBytesIns_Inst_Sbox_6_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M9_U1 ( .a ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}), .b ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354]}), .c ({new_AGEMA_signal_7851, new_AGEMA_signal_7850, new_AGEMA_signal_7849, SubBytesIns_Inst_Sbox_6_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M10_U1 ( .a ({new_AGEMA_signal_7851, new_AGEMA_signal_7850, new_AGEMA_signal_7849, SubBytesIns_Inst_Sbox_6_M9}), .b ({new_AGEMA_signal_7200, new_AGEMA_signal_7199, new_AGEMA_signal_7198, SubBytesIns_Inst_Sbox_6_M6}), .c ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M11_U1 ( .a ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .b ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360]}), .c ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_6_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M12_U1 ( .a ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}), .b ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366]}), .c ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_6_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M13_U1 ( .a ({new_AGEMA_signal_7209, new_AGEMA_signal_7208, new_AGEMA_signal_7207, SubBytesIns_Inst_Sbox_6_M12}), .b ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, SubBytesIns_Inst_Sbox_6_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M14_U1 ( .a ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372]}), .c ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, new_AGEMA_signal_7855, SubBytesIns_Inst_Sbox_6_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M15_U1 ( .a ({new_AGEMA_signal_7857, new_AGEMA_signal_7856, new_AGEMA_signal_7855, SubBytesIns_Inst_Sbox_6_M14}), .b ({new_AGEMA_signal_7206, new_AGEMA_signal_7205, new_AGEMA_signal_7204, SubBytesIns_Inst_Sbox_6_M11}), .c ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, new_AGEMA_signal_8254, SubBytesIns_Inst_Sbox_6_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M16_U1 ( .a ({new_AGEMA_signal_7842, new_AGEMA_signal_7841, new_AGEMA_signal_7840, SubBytesIns_Inst_Sbox_6_M3}), .b ({new_AGEMA_signal_7839, new_AGEMA_signal_7838, new_AGEMA_signal_7837, SubBytesIns_Inst_Sbox_6_M2}), .c ({new_AGEMA_signal_8259, new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M17_U1 ( .a ({new_AGEMA_signal_7845, new_AGEMA_signal_7844, new_AGEMA_signal_7843, SubBytesIns_Inst_Sbox_6_M5}), .b ({new_AGEMA_signal_7833, new_AGEMA_signal_7832, new_AGEMA_signal_7831, SubBytesIns_Inst_Sbox_6_T24}), .c ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, new_AGEMA_signal_8260, SubBytesIns_Inst_Sbox_6_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M18_U1 ( .a ({new_AGEMA_signal_7848, new_AGEMA_signal_7847, new_AGEMA_signal_7846, SubBytesIns_Inst_Sbox_6_M8}), .b ({new_AGEMA_signal_7203, new_AGEMA_signal_7202, new_AGEMA_signal_7201, SubBytesIns_Inst_Sbox_6_M7}), .c ({new_AGEMA_signal_8265, new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_6_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M19_U1 ( .a ({new_AGEMA_signal_8253, new_AGEMA_signal_8252, new_AGEMA_signal_8251, SubBytesIns_Inst_Sbox_6_M10}), .b ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, new_AGEMA_signal_8254, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_8523, new_AGEMA_signal_8522, new_AGEMA_signal_8521, SubBytesIns_Inst_Sbox_6_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M20_U1 ( .a ({new_AGEMA_signal_8259, new_AGEMA_signal_8258, new_AGEMA_signal_8257, SubBytesIns_Inst_Sbox_6_M16}), .b ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M21_U1 ( .a ({new_AGEMA_signal_8262, new_AGEMA_signal_8261, new_AGEMA_signal_8260, SubBytesIns_Inst_Sbox_6_M17}), .b ({new_AGEMA_signal_8256, new_AGEMA_signal_8255, new_AGEMA_signal_8254, SubBytesIns_Inst_Sbox_6_M15}), .c ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M22_U1 ( .a ({new_AGEMA_signal_8265, new_AGEMA_signal_8264, new_AGEMA_signal_8263, SubBytesIns_Inst_Sbox_6_M18}), .b ({new_AGEMA_signal_7854, new_AGEMA_signal_7853, new_AGEMA_signal_7852, SubBytesIns_Inst_Sbox_6_M13}), .c ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M23_U1 ( .a ({new_AGEMA_signal_8523, new_AGEMA_signal_8522, new_AGEMA_signal_8521, SubBytesIns_Inst_Sbox_6_M19}), .b ({new_AGEMA_signal_7836, new_AGEMA_signal_7835, new_AGEMA_signal_7834, SubBytesIns_Inst_Sbox_6_T25}), .c ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M24_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}), .c ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, new_AGEMA_signal_9031, SubBytesIns_Inst_Sbox_6_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M27_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}), .c ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_6_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M1_U1 ( .a ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_7_T13}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378]}), .c ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_7_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M2_U1 ( .a ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_7_T23}), .b ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .c ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, new_AGEMA_signal_7864, SubBytesIns_Inst_Sbox_7_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M3_U1 ( .a ({new_AGEMA_signal_7218, new_AGEMA_signal_7217, new_AGEMA_signal_7216, SubBytesIns_Inst_Sbox_7_T14}), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_7869, new_AGEMA_signal_7868, new_AGEMA_signal_7867, SubBytesIns_Inst_Sbox_7_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M4_U1 ( .a ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390]}), .c ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_7_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M5_U1 ( .a ({new_AGEMA_signal_7236, new_AGEMA_signal_7235, new_AGEMA_signal_7234, SubBytesIns_Inst_Sbox_7_M4}), .b ({new_AGEMA_signal_7233, new_AGEMA_signal_7232, new_AGEMA_signal_7231, SubBytesIns_Inst_Sbox_7_M1}), .c ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, new_AGEMA_signal_7870, SubBytesIns_Inst_Sbox_7_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M6_U1 ( .a ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396]}), .c ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_7_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M7_U1 ( .a ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}), .b ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402]}), .c ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_7_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M8_U1 ( .a ({new_AGEMA_signal_7230, new_AGEMA_signal_7229, new_AGEMA_signal_7228, SubBytesIns_Inst_Sbox_7_T26}), .b ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_7_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M9_U1 ( .a ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}), .b ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408]}), .c ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, new_AGEMA_signal_7876, SubBytesIns_Inst_Sbox_7_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M10_U1 ( .a ({new_AGEMA_signal_7878, new_AGEMA_signal_7877, new_AGEMA_signal_7876, SubBytesIns_Inst_Sbox_7_M9}), .b ({new_AGEMA_signal_7239, new_AGEMA_signal_7238, new_AGEMA_signal_7237, SubBytesIns_Inst_Sbox_7_M6}), .c ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, new_AGEMA_signal_8266, SubBytesIns_Inst_Sbox_7_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M11_U1 ( .a ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .b ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414]}), .c ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_7_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M12_U1 ( .a ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}), .b ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420]}), .c ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_7_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M13_U1 ( .a ({new_AGEMA_signal_7248, new_AGEMA_signal_7247, new_AGEMA_signal_7246, SubBytesIns_Inst_Sbox_7_M12}), .b ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_7_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M14_U1 ( .a ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .b ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426]}), .c ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, new_AGEMA_signal_7882, SubBytesIns_Inst_Sbox_7_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M15_U1 ( .a ({new_AGEMA_signal_7884, new_AGEMA_signal_7883, new_AGEMA_signal_7882, SubBytesIns_Inst_Sbox_7_M14}), .b ({new_AGEMA_signal_7245, new_AGEMA_signal_7244, new_AGEMA_signal_7243, SubBytesIns_Inst_Sbox_7_M11}), .c ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M16_U1 ( .a ({new_AGEMA_signal_7869, new_AGEMA_signal_7868, new_AGEMA_signal_7867, SubBytesIns_Inst_Sbox_7_M3}), .b ({new_AGEMA_signal_7866, new_AGEMA_signal_7865, new_AGEMA_signal_7864, SubBytesIns_Inst_Sbox_7_M2}), .c ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, new_AGEMA_signal_8272, SubBytesIns_Inst_Sbox_7_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M17_U1 ( .a ({new_AGEMA_signal_7872, new_AGEMA_signal_7871, new_AGEMA_signal_7870, SubBytesIns_Inst_Sbox_7_M5}), .b ({new_AGEMA_signal_7860, new_AGEMA_signal_7859, new_AGEMA_signal_7858, SubBytesIns_Inst_Sbox_7_T24}), .c ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M18_U1 ( .a ({new_AGEMA_signal_7875, new_AGEMA_signal_7874, new_AGEMA_signal_7873, SubBytesIns_Inst_Sbox_7_M8}), .b ({new_AGEMA_signal_7242, new_AGEMA_signal_7241, new_AGEMA_signal_7240, SubBytesIns_Inst_Sbox_7_M7}), .c ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, new_AGEMA_signal_8278, SubBytesIns_Inst_Sbox_7_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M19_U1 ( .a ({new_AGEMA_signal_8268, new_AGEMA_signal_8267, new_AGEMA_signal_8266, SubBytesIns_Inst_Sbox_7_M10}), .b ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_8535, new_AGEMA_signal_8534, new_AGEMA_signal_8533, SubBytesIns_Inst_Sbox_7_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M20_U1 ( .a ({new_AGEMA_signal_8274, new_AGEMA_signal_8273, new_AGEMA_signal_8272, SubBytesIns_Inst_Sbox_7_M16}), .b ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M21_U1 ( .a ({new_AGEMA_signal_8277, new_AGEMA_signal_8276, new_AGEMA_signal_8275, SubBytesIns_Inst_Sbox_7_M17}), .b ({new_AGEMA_signal_8271, new_AGEMA_signal_8270, new_AGEMA_signal_8269, SubBytesIns_Inst_Sbox_7_M15}), .c ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M22_U1 ( .a ({new_AGEMA_signal_8280, new_AGEMA_signal_8279, new_AGEMA_signal_8278, SubBytesIns_Inst_Sbox_7_M18}), .b ({new_AGEMA_signal_7881, new_AGEMA_signal_7880, new_AGEMA_signal_7879, SubBytesIns_Inst_Sbox_7_M13}), .c ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M23_U1 ( .a ({new_AGEMA_signal_8535, new_AGEMA_signal_8534, new_AGEMA_signal_8533, SubBytesIns_Inst_Sbox_7_M19}), .b ({new_AGEMA_signal_7863, new_AGEMA_signal_7862, new_AGEMA_signal_7861, SubBytesIns_Inst_Sbox_7_T25}), .c ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M24_U1 ( .a ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}), .c ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, new_AGEMA_signal_9046, SubBytesIns_Inst_Sbox_7_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M27_U1 ( .a ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}), .c ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_7_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M1_U1 ( .a ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_8_T13}), .b ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .c ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M2_U1 ( .a ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, SubBytesIns_Inst_Sbox_8_T23}), .b ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438]}), .c ({new_AGEMA_signal_7893, new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_8_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M3_U1 ( .a ({new_AGEMA_signal_7257, new_AGEMA_signal_7256, new_AGEMA_signal_7255, SubBytesIns_Inst_Sbox_8_T14}), .b ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, new_AGEMA_signal_7894, SubBytesIns_Inst_Sbox_8_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M4_U1 ( .a ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444]}), .c ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M5_U1 ( .a ({new_AGEMA_signal_7275, new_AGEMA_signal_7274, new_AGEMA_signal_7273, SubBytesIns_Inst_Sbox_8_M4}), .b ({new_AGEMA_signal_7272, new_AGEMA_signal_7271, new_AGEMA_signal_7270, SubBytesIns_Inst_Sbox_8_M1}), .c ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_8_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M6_U1 ( .a ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450]}), .c ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_8_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M7_U1 ( .a ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}), .b ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456]}), .c ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_8_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M8_U1 ( .a ({new_AGEMA_signal_7269, new_AGEMA_signal_7268, new_AGEMA_signal_7267, SubBytesIns_Inst_Sbox_8_T26}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, new_AGEMA_signal_7900, SubBytesIns_Inst_Sbox_8_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M9_U1 ( .a ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462]}), .c ({new_AGEMA_signal_7905, new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_8_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M10_U1 ( .a ({new_AGEMA_signal_7905, new_AGEMA_signal_7904, new_AGEMA_signal_7903, SubBytesIns_Inst_Sbox_8_M9}), .b ({new_AGEMA_signal_7278, new_AGEMA_signal_7277, new_AGEMA_signal_7276, SubBytesIns_Inst_Sbox_8_M6}), .c ({new_AGEMA_signal_8283, new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_8_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M11_U1 ( .a ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .b ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468]}), .c ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_8_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M12_U1 ( .a ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}), .b ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474]}), .c ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_8_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M13_U1 ( .a ({new_AGEMA_signal_7287, new_AGEMA_signal_7286, new_AGEMA_signal_7285, SubBytesIns_Inst_Sbox_8_M12}), .b ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, SubBytesIns_Inst_Sbox_8_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M14_U1 ( .a ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .b ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .c ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_8_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M15_U1 ( .a ({new_AGEMA_signal_7911, new_AGEMA_signal_7910, new_AGEMA_signal_7909, SubBytesIns_Inst_Sbox_8_M14}), .b ({new_AGEMA_signal_7284, new_AGEMA_signal_7283, new_AGEMA_signal_7282, SubBytesIns_Inst_Sbox_8_M11}), .c ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, new_AGEMA_signal_8284, SubBytesIns_Inst_Sbox_8_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M16_U1 ( .a ({new_AGEMA_signal_7896, new_AGEMA_signal_7895, new_AGEMA_signal_7894, SubBytesIns_Inst_Sbox_8_M3}), .b ({new_AGEMA_signal_7893, new_AGEMA_signal_7892, new_AGEMA_signal_7891, SubBytesIns_Inst_Sbox_8_M2}), .c ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M17_U1 ( .a ({new_AGEMA_signal_7899, new_AGEMA_signal_7898, new_AGEMA_signal_7897, SubBytesIns_Inst_Sbox_8_M5}), .b ({new_AGEMA_signal_7887, new_AGEMA_signal_7886, new_AGEMA_signal_7885, SubBytesIns_Inst_Sbox_8_T24}), .c ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, new_AGEMA_signal_8290, SubBytesIns_Inst_Sbox_8_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M18_U1 ( .a ({new_AGEMA_signal_7902, new_AGEMA_signal_7901, new_AGEMA_signal_7900, SubBytesIns_Inst_Sbox_8_M8}), .b ({new_AGEMA_signal_7281, new_AGEMA_signal_7280, new_AGEMA_signal_7279, SubBytesIns_Inst_Sbox_8_M7}), .c ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M19_U1 ( .a ({new_AGEMA_signal_8283, new_AGEMA_signal_8282, new_AGEMA_signal_8281, SubBytesIns_Inst_Sbox_8_M10}), .b ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, new_AGEMA_signal_8284, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_8547, new_AGEMA_signal_8546, new_AGEMA_signal_8545, SubBytesIns_Inst_Sbox_8_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M20_U1 ( .a ({new_AGEMA_signal_8289, new_AGEMA_signal_8288, new_AGEMA_signal_8287, SubBytesIns_Inst_Sbox_8_M16}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M21_U1 ( .a ({new_AGEMA_signal_8292, new_AGEMA_signal_8291, new_AGEMA_signal_8290, SubBytesIns_Inst_Sbox_8_M17}), .b ({new_AGEMA_signal_8286, new_AGEMA_signal_8285, new_AGEMA_signal_8284, SubBytesIns_Inst_Sbox_8_M15}), .c ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M22_U1 ( .a ({new_AGEMA_signal_8295, new_AGEMA_signal_8294, new_AGEMA_signal_8293, SubBytesIns_Inst_Sbox_8_M18}), .b ({new_AGEMA_signal_7908, new_AGEMA_signal_7907, new_AGEMA_signal_7906, SubBytesIns_Inst_Sbox_8_M13}), .c ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M23_U1 ( .a ({new_AGEMA_signal_8547, new_AGEMA_signal_8546, new_AGEMA_signal_8545, SubBytesIns_Inst_Sbox_8_M19}), .b ({new_AGEMA_signal_7890, new_AGEMA_signal_7889, new_AGEMA_signal_7888, SubBytesIns_Inst_Sbox_8_T25}), .c ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M24_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}), .c ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_8_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M27_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}), .c ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_8_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M1_U1 ( .a ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_9_T13}), .b ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486]}), .c ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_9_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M2_U1 ( .a ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_9_T23}), .b ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492]}), .c ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, new_AGEMA_signal_7918, SubBytesIns_Inst_Sbox_9_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M3_U1 ( .a ({new_AGEMA_signal_7296, new_AGEMA_signal_7295, new_AGEMA_signal_7294, SubBytesIns_Inst_Sbox_9_T14}), .b ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_9_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M4_U1 ( .a ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498]}), .c ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_9_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M5_U1 ( .a ({new_AGEMA_signal_7314, new_AGEMA_signal_7313, new_AGEMA_signal_7312, SubBytesIns_Inst_Sbox_9_M4}), .b ({new_AGEMA_signal_7311, new_AGEMA_signal_7310, new_AGEMA_signal_7309, SubBytesIns_Inst_Sbox_9_M1}), .c ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, new_AGEMA_signal_7924, SubBytesIns_Inst_Sbox_9_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M6_U1 ( .a ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504]}), .c ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_9_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M7_U1 ( .a ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}), .b ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510]}), .c ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_9_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M8_U1 ( .a ({new_AGEMA_signal_7308, new_AGEMA_signal_7307, new_AGEMA_signal_7306, SubBytesIns_Inst_Sbox_9_T26}), .b ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_9_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M9_U1 ( .a ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516]}), .c ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, new_AGEMA_signal_7930, SubBytesIns_Inst_Sbox_9_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M10_U1 ( .a ({new_AGEMA_signal_7932, new_AGEMA_signal_7931, new_AGEMA_signal_7930, SubBytesIns_Inst_Sbox_9_M9}), .b ({new_AGEMA_signal_7317, new_AGEMA_signal_7316, new_AGEMA_signal_7315, SubBytesIns_Inst_Sbox_9_M6}), .c ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, new_AGEMA_signal_8296, SubBytesIns_Inst_Sbox_9_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M11_U1 ( .a ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .b ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522]}), .c ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_9_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M12_U1 ( .a ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}), .b ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .c ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_9_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M13_U1 ( .a ({new_AGEMA_signal_7326, new_AGEMA_signal_7325, new_AGEMA_signal_7324, SubBytesIns_Inst_Sbox_9_M12}), .b ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_9_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M14_U1 ( .a ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .b ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534]}), .c ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, new_AGEMA_signal_7936, SubBytesIns_Inst_Sbox_9_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M15_U1 ( .a ({new_AGEMA_signal_7938, new_AGEMA_signal_7937, new_AGEMA_signal_7936, SubBytesIns_Inst_Sbox_9_M14}), .b ({new_AGEMA_signal_7323, new_AGEMA_signal_7322, new_AGEMA_signal_7321, SubBytesIns_Inst_Sbox_9_M11}), .c ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_9_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M16_U1 ( .a ({new_AGEMA_signal_7923, new_AGEMA_signal_7922, new_AGEMA_signal_7921, SubBytesIns_Inst_Sbox_9_M3}), .b ({new_AGEMA_signal_7920, new_AGEMA_signal_7919, new_AGEMA_signal_7918, SubBytesIns_Inst_Sbox_9_M2}), .c ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, new_AGEMA_signal_8302, SubBytesIns_Inst_Sbox_9_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M17_U1 ( .a ({new_AGEMA_signal_7926, new_AGEMA_signal_7925, new_AGEMA_signal_7924, SubBytesIns_Inst_Sbox_9_M5}), .b ({new_AGEMA_signal_7914, new_AGEMA_signal_7913, new_AGEMA_signal_7912, SubBytesIns_Inst_Sbox_9_T24}), .c ({new_AGEMA_signal_8307, new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_9_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M18_U1 ( .a ({new_AGEMA_signal_7929, new_AGEMA_signal_7928, new_AGEMA_signal_7927, SubBytesIns_Inst_Sbox_9_M8}), .b ({new_AGEMA_signal_7320, new_AGEMA_signal_7319, new_AGEMA_signal_7318, SubBytesIns_Inst_Sbox_9_M7}), .c ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, new_AGEMA_signal_8308, SubBytesIns_Inst_Sbox_9_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M19_U1 ( .a ({new_AGEMA_signal_8298, new_AGEMA_signal_8297, new_AGEMA_signal_8296, SubBytesIns_Inst_Sbox_9_M10}), .b ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, new_AGEMA_signal_8557, SubBytesIns_Inst_Sbox_9_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M20_U1 ( .a ({new_AGEMA_signal_8304, new_AGEMA_signal_8303, new_AGEMA_signal_8302, SubBytesIns_Inst_Sbox_9_M16}), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M21_U1 ( .a ({new_AGEMA_signal_8307, new_AGEMA_signal_8306, new_AGEMA_signal_8305, SubBytesIns_Inst_Sbox_9_M17}), .b ({new_AGEMA_signal_8301, new_AGEMA_signal_8300, new_AGEMA_signal_8299, SubBytesIns_Inst_Sbox_9_M15}), .c ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M22_U1 ( .a ({new_AGEMA_signal_8310, new_AGEMA_signal_8309, new_AGEMA_signal_8308, SubBytesIns_Inst_Sbox_9_M18}), .b ({new_AGEMA_signal_7935, new_AGEMA_signal_7934, new_AGEMA_signal_7933, SubBytesIns_Inst_Sbox_9_M13}), .c ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M23_U1 ( .a ({new_AGEMA_signal_8559, new_AGEMA_signal_8558, new_AGEMA_signal_8557, SubBytesIns_Inst_Sbox_9_M19}), .b ({new_AGEMA_signal_7917, new_AGEMA_signal_7916, new_AGEMA_signal_7915, SubBytesIns_Inst_Sbox_9_T25}), .c ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M24_U1 ( .a ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}), .c ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, new_AGEMA_signal_9076, SubBytesIns_Inst_Sbox_9_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M27_U1 ( .a ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}), .c ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M1_U1 ( .a ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_10_T13}), .b ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540]}), .c ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_10_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M2_U1 ( .a ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_10_T23}), .b ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546]}), .c ({new_AGEMA_signal_7947, new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_10_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M3_U1 ( .a ({new_AGEMA_signal_7335, new_AGEMA_signal_7334, new_AGEMA_signal_7333, SubBytesIns_Inst_Sbox_10_T14}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, new_AGEMA_signal_7948, SubBytesIns_Inst_Sbox_10_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M4_U1 ( .a ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552]}), .c ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_10_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M5_U1 ( .a ({new_AGEMA_signal_7353, new_AGEMA_signal_7352, new_AGEMA_signal_7351, SubBytesIns_Inst_Sbox_10_M4}), .b ({new_AGEMA_signal_7350, new_AGEMA_signal_7349, new_AGEMA_signal_7348, SubBytesIns_Inst_Sbox_10_M1}), .c ({new_AGEMA_signal_7953, new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M6_U1 ( .a ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558]}), .c ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, SubBytesIns_Inst_Sbox_10_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M7_U1 ( .a ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}), .b ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564]}), .c ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_10_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M8_U1 ( .a ({new_AGEMA_signal_7347, new_AGEMA_signal_7346, new_AGEMA_signal_7345, SubBytesIns_Inst_Sbox_10_T26}), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, new_AGEMA_signal_7954, SubBytesIns_Inst_Sbox_10_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M9_U1 ( .a ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570]}), .c ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_10_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M10_U1 ( .a ({new_AGEMA_signal_7959, new_AGEMA_signal_7958, new_AGEMA_signal_7957, SubBytesIns_Inst_Sbox_10_M9}), .b ({new_AGEMA_signal_7356, new_AGEMA_signal_7355, new_AGEMA_signal_7354, SubBytesIns_Inst_Sbox_10_M6}), .c ({new_AGEMA_signal_8313, new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_10_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M11_U1 ( .a ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .b ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .c ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, SubBytesIns_Inst_Sbox_10_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M12_U1 ( .a ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}), .b ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582]}), .c ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_10_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M13_U1 ( .a ({new_AGEMA_signal_7365, new_AGEMA_signal_7364, new_AGEMA_signal_7363, SubBytesIns_Inst_Sbox_10_M12}), .b ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, SubBytesIns_Inst_Sbox_10_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M14_U1 ( .a ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588]}), .c ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_10_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M15_U1 ( .a ({new_AGEMA_signal_7965, new_AGEMA_signal_7964, new_AGEMA_signal_7963, SubBytesIns_Inst_Sbox_10_M14}), .b ({new_AGEMA_signal_7362, new_AGEMA_signal_7361, new_AGEMA_signal_7360, SubBytesIns_Inst_Sbox_10_M11}), .c ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, new_AGEMA_signal_8314, SubBytesIns_Inst_Sbox_10_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M16_U1 ( .a ({new_AGEMA_signal_7950, new_AGEMA_signal_7949, new_AGEMA_signal_7948, SubBytesIns_Inst_Sbox_10_M3}), .b ({new_AGEMA_signal_7947, new_AGEMA_signal_7946, new_AGEMA_signal_7945, SubBytesIns_Inst_Sbox_10_M2}), .c ({new_AGEMA_signal_8319, new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_10_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M17_U1 ( .a ({new_AGEMA_signal_7953, new_AGEMA_signal_7952, new_AGEMA_signal_7951, SubBytesIns_Inst_Sbox_10_M5}), .b ({new_AGEMA_signal_7941, new_AGEMA_signal_7940, new_AGEMA_signal_7939, SubBytesIns_Inst_Sbox_10_T24}), .c ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, new_AGEMA_signal_8320, SubBytesIns_Inst_Sbox_10_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M18_U1 ( .a ({new_AGEMA_signal_7956, new_AGEMA_signal_7955, new_AGEMA_signal_7954, SubBytesIns_Inst_Sbox_10_M8}), .b ({new_AGEMA_signal_7359, new_AGEMA_signal_7358, new_AGEMA_signal_7357, SubBytesIns_Inst_Sbox_10_M7}), .c ({new_AGEMA_signal_8325, new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_10_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M19_U1 ( .a ({new_AGEMA_signal_8313, new_AGEMA_signal_8312, new_AGEMA_signal_8311, SubBytesIns_Inst_Sbox_10_M10}), .b ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, new_AGEMA_signal_8314, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_8571, new_AGEMA_signal_8570, new_AGEMA_signal_8569, SubBytesIns_Inst_Sbox_10_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M20_U1 ( .a ({new_AGEMA_signal_8319, new_AGEMA_signal_8318, new_AGEMA_signal_8317, SubBytesIns_Inst_Sbox_10_M16}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M21_U1 ( .a ({new_AGEMA_signal_8322, new_AGEMA_signal_8321, new_AGEMA_signal_8320, SubBytesIns_Inst_Sbox_10_M17}), .b ({new_AGEMA_signal_8316, new_AGEMA_signal_8315, new_AGEMA_signal_8314, SubBytesIns_Inst_Sbox_10_M15}), .c ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M22_U1 ( .a ({new_AGEMA_signal_8325, new_AGEMA_signal_8324, new_AGEMA_signal_8323, SubBytesIns_Inst_Sbox_10_M18}), .b ({new_AGEMA_signal_7962, new_AGEMA_signal_7961, new_AGEMA_signal_7960, SubBytesIns_Inst_Sbox_10_M13}), .c ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M23_U1 ( .a ({new_AGEMA_signal_8571, new_AGEMA_signal_8570, new_AGEMA_signal_8569, SubBytesIns_Inst_Sbox_10_M19}), .b ({new_AGEMA_signal_7944, new_AGEMA_signal_7943, new_AGEMA_signal_7942, SubBytesIns_Inst_Sbox_10_T25}), .c ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M24_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}), .c ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_10_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M27_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}), .c ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M1_U1 ( .a ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_11_T13}), .b ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594]}), .c ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_11_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M2_U1 ( .a ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_11_T23}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600]}), .c ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, new_AGEMA_signal_7972, SubBytesIns_Inst_Sbox_11_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M3_U1 ( .a ({new_AGEMA_signal_7374, new_AGEMA_signal_7373, new_AGEMA_signal_7372, SubBytesIns_Inst_Sbox_11_T14}), .b ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_11_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M4_U1 ( .a ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606]}), .c ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, new_AGEMA_signal_7390, SubBytesIns_Inst_Sbox_11_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M5_U1 ( .a ({new_AGEMA_signal_7392, new_AGEMA_signal_7391, new_AGEMA_signal_7390, SubBytesIns_Inst_Sbox_11_M4}), .b ({new_AGEMA_signal_7389, new_AGEMA_signal_7388, new_AGEMA_signal_7387, SubBytesIns_Inst_Sbox_11_M1}), .c ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, new_AGEMA_signal_7978, SubBytesIns_Inst_Sbox_11_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M6_U1 ( .a ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612]}), .c ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_11_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M7_U1 ( .a ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}), .b ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618]}), .c ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, new_AGEMA_signal_7396, SubBytesIns_Inst_Sbox_11_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M8_U1 ( .a ({new_AGEMA_signal_7386, new_AGEMA_signal_7385, new_AGEMA_signal_7384, SubBytesIns_Inst_Sbox_11_T26}), .b ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_7983, new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_11_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M9_U1 ( .a ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .c ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, new_AGEMA_signal_7984, SubBytesIns_Inst_Sbox_11_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M10_U1 ( .a ({new_AGEMA_signal_7986, new_AGEMA_signal_7985, new_AGEMA_signal_7984, SubBytesIns_Inst_Sbox_11_M9}), .b ({new_AGEMA_signal_7395, new_AGEMA_signal_7394, new_AGEMA_signal_7393, SubBytesIns_Inst_Sbox_11_M6}), .c ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, new_AGEMA_signal_8326, SubBytesIns_Inst_Sbox_11_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M11_U1 ( .a ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .b ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630]}), .c ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M12_U1 ( .a ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}), .b ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636]}), .c ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, new_AGEMA_signal_7402, SubBytesIns_Inst_Sbox_11_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M13_U1 ( .a ({new_AGEMA_signal_7404, new_AGEMA_signal_7403, new_AGEMA_signal_7402, SubBytesIns_Inst_Sbox_11_M12}), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_11_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M14_U1 ( .a ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642]}), .c ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, new_AGEMA_signal_7990, SubBytesIns_Inst_Sbox_11_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M15_U1 ( .a ({new_AGEMA_signal_7992, new_AGEMA_signal_7991, new_AGEMA_signal_7990, SubBytesIns_Inst_Sbox_11_M14}), .b ({new_AGEMA_signal_7401, new_AGEMA_signal_7400, new_AGEMA_signal_7399, SubBytesIns_Inst_Sbox_11_M11}), .c ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_11_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M16_U1 ( .a ({new_AGEMA_signal_7977, new_AGEMA_signal_7976, new_AGEMA_signal_7975, SubBytesIns_Inst_Sbox_11_M3}), .b ({new_AGEMA_signal_7974, new_AGEMA_signal_7973, new_AGEMA_signal_7972, SubBytesIns_Inst_Sbox_11_M2}), .c ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, new_AGEMA_signal_8332, SubBytesIns_Inst_Sbox_11_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M17_U1 ( .a ({new_AGEMA_signal_7980, new_AGEMA_signal_7979, new_AGEMA_signal_7978, SubBytesIns_Inst_Sbox_11_M5}), .b ({new_AGEMA_signal_7968, new_AGEMA_signal_7967, new_AGEMA_signal_7966, SubBytesIns_Inst_Sbox_11_T24}), .c ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_11_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M18_U1 ( .a ({new_AGEMA_signal_7983, new_AGEMA_signal_7982, new_AGEMA_signal_7981, SubBytesIns_Inst_Sbox_11_M8}), .b ({new_AGEMA_signal_7398, new_AGEMA_signal_7397, new_AGEMA_signal_7396, SubBytesIns_Inst_Sbox_11_M7}), .c ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, new_AGEMA_signal_8338, SubBytesIns_Inst_Sbox_11_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M19_U1 ( .a ({new_AGEMA_signal_8328, new_AGEMA_signal_8327, new_AGEMA_signal_8326, SubBytesIns_Inst_Sbox_11_M10}), .b ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_8583, new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_11_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M20_U1 ( .a ({new_AGEMA_signal_8334, new_AGEMA_signal_8333, new_AGEMA_signal_8332, SubBytesIns_Inst_Sbox_11_M16}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M21_U1 ( .a ({new_AGEMA_signal_8337, new_AGEMA_signal_8336, new_AGEMA_signal_8335, SubBytesIns_Inst_Sbox_11_M17}), .b ({new_AGEMA_signal_8331, new_AGEMA_signal_8330, new_AGEMA_signal_8329, SubBytesIns_Inst_Sbox_11_M15}), .c ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M22_U1 ( .a ({new_AGEMA_signal_8340, new_AGEMA_signal_8339, new_AGEMA_signal_8338, SubBytesIns_Inst_Sbox_11_M18}), .b ({new_AGEMA_signal_7989, new_AGEMA_signal_7988, new_AGEMA_signal_7987, SubBytesIns_Inst_Sbox_11_M13}), .c ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M23_U1 ( .a ({new_AGEMA_signal_8583, new_AGEMA_signal_8582, new_AGEMA_signal_8581, SubBytesIns_Inst_Sbox_11_M19}), .b ({new_AGEMA_signal_7971, new_AGEMA_signal_7970, new_AGEMA_signal_7969, SubBytesIns_Inst_Sbox_11_T25}), .c ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M24_U1 ( .a ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}), .c ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, new_AGEMA_signal_9106, SubBytesIns_Inst_Sbox_11_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M27_U1 ( .a ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}), .c ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_11_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M1_U1 ( .a ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_12_T13}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648]}), .c ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, SubBytesIns_Inst_Sbox_12_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M2_U1 ( .a ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, SubBytesIns_Inst_Sbox_12_T23}), .b ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654]}), .c ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, new_AGEMA_signal_7999, SubBytesIns_Inst_Sbox_12_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M3_U1 ( .a ({new_AGEMA_signal_7413, new_AGEMA_signal_7412, new_AGEMA_signal_7411, SubBytesIns_Inst_Sbox_12_T14}), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, new_AGEMA_signal_8002, SubBytesIns_Inst_Sbox_12_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M4_U1 ( .a ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660]}), .c ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_12_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M5_U1 ( .a ({new_AGEMA_signal_7431, new_AGEMA_signal_7430, new_AGEMA_signal_7429, SubBytesIns_Inst_Sbox_12_M4}), .b ({new_AGEMA_signal_7428, new_AGEMA_signal_7427, new_AGEMA_signal_7426, SubBytesIns_Inst_Sbox_12_M1}), .c ({new_AGEMA_signal_8007, new_AGEMA_signal_8006, new_AGEMA_signal_8005, SubBytesIns_Inst_Sbox_12_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M6_U1 ( .a ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666]}), .c ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, SubBytesIns_Inst_Sbox_12_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M7_U1 ( .a ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}), .b ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .c ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_12_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M8_U1 ( .a ({new_AGEMA_signal_7425, new_AGEMA_signal_7424, new_AGEMA_signal_7423, SubBytesIns_Inst_Sbox_12_T26}), .b ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, new_AGEMA_signal_8008, SubBytesIns_Inst_Sbox_12_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M9_U1 ( .a ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678]}), .c ({new_AGEMA_signal_8013, new_AGEMA_signal_8012, new_AGEMA_signal_8011, SubBytesIns_Inst_Sbox_12_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M10_U1 ( .a ({new_AGEMA_signal_8013, new_AGEMA_signal_8012, new_AGEMA_signal_8011, SubBytesIns_Inst_Sbox_12_M9}), .b ({new_AGEMA_signal_7434, new_AGEMA_signal_7433, new_AGEMA_signal_7432, SubBytesIns_Inst_Sbox_12_M6}), .c ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_12_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M11_U1 ( .a ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .b ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684]}), .c ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, SubBytesIns_Inst_Sbox_12_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M12_U1 ( .a ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}), .b ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690]}), .c ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, new_AGEMA_signal_7441, SubBytesIns_Inst_Sbox_12_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M13_U1 ( .a ({new_AGEMA_signal_7443, new_AGEMA_signal_7442, new_AGEMA_signal_7441, SubBytesIns_Inst_Sbox_12_M12}), .b ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, SubBytesIns_Inst_Sbox_12_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M14_U1 ( .a ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696]}), .c ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, new_AGEMA_signal_8017, SubBytesIns_Inst_Sbox_12_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M15_U1 ( .a ({new_AGEMA_signal_8019, new_AGEMA_signal_8018, new_AGEMA_signal_8017, SubBytesIns_Inst_Sbox_12_M14}), .b ({new_AGEMA_signal_7440, new_AGEMA_signal_7439, new_AGEMA_signal_7438, SubBytesIns_Inst_Sbox_12_M11}), .c ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, new_AGEMA_signal_8344, SubBytesIns_Inst_Sbox_12_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M16_U1 ( .a ({new_AGEMA_signal_8004, new_AGEMA_signal_8003, new_AGEMA_signal_8002, SubBytesIns_Inst_Sbox_12_M3}), .b ({new_AGEMA_signal_8001, new_AGEMA_signal_8000, new_AGEMA_signal_7999, SubBytesIns_Inst_Sbox_12_M2}), .c ({new_AGEMA_signal_8349, new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_12_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M17_U1 ( .a ({new_AGEMA_signal_8007, new_AGEMA_signal_8006, new_AGEMA_signal_8005, SubBytesIns_Inst_Sbox_12_M5}), .b ({new_AGEMA_signal_7995, new_AGEMA_signal_7994, new_AGEMA_signal_7993, SubBytesIns_Inst_Sbox_12_T24}), .c ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, new_AGEMA_signal_8350, SubBytesIns_Inst_Sbox_12_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M18_U1 ( .a ({new_AGEMA_signal_8010, new_AGEMA_signal_8009, new_AGEMA_signal_8008, SubBytesIns_Inst_Sbox_12_M8}), .b ({new_AGEMA_signal_7437, new_AGEMA_signal_7436, new_AGEMA_signal_7435, SubBytesIns_Inst_Sbox_12_M7}), .c ({new_AGEMA_signal_8355, new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_12_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M19_U1 ( .a ({new_AGEMA_signal_8343, new_AGEMA_signal_8342, new_AGEMA_signal_8341, SubBytesIns_Inst_Sbox_12_M10}), .b ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, new_AGEMA_signal_8344, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_8595, new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_12_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M20_U1 ( .a ({new_AGEMA_signal_8349, new_AGEMA_signal_8348, new_AGEMA_signal_8347, SubBytesIns_Inst_Sbox_12_M16}), .b ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M21_U1 ( .a ({new_AGEMA_signal_8352, new_AGEMA_signal_8351, new_AGEMA_signal_8350, SubBytesIns_Inst_Sbox_12_M17}), .b ({new_AGEMA_signal_8346, new_AGEMA_signal_8345, new_AGEMA_signal_8344, SubBytesIns_Inst_Sbox_12_M15}), .c ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M22_U1 ( .a ({new_AGEMA_signal_8355, new_AGEMA_signal_8354, new_AGEMA_signal_8353, SubBytesIns_Inst_Sbox_12_M18}), .b ({new_AGEMA_signal_8016, new_AGEMA_signal_8015, new_AGEMA_signal_8014, SubBytesIns_Inst_Sbox_12_M13}), .c ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M23_U1 ( .a ({new_AGEMA_signal_8595, new_AGEMA_signal_8594, new_AGEMA_signal_8593, SubBytesIns_Inst_Sbox_12_M19}), .b ({new_AGEMA_signal_7998, new_AGEMA_signal_7997, new_AGEMA_signal_7996, SubBytesIns_Inst_Sbox_12_T25}), .c ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M24_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}), .c ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_12_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M27_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}), .c ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_12_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M1_U1 ( .a ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_13_T13}), .b ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702]}), .c ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, SubBytesIns_Inst_Sbox_13_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M2_U1 ( .a ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, SubBytesIns_Inst_Sbox_13_T23}), .b ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708]}), .c ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, new_AGEMA_signal_8026, SubBytesIns_Inst_Sbox_13_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M3_U1 ( .a ({new_AGEMA_signal_7452, new_AGEMA_signal_7451, new_AGEMA_signal_7450, SubBytesIns_Inst_Sbox_13_T14}), .b ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, new_AGEMA_signal_8029, SubBytesIns_Inst_Sbox_13_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M4_U1 ( .a ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714]}), .c ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, new_AGEMA_signal_7468, SubBytesIns_Inst_Sbox_13_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M5_U1 ( .a ({new_AGEMA_signal_7470, new_AGEMA_signal_7469, new_AGEMA_signal_7468, SubBytesIns_Inst_Sbox_13_M4}), .b ({new_AGEMA_signal_7467, new_AGEMA_signal_7466, new_AGEMA_signal_7465, SubBytesIns_Inst_Sbox_13_M1}), .c ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, new_AGEMA_signal_8032, SubBytesIns_Inst_Sbox_13_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M6_U1 ( .a ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .c ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, SubBytesIns_Inst_Sbox_13_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M7_U1 ( .a ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}), .b ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726]}), .c ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, new_AGEMA_signal_7474, SubBytesIns_Inst_Sbox_13_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M8_U1 ( .a ({new_AGEMA_signal_7464, new_AGEMA_signal_7463, new_AGEMA_signal_7462, SubBytesIns_Inst_Sbox_13_T26}), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_8037, new_AGEMA_signal_8036, new_AGEMA_signal_8035, SubBytesIns_Inst_Sbox_13_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M9_U1 ( .a ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}), .b ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732]}), .c ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, new_AGEMA_signal_8038, SubBytesIns_Inst_Sbox_13_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M10_U1 ( .a ({new_AGEMA_signal_8040, new_AGEMA_signal_8039, new_AGEMA_signal_8038, SubBytesIns_Inst_Sbox_13_M9}), .b ({new_AGEMA_signal_7473, new_AGEMA_signal_7472, new_AGEMA_signal_7471, SubBytesIns_Inst_Sbox_13_M6}), .c ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, new_AGEMA_signal_8356, SubBytesIns_Inst_Sbox_13_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M11_U1 ( .a ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .b ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738]}), .c ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_13_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M12_U1 ( .a ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}), .b ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744]}), .c ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, new_AGEMA_signal_7480, SubBytesIns_Inst_Sbox_13_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M13_U1 ( .a ({new_AGEMA_signal_7482, new_AGEMA_signal_7481, new_AGEMA_signal_7480, SubBytesIns_Inst_Sbox_13_M12}), .b ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, new_AGEMA_signal_8041, SubBytesIns_Inst_Sbox_13_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M14_U1 ( .a ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750]}), .c ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, new_AGEMA_signal_8044, SubBytesIns_Inst_Sbox_13_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M15_U1 ( .a ({new_AGEMA_signal_8046, new_AGEMA_signal_8045, new_AGEMA_signal_8044, SubBytesIns_Inst_Sbox_13_M14}), .b ({new_AGEMA_signal_7479, new_AGEMA_signal_7478, new_AGEMA_signal_7477, SubBytesIns_Inst_Sbox_13_M11}), .c ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_13_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M16_U1 ( .a ({new_AGEMA_signal_8031, new_AGEMA_signal_8030, new_AGEMA_signal_8029, SubBytesIns_Inst_Sbox_13_M3}), .b ({new_AGEMA_signal_8028, new_AGEMA_signal_8027, new_AGEMA_signal_8026, SubBytesIns_Inst_Sbox_13_M2}), .c ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, new_AGEMA_signal_8362, SubBytesIns_Inst_Sbox_13_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M17_U1 ( .a ({new_AGEMA_signal_8034, new_AGEMA_signal_8033, new_AGEMA_signal_8032, SubBytesIns_Inst_Sbox_13_M5}), .b ({new_AGEMA_signal_8022, new_AGEMA_signal_8021, new_AGEMA_signal_8020, SubBytesIns_Inst_Sbox_13_T24}), .c ({new_AGEMA_signal_8367, new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_13_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M18_U1 ( .a ({new_AGEMA_signal_8037, new_AGEMA_signal_8036, new_AGEMA_signal_8035, SubBytesIns_Inst_Sbox_13_M8}), .b ({new_AGEMA_signal_7476, new_AGEMA_signal_7475, new_AGEMA_signal_7474, SubBytesIns_Inst_Sbox_13_M7}), .c ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, new_AGEMA_signal_8368, SubBytesIns_Inst_Sbox_13_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M19_U1 ( .a ({new_AGEMA_signal_8358, new_AGEMA_signal_8357, new_AGEMA_signal_8356, SubBytesIns_Inst_Sbox_13_M10}), .b ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_13_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M20_U1 ( .a ({new_AGEMA_signal_8364, new_AGEMA_signal_8363, new_AGEMA_signal_8362, SubBytesIns_Inst_Sbox_13_M16}), .b ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, new_AGEMA_signal_8041, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M21_U1 ( .a ({new_AGEMA_signal_8367, new_AGEMA_signal_8366, new_AGEMA_signal_8365, SubBytesIns_Inst_Sbox_13_M17}), .b ({new_AGEMA_signal_8361, new_AGEMA_signal_8360, new_AGEMA_signal_8359, SubBytesIns_Inst_Sbox_13_M15}), .c ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M22_U1 ( .a ({new_AGEMA_signal_8370, new_AGEMA_signal_8369, new_AGEMA_signal_8368, SubBytesIns_Inst_Sbox_13_M18}), .b ({new_AGEMA_signal_8043, new_AGEMA_signal_8042, new_AGEMA_signal_8041, SubBytesIns_Inst_Sbox_13_M13}), .c ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M23_U1 ( .a ({new_AGEMA_signal_8607, new_AGEMA_signal_8606, new_AGEMA_signal_8605, SubBytesIns_Inst_Sbox_13_M19}), .b ({new_AGEMA_signal_8025, new_AGEMA_signal_8024, new_AGEMA_signal_8023, SubBytesIns_Inst_Sbox_13_T25}), .c ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M24_U1 ( .a ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}), .c ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, new_AGEMA_signal_9136, SubBytesIns_Inst_Sbox_13_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M27_U1 ( .a ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}), .c ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_13_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M1_U1 ( .a ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_T13}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756]}), .c ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, SubBytesIns_Inst_Sbox_14_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M2_U1 ( .a ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, SubBytesIns_Inst_Sbox_14_T23}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762]}), .c ({new_AGEMA_signal_8055, new_AGEMA_signal_8054, new_AGEMA_signal_8053, SubBytesIns_Inst_Sbox_14_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M3_U1 ( .a ({new_AGEMA_signal_7491, new_AGEMA_signal_7490, new_AGEMA_signal_7489, SubBytesIns_Inst_Sbox_14_T14}), .b ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, new_AGEMA_signal_8056, SubBytesIns_Inst_Sbox_14_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M4_U1 ( .a ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .c ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_14_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M5_U1 ( .a ({new_AGEMA_signal_7509, new_AGEMA_signal_7508, new_AGEMA_signal_7507, SubBytesIns_Inst_Sbox_14_M4}), .b ({new_AGEMA_signal_7506, new_AGEMA_signal_7505, new_AGEMA_signal_7504, SubBytesIns_Inst_Sbox_14_M1}), .c ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, new_AGEMA_signal_8059, SubBytesIns_Inst_Sbox_14_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M6_U1 ( .a ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774]}), .c ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, SubBytesIns_Inst_Sbox_14_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M7_U1 ( .a ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}), .b ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780]}), .c ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_14_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M8_U1 ( .a ({new_AGEMA_signal_7503, new_AGEMA_signal_7502, new_AGEMA_signal_7501, SubBytesIns_Inst_Sbox_14_T26}), .b ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, new_AGEMA_signal_8062, SubBytesIns_Inst_Sbox_14_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M9_U1 ( .a ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786]}), .c ({new_AGEMA_signal_8067, new_AGEMA_signal_8066, new_AGEMA_signal_8065, SubBytesIns_Inst_Sbox_14_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M10_U1 ( .a ({new_AGEMA_signal_8067, new_AGEMA_signal_8066, new_AGEMA_signal_8065, SubBytesIns_Inst_Sbox_14_M9}), .b ({new_AGEMA_signal_7512, new_AGEMA_signal_7511, new_AGEMA_signal_7510, SubBytesIns_Inst_Sbox_14_M6}), .c ({new_AGEMA_signal_8373, new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_14_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M11_U1 ( .a ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .b ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792]}), .c ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, SubBytesIns_Inst_Sbox_14_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M12_U1 ( .a ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}), .b ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798]}), .c ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_14_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M13_U1 ( .a ({new_AGEMA_signal_7521, new_AGEMA_signal_7520, new_AGEMA_signal_7519, SubBytesIns_Inst_Sbox_14_M12}), .b ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, SubBytesIns_Inst_Sbox_14_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M14_U1 ( .a ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804]}), .c ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, new_AGEMA_signal_8071, SubBytesIns_Inst_Sbox_14_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M15_U1 ( .a ({new_AGEMA_signal_8073, new_AGEMA_signal_8072, new_AGEMA_signal_8071, SubBytesIns_Inst_Sbox_14_M14}), .b ({new_AGEMA_signal_7518, new_AGEMA_signal_7517, new_AGEMA_signal_7516, SubBytesIns_Inst_Sbox_14_M11}), .c ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, new_AGEMA_signal_8374, SubBytesIns_Inst_Sbox_14_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M16_U1 ( .a ({new_AGEMA_signal_8058, new_AGEMA_signal_8057, new_AGEMA_signal_8056, SubBytesIns_Inst_Sbox_14_M3}), .b ({new_AGEMA_signal_8055, new_AGEMA_signal_8054, new_AGEMA_signal_8053, SubBytesIns_Inst_Sbox_14_M2}), .c ({new_AGEMA_signal_8379, new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_14_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M17_U1 ( .a ({new_AGEMA_signal_8061, new_AGEMA_signal_8060, new_AGEMA_signal_8059, SubBytesIns_Inst_Sbox_14_M5}), .b ({new_AGEMA_signal_8049, new_AGEMA_signal_8048, new_AGEMA_signal_8047, SubBytesIns_Inst_Sbox_14_T24}), .c ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, new_AGEMA_signal_8380, SubBytesIns_Inst_Sbox_14_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M18_U1 ( .a ({new_AGEMA_signal_8064, new_AGEMA_signal_8063, new_AGEMA_signal_8062, SubBytesIns_Inst_Sbox_14_M8}), .b ({new_AGEMA_signal_7515, new_AGEMA_signal_7514, new_AGEMA_signal_7513, SubBytesIns_Inst_Sbox_14_M7}), .c ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_14_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M19_U1 ( .a ({new_AGEMA_signal_8373, new_AGEMA_signal_8372, new_AGEMA_signal_8371, SubBytesIns_Inst_Sbox_14_M10}), .b ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, new_AGEMA_signal_8374, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_8619, new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_14_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M20_U1 ( .a ({new_AGEMA_signal_8379, new_AGEMA_signal_8378, new_AGEMA_signal_8377, SubBytesIns_Inst_Sbox_14_M16}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M21_U1 ( .a ({new_AGEMA_signal_8382, new_AGEMA_signal_8381, new_AGEMA_signal_8380, SubBytesIns_Inst_Sbox_14_M17}), .b ({new_AGEMA_signal_8376, new_AGEMA_signal_8375, new_AGEMA_signal_8374, SubBytesIns_Inst_Sbox_14_M15}), .c ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M22_U1 ( .a ({new_AGEMA_signal_8385, new_AGEMA_signal_8384, new_AGEMA_signal_8383, SubBytesIns_Inst_Sbox_14_M18}), .b ({new_AGEMA_signal_8070, new_AGEMA_signal_8069, new_AGEMA_signal_8068, SubBytesIns_Inst_Sbox_14_M13}), .c ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M23_U1 ( .a ({new_AGEMA_signal_8619, new_AGEMA_signal_8618, new_AGEMA_signal_8617, SubBytesIns_Inst_Sbox_14_M19}), .b ({new_AGEMA_signal_8052, new_AGEMA_signal_8051, new_AGEMA_signal_8050, SubBytesIns_Inst_Sbox_14_T25}), .c ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M24_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}), .c ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_14_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M27_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}), .c ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_14_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M1_U1 ( .a ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_15_T13}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810]}), .c ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_15_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M2_U1 ( .a ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_15_T23}), .b ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .c ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, new_AGEMA_signal_8080, SubBytesIns_Inst_Sbox_15_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M3_U1 ( .a ({new_AGEMA_signal_7530, new_AGEMA_signal_7529, new_AGEMA_signal_7528, SubBytesIns_Inst_Sbox_15_T14}), .b ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, new_AGEMA_signal_8083, SubBytesIns_Inst_Sbox_15_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M4_U1 ( .a ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822]}), .c ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, new_AGEMA_signal_7546, SubBytesIns_Inst_Sbox_15_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M5_U1 ( .a ({new_AGEMA_signal_7548, new_AGEMA_signal_7547, new_AGEMA_signal_7546, SubBytesIns_Inst_Sbox_15_M4}), .b ({new_AGEMA_signal_7545, new_AGEMA_signal_7544, new_AGEMA_signal_7543, SubBytesIns_Inst_Sbox_15_M1}), .c ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, new_AGEMA_signal_8086, SubBytesIns_Inst_Sbox_15_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M6_U1 ( .a ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828]}), .c ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_15_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M7_U1 ( .a ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}), .b ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834]}), .c ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, new_AGEMA_signal_7552, SubBytesIns_Inst_Sbox_15_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M8_U1 ( .a ({new_AGEMA_signal_7542, new_AGEMA_signal_7541, new_AGEMA_signal_7540, SubBytesIns_Inst_Sbox_15_T26}), .b ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_8091, new_AGEMA_signal_8090, new_AGEMA_signal_8089, SubBytesIns_Inst_Sbox_15_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M9_U1 ( .a ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840]}), .c ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, new_AGEMA_signal_8092, SubBytesIns_Inst_Sbox_15_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M10_U1 ( .a ({new_AGEMA_signal_8094, new_AGEMA_signal_8093, new_AGEMA_signal_8092, SubBytesIns_Inst_Sbox_15_M9}), .b ({new_AGEMA_signal_7551, new_AGEMA_signal_7550, new_AGEMA_signal_7549, SubBytesIns_Inst_Sbox_15_M6}), .c ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, new_AGEMA_signal_8386, SubBytesIns_Inst_Sbox_15_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M11_U1 ( .a ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .b ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846]}), .c ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_15_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M12_U1 ( .a ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}), .b ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852]}), .c ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, new_AGEMA_signal_7558, SubBytesIns_Inst_Sbox_15_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M13_U1 ( .a ({new_AGEMA_signal_7560, new_AGEMA_signal_7559, new_AGEMA_signal_7558, SubBytesIns_Inst_Sbox_15_M12}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_15_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M14_U1 ( .a ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858]}), .c ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, new_AGEMA_signal_8098, SubBytesIns_Inst_Sbox_15_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M15_U1 ( .a ({new_AGEMA_signal_8100, new_AGEMA_signal_8099, new_AGEMA_signal_8098, SubBytesIns_Inst_Sbox_15_M14}), .b ({new_AGEMA_signal_7557, new_AGEMA_signal_7556, new_AGEMA_signal_7555, SubBytesIns_Inst_Sbox_15_M11}), .c ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_15_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M16_U1 ( .a ({new_AGEMA_signal_8085, new_AGEMA_signal_8084, new_AGEMA_signal_8083, SubBytesIns_Inst_Sbox_15_M3}), .b ({new_AGEMA_signal_8082, new_AGEMA_signal_8081, new_AGEMA_signal_8080, SubBytesIns_Inst_Sbox_15_M2}), .c ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, new_AGEMA_signal_8392, SubBytesIns_Inst_Sbox_15_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M17_U1 ( .a ({new_AGEMA_signal_8088, new_AGEMA_signal_8087, new_AGEMA_signal_8086, SubBytesIns_Inst_Sbox_15_M5}), .b ({new_AGEMA_signal_8076, new_AGEMA_signal_8075, new_AGEMA_signal_8074, SubBytesIns_Inst_Sbox_15_T24}), .c ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_15_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M18_U1 ( .a ({new_AGEMA_signal_8091, new_AGEMA_signal_8090, new_AGEMA_signal_8089, SubBytesIns_Inst_Sbox_15_M8}), .b ({new_AGEMA_signal_7554, new_AGEMA_signal_7553, new_AGEMA_signal_7552, SubBytesIns_Inst_Sbox_15_M7}), .c ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, new_AGEMA_signal_8398, SubBytesIns_Inst_Sbox_15_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M19_U1 ( .a ({new_AGEMA_signal_8388, new_AGEMA_signal_8387, new_AGEMA_signal_8386, SubBytesIns_Inst_Sbox_15_M10}), .b ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_15_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M20_U1 ( .a ({new_AGEMA_signal_8394, new_AGEMA_signal_8393, new_AGEMA_signal_8392, SubBytesIns_Inst_Sbox_15_M16}), .b ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M21_U1 ( .a ({new_AGEMA_signal_8397, new_AGEMA_signal_8396, new_AGEMA_signal_8395, SubBytesIns_Inst_Sbox_15_M17}), .b ({new_AGEMA_signal_8391, new_AGEMA_signal_8390, new_AGEMA_signal_8389, SubBytesIns_Inst_Sbox_15_M15}), .c ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M22_U1 ( .a ({new_AGEMA_signal_8400, new_AGEMA_signal_8399, new_AGEMA_signal_8398, SubBytesIns_Inst_Sbox_15_M18}), .b ({new_AGEMA_signal_8097, new_AGEMA_signal_8096, new_AGEMA_signal_8095, SubBytesIns_Inst_Sbox_15_M13}), .c ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M23_U1 ( .a ({new_AGEMA_signal_8631, new_AGEMA_signal_8630, new_AGEMA_signal_8629, SubBytesIns_Inst_Sbox_15_M19}), .b ({new_AGEMA_signal_8079, new_AGEMA_signal_8078, new_AGEMA_signal_8077, SubBytesIns_Inst_Sbox_15_T25}), .c ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M24_U1 ( .a ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}), .c ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, new_AGEMA_signal_9166, SubBytesIns_Inst_Sbox_15_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M27_U1 ( .a ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}), .c ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_15_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M1_U1 ( .a ({new_AGEMA_signal_6309, new_AGEMA_signal_6308, new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .c ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M2_U1 ( .a ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .b ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870]}), .c ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, new_AGEMA_signal_7567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M3_U1 ( .a ({new_AGEMA_signal_6789, new_AGEMA_signal_6788, new_AGEMA_signal_6787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T14}), .b ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, new_AGEMA_signal_7570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M4_U1 ( .a ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .clk (clk), .r ({Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876]}), .c ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M5_U1 ( .a ({new_AGEMA_signal_6807, new_AGEMA_signal_6806, new_AGEMA_signal_6805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M4}), .b ({new_AGEMA_signal_6804, new_AGEMA_signal_6803, new_AGEMA_signal_6802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M1}), .c ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, new_AGEMA_signal_7573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M6_U1 ( .a ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882]}), .c ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M7_U1 ( .a ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .b ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888]}), .c ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M8_U1 ( .a ({new_AGEMA_signal_6801, new_AGEMA_signal_6800, new_AGEMA_signal_6799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T26}), .b ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, new_AGEMA_signal_7576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M9_U1 ( .a ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894]}), .c ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, new_AGEMA_signal_7579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M10_U1 ( .a ({new_AGEMA_signal_7581, new_AGEMA_signal_7580, new_AGEMA_signal_7579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M9}), .b ({new_AGEMA_signal_6810, new_AGEMA_signal_6809, new_AGEMA_signal_6808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M6}), .c ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, new_AGEMA_signal_8101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M11_U1 ( .a ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900]}), .c ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M12_U1 ( .a ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906]}), .c ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M13_U1 ( .a ({new_AGEMA_signal_6819, new_AGEMA_signal_6818, new_AGEMA_signal_6817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M12}), .b ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M14_U1 ( .a ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .b ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .c ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, new_AGEMA_signal_7585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M15_U1 ( .a ({new_AGEMA_signal_7587, new_AGEMA_signal_7586, new_AGEMA_signal_7585, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M14}), .b ({new_AGEMA_signal_6816, new_AGEMA_signal_6815, new_AGEMA_signal_6814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M11}), .c ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M16_U1 ( .a ({new_AGEMA_signal_7572, new_AGEMA_signal_7571, new_AGEMA_signal_7570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M3}), .b ({new_AGEMA_signal_7569, new_AGEMA_signal_7568, new_AGEMA_signal_7567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M2}), .c ({new_AGEMA_signal_8109, new_AGEMA_signal_8108, new_AGEMA_signal_8107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M17_U1 ( .a ({new_AGEMA_signal_7575, new_AGEMA_signal_7574, new_AGEMA_signal_7573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M5}), .b ({new_AGEMA_signal_7563, new_AGEMA_signal_7562, new_AGEMA_signal_7561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T24}), .c ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, new_AGEMA_signal_8110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M18_U1 ( .a ({new_AGEMA_signal_7578, new_AGEMA_signal_7577, new_AGEMA_signal_7576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M8}), .b ({new_AGEMA_signal_6813, new_AGEMA_signal_6812, new_AGEMA_signal_6811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M7}), .c ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, new_AGEMA_signal_8113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M19_U1 ( .a ({new_AGEMA_signal_8103, new_AGEMA_signal_8102, new_AGEMA_signal_8101, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M10}), .b ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8403, new_AGEMA_signal_8402, new_AGEMA_signal_8401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M20_U1 ( .a ({new_AGEMA_signal_8109, new_AGEMA_signal_8108, new_AGEMA_signal_8107, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M16}), .b ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M21_U1 ( .a ({new_AGEMA_signal_8112, new_AGEMA_signal_8111, new_AGEMA_signal_8110, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M17}), .b ({new_AGEMA_signal_8106, new_AGEMA_signal_8105, new_AGEMA_signal_8104, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M15}), .c ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M22_U1 ( .a ({new_AGEMA_signal_8115, new_AGEMA_signal_8114, new_AGEMA_signal_8113, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M18}), .b ({new_AGEMA_signal_7584, new_AGEMA_signal_7583, new_AGEMA_signal_7582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M13}), .c ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M23_U1 ( .a ({new_AGEMA_signal_8403, new_AGEMA_signal_8402, new_AGEMA_signal_8401, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M19}), .b ({new_AGEMA_signal_7566, new_AGEMA_signal_7565, new_AGEMA_signal_7564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T25}), .c ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M24_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .c ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, new_AGEMA_signal_8881, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M27_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .c ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, new_AGEMA_signal_8647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M1_U1 ( .a ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918]}), .c ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M2_U1 ( .a ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .b ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924]}), .c ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, new_AGEMA_signal_7594, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M3_U1 ( .a ({new_AGEMA_signal_6828, new_AGEMA_signal_6827, new_AGEMA_signal_6826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T14}), .b ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, new_AGEMA_signal_7597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M4_U1 ( .a ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .clk (clk), .r ({Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930]}), .c ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, new_AGEMA_signal_6844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M5_U1 ( .a ({new_AGEMA_signal_6846, new_AGEMA_signal_6845, new_AGEMA_signal_6844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M4}), .b ({new_AGEMA_signal_6843, new_AGEMA_signal_6842, new_AGEMA_signal_6841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M1}), .c ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, new_AGEMA_signal_7600, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M6_U1 ( .a ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936]}), .c ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M7_U1 ( .a ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942]}), .c ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, new_AGEMA_signal_6850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M8_U1 ( .a ({new_AGEMA_signal_6840, new_AGEMA_signal_6839, new_AGEMA_signal_6838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T26}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, new_AGEMA_signal_7603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M9_U1 ( .a ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948]}), .c ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, new_AGEMA_signal_7606, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M10_U1 ( .a ({new_AGEMA_signal_7608, new_AGEMA_signal_7607, new_AGEMA_signal_7606, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M9}), .b ({new_AGEMA_signal_6849, new_AGEMA_signal_6848, new_AGEMA_signal_6847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M6}), .c ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, new_AGEMA_signal_8116, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M11_U1 ( .a ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .b ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954]}), .c ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M12_U1 ( .a ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .b ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .c ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, new_AGEMA_signal_6856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M13_U1 ( .a ({new_AGEMA_signal_6858, new_AGEMA_signal_6857, new_AGEMA_signal_6856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M12}), .b ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, new_AGEMA_signal_7609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M14_U1 ( .a ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966]}), .c ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, new_AGEMA_signal_7612, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M15_U1 ( .a ({new_AGEMA_signal_7614, new_AGEMA_signal_7613, new_AGEMA_signal_7612, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M14}), .b ({new_AGEMA_signal_6855, new_AGEMA_signal_6854, new_AGEMA_signal_6853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M11}), .c ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M16_U1 ( .a ({new_AGEMA_signal_7599, new_AGEMA_signal_7598, new_AGEMA_signal_7597, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M3}), .b ({new_AGEMA_signal_7596, new_AGEMA_signal_7595, new_AGEMA_signal_7594, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M2}), .c ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, new_AGEMA_signal_8122, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M17_U1 ( .a ({new_AGEMA_signal_7602, new_AGEMA_signal_7601, new_AGEMA_signal_7600, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M5}), .b ({new_AGEMA_signal_7590, new_AGEMA_signal_7589, new_AGEMA_signal_7588, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T24}), .c ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, new_AGEMA_signal_8125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M18_U1 ( .a ({new_AGEMA_signal_7605, new_AGEMA_signal_7604, new_AGEMA_signal_7603, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M8}), .b ({new_AGEMA_signal_6852, new_AGEMA_signal_6851, new_AGEMA_signal_6850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M7}), .c ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, new_AGEMA_signal_8128, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M19_U1 ( .a ({new_AGEMA_signal_8118, new_AGEMA_signal_8117, new_AGEMA_signal_8116, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M10}), .b ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, new_AGEMA_signal_8413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M20_U1 ( .a ({new_AGEMA_signal_8124, new_AGEMA_signal_8123, new_AGEMA_signal_8122, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M16}), .b ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, new_AGEMA_signal_7609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M21_U1 ( .a ({new_AGEMA_signal_8127, new_AGEMA_signal_8126, new_AGEMA_signal_8125, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M17}), .b ({new_AGEMA_signal_8121, new_AGEMA_signal_8120, new_AGEMA_signal_8119, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M15}), .c ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M22_U1 ( .a ({new_AGEMA_signal_8130, new_AGEMA_signal_8129, new_AGEMA_signal_8128, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M18}), .b ({new_AGEMA_signal_7611, new_AGEMA_signal_7610, new_AGEMA_signal_7609, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M13}), .c ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M23_U1 ( .a ({new_AGEMA_signal_8415, new_AGEMA_signal_8414, new_AGEMA_signal_8413, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M19}), .b ({new_AGEMA_signal_7593, new_AGEMA_signal_7592, new_AGEMA_signal_7591, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T25}), .c ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M24_U1 ( .a ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .c ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, new_AGEMA_signal_8896, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M27_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .c ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, new_AGEMA_signal_8659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M1_U1 ( .a ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972]}), .c ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M2_U1 ( .a ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .b ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978]}), .c ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, new_AGEMA_signal_7621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M3_U1 ( .a ({new_AGEMA_signal_6867, new_AGEMA_signal_6866, new_AGEMA_signal_6865, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T14}), .b ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, new_AGEMA_signal_7624, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M4_U1 ( .a ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .clk (clk), .r ({Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984]}), .c ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, new_AGEMA_signal_6883, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M5_U1 ( .a ({new_AGEMA_signal_6885, new_AGEMA_signal_6884, new_AGEMA_signal_6883, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M4}), .b ({new_AGEMA_signal_6882, new_AGEMA_signal_6881, new_AGEMA_signal_6880, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M1}), .c ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, new_AGEMA_signal_7627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M6_U1 ( .a ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990]}), .c ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M7_U1 ( .a ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .b ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996]}), .c ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, new_AGEMA_signal_6889, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M8_U1 ( .a ({new_AGEMA_signal_6879, new_AGEMA_signal_6878, new_AGEMA_signal_6877, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T26}), .b ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, new_AGEMA_signal_7630, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M9_U1 ( .a ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002]}), .c ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, new_AGEMA_signal_7633, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M10_U1 ( .a ({new_AGEMA_signal_7635, new_AGEMA_signal_7634, new_AGEMA_signal_7633, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M9}), .b ({new_AGEMA_signal_6888, new_AGEMA_signal_6887, new_AGEMA_signal_6886, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M6}), .c ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, new_AGEMA_signal_8131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M11_U1 ( .a ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .b ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .c ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M12_U1 ( .a ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014]}), .c ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, new_AGEMA_signal_6895, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M13_U1 ( .a ({new_AGEMA_signal_6897, new_AGEMA_signal_6896, new_AGEMA_signal_6895, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M12}), .b ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M14_U1 ( .a ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020]}), .c ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M15_U1 ( .a ({new_AGEMA_signal_7641, new_AGEMA_signal_7640, new_AGEMA_signal_7639, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M14}), .b ({new_AGEMA_signal_6894, new_AGEMA_signal_6893, new_AGEMA_signal_6892, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M11}), .c ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M16_U1 ( .a ({new_AGEMA_signal_7626, new_AGEMA_signal_7625, new_AGEMA_signal_7624, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M3}), .b ({new_AGEMA_signal_7623, new_AGEMA_signal_7622, new_AGEMA_signal_7621, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M2}), .c ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, new_AGEMA_signal_8137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M17_U1 ( .a ({new_AGEMA_signal_7629, new_AGEMA_signal_7628, new_AGEMA_signal_7627, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M5}), .b ({new_AGEMA_signal_7617, new_AGEMA_signal_7616, new_AGEMA_signal_7615, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T24}), .c ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, new_AGEMA_signal_8140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M18_U1 ( .a ({new_AGEMA_signal_7632, new_AGEMA_signal_7631, new_AGEMA_signal_7630, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M8}), .b ({new_AGEMA_signal_6891, new_AGEMA_signal_6890, new_AGEMA_signal_6889, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M7}), .c ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, new_AGEMA_signal_8143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M19_U1 ( .a ({new_AGEMA_signal_8133, new_AGEMA_signal_8132, new_AGEMA_signal_8131, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M10}), .b ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8427, new_AGEMA_signal_8426, new_AGEMA_signal_8425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M20_U1 ( .a ({new_AGEMA_signal_8139, new_AGEMA_signal_8138, new_AGEMA_signal_8137, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M16}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M21_U1 ( .a ({new_AGEMA_signal_8142, new_AGEMA_signal_8141, new_AGEMA_signal_8140, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M17}), .b ({new_AGEMA_signal_8136, new_AGEMA_signal_8135, new_AGEMA_signal_8134, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M15}), .c ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M22_U1 ( .a ({new_AGEMA_signal_8145, new_AGEMA_signal_8144, new_AGEMA_signal_8143, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M18}), .b ({new_AGEMA_signal_7638, new_AGEMA_signal_7637, new_AGEMA_signal_7636, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M13}), .c ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M23_U1 ( .a ({new_AGEMA_signal_8427, new_AGEMA_signal_8426, new_AGEMA_signal_8425, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M19}), .b ({new_AGEMA_signal_7620, new_AGEMA_signal_7619, new_AGEMA_signal_7618, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T25}), .c ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M24_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .c ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, new_AGEMA_signal_8911, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M27_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .c ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, new_AGEMA_signal_8671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M1_U1 ( .a ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026]}), .c ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M2_U1 ( .a ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .b ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032]}), .c ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, new_AGEMA_signal_7648, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M3_U1 ( .a ({new_AGEMA_signal_6906, new_AGEMA_signal_6905, new_AGEMA_signal_6904, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T14}), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M4_U1 ( .a ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .clk (clk), .r ({Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038]}), .c ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, new_AGEMA_signal_6922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M5_U1 ( .a ({new_AGEMA_signal_6924, new_AGEMA_signal_6923, new_AGEMA_signal_6922, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M4}), .b ({new_AGEMA_signal_6921, new_AGEMA_signal_6920, new_AGEMA_signal_6919, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M1}), .c ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, new_AGEMA_signal_7654, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M6_U1 ( .a ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044]}), .c ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M7_U1 ( .a ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050]}), .c ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, new_AGEMA_signal_6928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M8_U1 ( .a ({new_AGEMA_signal_6918, new_AGEMA_signal_6917, new_AGEMA_signal_6916, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T26}), .b ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M9_U1 ( .a ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .b ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056]}), .c ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, new_AGEMA_signal_7660, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M10_U1 ( .a ({new_AGEMA_signal_7662, new_AGEMA_signal_7661, new_AGEMA_signal_7660, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M9}), .b ({new_AGEMA_signal_6927, new_AGEMA_signal_6926, new_AGEMA_signal_6925, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M6}), .c ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, new_AGEMA_signal_8146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M11_U1 ( .a ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .b ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062]}), .c ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M12_U1 ( .a ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .b ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068]}), .c ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, new_AGEMA_signal_6934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M13_U1 ( .a ({new_AGEMA_signal_6936, new_AGEMA_signal_6935, new_AGEMA_signal_6934, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M12}), .b ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M14_U1 ( .a ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074]}), .c ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, new_AGEMA_signal_7666, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M15_U1 ( .a ({new_AGEMA_signal_7668, new_AGEMA_signal_7667, new_AGEMA_signal_7666, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M14}), .b ({new_AGEMA_signal_6933, new_AGEMA_signal_6932, new_AGEMA_signal_6931, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M11}), .c ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M16_U1 ( .a ({new_AGEMA_signal_7653, new_AGEMA_signal_7652, new_AGEMA_signal_7651, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M3}), .b ({new_AGEMA_signal_7650, new_AGEMA_signal_7649, new_AGEMA_signal_7648, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M2}), .c ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, new_AGEMA_signal_8152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M17_U1 ( .a ({new_AGEMA_signal_7656, new_AGEMA_signal_7655, new_AGEMA_signal_7654, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M5}), .b ({new_AGEMA_signal_7644, new_AGEMA_signal_7643, new_AGEMA_signal_7642, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T24}), .c ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, new_AGEMA_signal_8155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M18_U1 ( .a ({new_AGEMA_signal_7659, new_AGEMA_signal_7658, new_AGEMA_signal_7657, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M8}), .b ({new_AGEMA_signal_6930, new_AGEMA_signal_6929, new_AGEMA_signal_6928, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M7}), .c ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, new_AGEMA_signal_8158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M19_U1 ( .a ({new_AGEMA_signal_8148, new_AGEMA_signal_8147, new_AGEMA_signal_8146, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M10}), .b ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, new_AGEMA_signal_8437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M20_U1 ( .a ({new_AGEMA_signal_8154, new_AGEMA_signal_8153, new_AGEMA_signal_8152, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M16}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M21_U1 ( .a ({new_AGEMA_signal_8157, new_AGEMA_signal_8156, new_AGEMA_signal_8155, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M17}), .b ({new_AGEMA_signal_8151, new_AGEMA_signal_8150, new_AGEMA_signal_8149, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M15}), .c ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M22_U1 ( .a ({new_AGEMA_signal_8160, new_AGEMA_signal_8159, new_AGEMA_signal_8158, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M18}), .b ({new_AGEMA_signal_7665, new_AGEMA_signal_7664, new_AGEMA_signal_7663, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M13}), .c ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M23_U1 ( .a ({new_AGEMA_signal_8439, new_AGEMA_signal_8438, new_AGEMA_signal_8437, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M19}), .b ({new_AGEMA_signal_7647, new_AGEMA_signal_7646, new_AGEMA_signal_7645, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T25}), .c ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M24_U1 ( .a ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .c ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, new_AGEMA_signal_8926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M27_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .c ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, new_AGEMA_signal_8683, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080]}), .c ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, new_AGEMA_signal_8944, SubBytesIns_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_8454, new_AGEMA_signal_8453, new_AGEMA_signal_8452, SubBytesIns_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086]}), .c ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, new_AGEMA_signal_8950, SubBytesIns_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8955, new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_8460, new_AGEMA_signal_8459, new_AGEMA_signal_8458, SubBytesIns_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092]}), .c ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, new_AGEMA_signal_8698, SubBytesIns_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_8694, new_AGEMA_signal_8693, new_AGEMA_signal_8692, SubBytesIns_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_9255, new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098]}), .c ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8961, new_AGEMA_signal_8960, new_AGEMA_signal_8959, SubBytesIns_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, new_AGEMA_signal_8962, SubBytesIns_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_8466, new_AGEMA_signal_8465, new_AGEMA_signal_8464, SubBytesIns_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104]}), .c ({new_AGEMA_signal_8967, new_AGEMA_signal_8966, new_AGEMA_signal_8965, SubBytesIns_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, new_AGEMA_signal_8968, SubBytesIns_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_8472, new_AGEMA_signal_8471, new_AGEMA_signal_8470, SubBytesIns_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110]}), .c ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, new_AGEMA_signal_8710, SubBytesIns_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, new_AGEMA_signal_8956, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_8706, new_AGEMA_signal_8705, new_AGEMA_signal_8704, SubBytesIns_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, new_AGEMA_signal_9268, SubBytesIns_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116]}), .c ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, new_AGEMA_signal_8974, SubBytesIns_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, new_AGEMA_signal_8977, SubBytesIns_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_8478, new_AGEMA_signal_8477, new_AGEMA_signal_8476, SubBytesIns_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122]}), .c ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, new_AGEMA_signal_8980, SubBytesIns_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8985, new_AGEMA_signal_8984, new_AGEMA_signal_8983, SubBytesIns_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_8484, new_AGEMA_signal_8483, new_AGEMA_signal_8482, SubBytesIns_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128]}), .c ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, new_AGEMA_signal_8722, SubBytesIns_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, new_AGEMA_signal_8971, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_8718, new_AGEMA_signal_8717, new_AGEMA_signal_8716, SubBytesIns_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_9285, new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134]}), .c ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8991, new_AGEMA_signal_8990, new_AGEMA_signal_8989, SubBytesIns_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, new_AGEMA_signal_8992, SubBytesIns_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_8490, new_AGEMA_signal_8489, new_AGEMA_signal_8488, SubBytesIns_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140]}), .c ({new_AGEMA_signal_8997, new_AGEMA_signal_8996, new_AGEMA_signal_8995, SubBytesIns_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, new_AGEMA_signal_8998, SubBytesIns_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_8496, new_AGEMA_signal_8495, new_AGEMA_signal_8494, SubBytesIns_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146]}), .c ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, new_AGEMA_signal_8734, SubBytesIns_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, new_AGEMA_signal_8986, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_8730, new_AGEMA_signal_8729, new_AGEMA_signal_8728, SubBytesIns_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, new_AGEMA_signal_9298, SubBytesIns_Inst_Sbox_3_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M25_U1 ( .a ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}), .b ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}), .clk (clk), .r ({Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152]}), .c ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M26_U1 ( .a ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, new_AGEMA_signal_9004, SubBytesIns_Inst_Sbox_4_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M28_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9009, new_AGEMA_signal_9008, new_AGEMA_signal_9007, SubBytesIns_Inst_Sbox_4_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M31_U1 ( .a ({new_AGEMA_signal_8502, new_AGEMA_signal_8501, new_AGEMA_signal_8500, SubBytesIns_Inst_Sbox_4_M20}), .b ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}), .clk (clk), .r ({Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158]}), .c ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, new_AGEMA_signal_9010, SubBytesIns_Inst_Sbox_4_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M33_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_4_M27}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9015, new_AGEMA_signal_9014, new_AGEMA_signal_9013, SubBytesIns_Inst_Sbox_4_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M34_U1 ( .a ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_8508, new_AGEMA_signal_8507, new_AGEMA_signal_8506, SubBytesIns_Inst_Sbox_4_M22}), .clk (clk), .r ({Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164]}), .c ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, new_AGEMA_signal_8746, SubBytesIns_Inst_Sbox_4_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M36_U1 ( .a ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, new_AGEMA_signal_9001, SubBytesIns_Inst_Sbox_4_M24}), .b ({new_AGEMA_signal_8742, new_AGEMA_signal_8741, new_AGEMA_signal_8740, SubBytesIns_Inst_Sbox_4_M25}), .c ({new_AGEMA_signal_9315, new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_4_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M25_U1 ( .a ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}), .b ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}), .clk (clk), .r ({Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170]}), .c ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M26_U1 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, new_AGEMA_signal_9019, SubBytesIns_Inst_Sbox_5_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M28_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, new_AGEMA_signal_9022, SubBytesIns_Inst_Sbox_5_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M31_U1 ( .a ({new_AGEMA_signal_8514, new_AGEMA_signal_8513, new_AGEMA_signal_8512, SubBytesIns_Inst_Sbox_5_M20}), .b ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}), .clk (clk), .r ({Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176]}), .c ({new_AGEMA_signal_9027, new_AGEMA_signal_9026, new_AGEMA_signal_9025, SubBytesIns_Inst_Sbox_5_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M33_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_5_M27}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, new_AGEMA_signal_9028, SubBytesIns_Inst_Sbox_5_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M34_U1 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_8520, new_AGEMA_signal_8519, new_AGEMA_signal_8518, SubBytesIns_Inst_Sbox_5_M22}), .clk (clk), .r ({Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182]}), .c ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, new_AGEMA_signal_8758, SubBytesIns_Inst_Sbox_5_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M36_U1 ( .a ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, new_AGEMA_signal_9016, SubBytesIns_Inst_Sbox_5_M24}), .b ({new_AGEMA_signal_8754, new_AGEMA_signal_8753, new_AGEMA_signal_8752, SubBytesIns_Inst_Sbox_5_M25}), .c ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, new_AGEMA_signal_9328, SubBytesIns_Inst_Sbox_5_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M25_U1 ( .a ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}), .b ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}), .clk (clk), .r ({Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188]}), .c ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M26_U1 ( .a ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, new_AGEMA_signal_9034, SubBytesIns_Inst_Sbox_6_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M28_U1 ( .a ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_6_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M31_U1 ( .a ({new_AGEMA_signal_8526, new_AGEMA_signal_8525, new_AGEMA_signal_8524, SubBytesIns_Inst_Sbox_6_M20}), .b ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}), .clk (clk), .r ({Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194]}), .c ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, new_AGEMA_signal_9040, SubBytesIns_Inst_Sbox_6_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M33_U1 ( .a ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_6_M27}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9045, new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_6_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M34_U1 ( .a ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_8532, new_AGEMA_signal_8531, new_AGEMA_signal_8530, SubBytesIns_Inst_Sbox_6_M22}), .clk (clk), .r ({Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200]}), .c ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, new_AGEMA_signal_8770, SubBytesIns_Inst_Sbox_6_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M36_U1 ( .a ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, new_AGEMA_signal_9031, SubBytesIns_Inst_Sbox_6_M24}), .b ({new_AGEMA_signal_8766, new_AGEMA_signal_8765, new_AGEMA_signal_8764, SubBytesIns_Inst_Sbox_6_M25}), .c ({new_AGEMA_signal_9345, new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_6_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M25_U1 ( .a ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}), .b ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}), .clk (clk), .r ({Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206]}), .c ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M26_U1 ( .a ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9051, new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_7_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M28_U1 ( .a ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, new_AGEMA_signal_9052, SubBytesIns_Inst_Sbox_7_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M31_U1 ( .a ({new_AGEMA_signal_8538, new_AGEMA_signal_8537, new_AGEMA_signal_8536, SubBytesIns_Inst_Sbox_7_M20}), .b ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}), .clk (clk), .r ({Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212]}), .c ({new_AGEMA_signal_9057, new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_7_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M33_U1 ( .a ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_7_M27}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, new_AGEMA_signal_9058, SubBytesIns_Inst_Sbox_7_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M34_U1 ( .a ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_8544, new_AGEMA_signal_8543, new_AGEMA_signal_8542, SubBytesIns_Inst_Sbox_7_M22}), .clk (clk), .r ({Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218]}), .c ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, new_AGEMA_signal_8782, SubBytesIns_Inst_Sbox_7_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M36_U1 ( .a ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, new_AGEMA_signal_9046, SubBytesIns_Inst_Sbox_7_M24}), .b ({new_AGEMA_signal_8778, new_AGEMA_signal_8777, new_AGEMA_signal_8776, SubBytesIns_Inst_Sbox_7_M25}), .c ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, new_AGEMA_signal_9358, SubBytesIns_Inst_Sbox_7_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M25_U1 ( .a ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}), .b ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}), .clk (clk), .r ({Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224]}), .c ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M26_U1 ( .a ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, new_AGEMA_signal_9064, SubBytesIns_Inst_Sbox_8_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M28_U1 ( .a ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9069, new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_8_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M31_U1 ( .a ({new_AGEMA_signal_8550, new_AGEMA_signal_8549, new_AGEMA_signal_8548, SubBytesIns_Inst_Sbox_8_M20}), .b ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}), .clk (clk), .r ({Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230]}), .c ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, new_AGEMA_signal_9070, SubBytesIns_Inst_Sbox_8_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M33_U1 ( .a ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_8_M27}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9075, new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_8_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M34_U1 ( .a ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_8556, new_AGEMA_signal_8555, new_AGEMA_signal_8554, SubBytesIns_Inst_Sbox_8_M22}), .clk (clk), .r ({Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236]}), .c ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, new_AGEMA_signal_8794, SubBytesIns_Inst_Sbox_8_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M36_U1 ( .a ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_8_M24}), .b ({new_AGEMA_signal_8790, new_AGEMA_signal_8789, new_AGEMA_signal_8788, SubBytesIns_Inst_Sbox_8_M25}), .c ({new_AGEMA_signal_9375, new_AGEMA_signal_9374, new_AGEMA_signal_9373, SubBytesIns_Inst_Sbox_8_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M25_U1 ( .a ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}), .b ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}), .clk (clk), .r ({Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242]}), .c ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M26_U1 ( .a ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9081, new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_9_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M28_U1 ( .a ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, new_AGEMA_signal_9082, SubBytesIns_Inst_Sbox_9_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M31_U1 ( .a ({new_AGEMA_signal_8562, new_AGEMA_signal_8561, new_AGEMA_signal_8560, SubBytesIns_Inst_Sbox_9_M20}), .b ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}), .clk (clk), .r ({Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248]}), .c ({new_AGEMA_signal_9087, new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_9_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M33_U1 ( .a ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M27}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, new_AGEMA_signal_9088, SubBytesIns_Inst_Sbox_9_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M34_U1 ( .a ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_8568, new_AGEMA_signal_8567, new_AGEMA_signal_8566, SubBytesIns_Inst_Sbox_9_M22}), .clk (clk), .r ({Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254]}), .c ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, new_AGEMA_signal_8806, SubBytesIns_Inst_Sbox_9_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M36_U1 ( .a ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, new_AGEMA_signal_9076, SubBytesIns_Inst_Sbox_9_M24}), .b ({new_AGEMA_signal_8802, new_AGEMA_signal_8801, new_AGEMA_signal_8800, SubBytesIns_Inst_Sbox_9_M25}), .c ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, new_AGEMA_signal_9388, SubBytesIns_Inst_Sbox_9_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M25_U1 ( .a ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}), .b ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}), .clk (clk), .r ({Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260]}), .c ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M26_U1 ( .a ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, new_AGEMA_signal_9094, SubBytesIns_Inst_Sbox_10_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M28_U1 ( .a ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_10_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M31_U1 ( .a ({new_AGEMA_signal_8574, new_AGEMA_signal_8573, new_AGEMA_signal_8572, SubBytesIns_Inst_Sbox_10_M20}), .b ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}), .clk (clk), .r ({Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266]}), .c ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, new_AGEMA_signal_9100, SubBytesIns_Inst_Sbox_10_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M33_U1 ( .a ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M27}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9105, new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_10_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M34_U1 ( .a ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_8580, new_AGEMA_signal_8579, new_AGEMA_signal_8578, SubBytesIns_Inst_Sbox_10_M22}), .clk (clk), .r ({Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272]}), .c ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, new_AGEMA_signal_8818, SubBytesIns_Inst_Sbox_10_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M36_U1 ( .a ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_10_M24}), .b ({new_AGEMA_signal_8814, new_AGEMA_signal_8813, new_AGEMA_signal_8812, SubBytesIns_Inst_Sbox_10_M25}), .c ({new_AGEMA_signal_9405, new_AGEMA_signal_9404, new_AGEMA_signal_9403, SubBytesIns_Inst_Sbox_10_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M25_U1 ( .a ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}), .b ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}), .clk (clk), .r ({Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278]}), .c ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M26_U1 ( .a ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_11_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M28_U1 ( .a ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, new_AGEMA_signal_9112, SubBytesIns_Inst_Sbox_11_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M31_U1 ( .a ({new_AGEMA_signal_8586, new_AGEMA_signal_8585, new_AGEMA_signal_8584, SubBytesIns_Inst_Sbox_11_M20}), .b ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}), .clk (clk), .r ({Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284]}), .c ({new_AGEMA_signal_9117, new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_11_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M33_U1 ( .a ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_11_M27}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, new_AGEMA_signal_9118, SubBytesIns_Inst_Sbox_11_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M34_U1 ( .a ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_8592, new_AGEMA_signal_8591, new_AGEMA_signal_8590, SubBytesIns_Inst_Sbox_11_M22}), .clk (clk), .r ({Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290]}), .c ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, new_AGEMA_signal_8830, SubBytesIns_Inst_Sbox_11_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M36_U1 ( .a ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, new_AGEMA_signal_9106, SubBytesIns_Inst_Sbox_11_M24}), .b ({new_AGEMA_signal_8826, new_AGEMA_signal_8825, new_AGEMA_signal_8824, SubBytesIns_Inst_Sbox_11_M25}), .c ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, new_AGEMA_signal_9418, SubBytesIns_Inst_Sbox_11_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M25_U1 ( .a ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}), .b ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}), .clk (clk), .r ({Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296]}), .c ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M26_U1 ( .a ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, new_AGEMA_signal_9124, SubBytesIns_Inst_Sbox_12_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M28_U1 ( .a ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_12_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M31_U1 ( .a ({new_AGEMA_signal_8598, new_AGEMA_signal_8597, new_AGEMA_signal_8596, SubBytesIns_Inst_Sbox_12_M20}), .b ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}), .clk (clk), .r ({Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302]}), .c ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, new_AGEMA_signal_9130, SubBytesIns_Inst_Sbox_12_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M33_U1 ( .a ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_12_M27}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9135, new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_12_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M34_U1 ( .a ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_8604, new_AGEMA_signal_8603, new_AGEMA_signal_8602, SubBytesIns_Inst_Sbox_12_M22}), .clk (clk), .r ({Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308]}), .c ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, new_AGEMA_signal_8842, SubBytesIns_Inst_Sbox_12_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M36_U1 ( .a ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_12_M24}), .b ({new_AGEMA_signal_8838, new_AGEMA_signal_8837, new_AGEMA_signal_8836, SubBytesIns_Inst_Sbox_12_M25}), .c ({new_AGEMA_signal_9435, new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_12_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M25_U1 ( .a ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}), .b ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}), .clk (clk), .r ({Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314]}), .c ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M26_U1 ( .a ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9141, new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_13_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M28_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, new_AGEMA_signal_9142, SubBytesIns_Inst_Sbox_13_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M31_U1 ( .a ({new_AGEMA_signal_8610, new_AGEMA_signal_8609, new_AGEMA_signal_8608, SubBytesIns_Inst_Sbox_13_M20}), .b ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}), .clk (clk), .r ({Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320]}), .c ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_13_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M33_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_13_M27}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, new_AGEMA_signal_9148, SubBytesIns_Inst_Sbox_13_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M34_U1 ( .a ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_8616, new_AGEMA_signal_8615, new_AGEMA_signal_8614, SubBytesIns_Inst_Sbox_13_M22}), .clk (clk), .r ({Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326]}), .c ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, new_AGEMA_signal_8854, SubBytesIns_Inst_Sbox_13_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M36_U1 ( .a ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, new_AGEMA_signal_9136, SubBytesIns_Inst_Sbox_13_M24}), .b ({new_AGEMA_signal_8850, new_AGEMA_signal_8849, new_AGEMA_signal_8848, SubBytesIns_Inst_Sbox_13_M25}), .c ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, new_AGEMA_signal_9448, SubBytesIns_Inst_Sbox_13_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M25_U1 ( .a ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}), .b ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}), .clk (clk), .r ({Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332]}), .c ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M26_U1 ( .a ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, new_AGEMA_signal_9154, SubBytesIns_Inst_Sbox_14_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M28_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9159, new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_14_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M31_U1 ( .a ({new_AGEMA_signal_8622, new_AGEMA_signal_8621, new_AGEMA_signal_8620, SubBytesIns_Inst_Sbox_14_M20}), .b ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}), .clk (clk), .r ({Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338]}), .c ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, new_AGEMA_signal_9160, SubBytesIns_Inst_Sbox_14_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M33_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_14_M27}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9165, new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_14_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M34_U1 ( .a ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_8628, new_AGEMA_signal_8627, new_AGEMA_signal_8626, SubBytesIns_Inst_Sbox_14_M22}), .clk (clk), .r ({Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344]}), .c ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, new_AGEMA_signal_8866, SubBytesIns_Inst_Sbox_14_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M36_U1 ( .a ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_14_M24}), .b ({new_AGEMA_signal_8862, new_AGEMA_signal_8861, new_AGEMA_signal_8860, SubBytesIns_Inst_Sbox_14_M25}), .c ({new_AGEMA_signal_9465, new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_14_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M25_U1 ( .a ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}), .b ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}), .clk (clk), .r ({Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350]}), .c ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M26_U1 ( .a ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_15_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M28_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, new_AGEMA_signal_9172, SubBytesIns_Inst_Sbox_15_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M31_U1 ( .a ({new_AGEMA_signal_8634, new_AGEMA_signal_8633, new_AGEMA_signal_8632, SubBytesIns_Inst_Sbox_15_M20}), .b ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}), .clk (clk), .r ({Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356]}), .c ({new_AGEMA_signal_9177, new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_15_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M33_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_15_M27}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, new_AGEMA_signal_9178, SubBytesIns_Inst_Sbox_15_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M34_U1 ( .a ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_8640, new_AGEMA_signal_8639, new_AGEMA_signal_8638, SubBytesIns_Inst_Sbox_15_M22}), .clk (clk), .r ({Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362]}), .c ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, new_AGEMA_signal_8878, SubBytesIns_Inst_Sbox_15_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M36_U1 ( .a ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, new_AGEMA_signal_9166, SubBytesIns_Inst_Sbox_15_M24}), .b ({new_AGEMA_signal_8874, new_AGEMA_signal_8873, new_AGEMA_signal_8872, SubBytesIns_Inst_Sbox_15_M25}), .c ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, new_AGEMA_signal_9478, SubBytesIns_Inst_Sbox_15_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M25_U1 ( .a ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .b ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .clk (clk), .r ({Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368]}), .c ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M26_U1 ( .a ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, new_AGEMA_signal_8884, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M28_U1 ( .a ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, new_AGEMA_signal_8887, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M31_U1 ( .a ({new_AGEMA_signal_8406, new_AGEMA_signal_8405, new_AGEMA_signal_8404, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M20}), .b ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .clk (clk), .r ({Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374]}), .c ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, new_AGEMA_signal_8890, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M33_U1 ( .a ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, new_AGEMA_signal_8647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_8895, new_AGEMA_signal_8894, new_AGEMA_signal_8893, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M34_U1 ( .a ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_8412, new_AGEMA_signal_8411, new_AGEMA_signal_8410, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M22}), .clk (clk), .r ({Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380]}), .c ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, new_AGEMA_signal_8650, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M36_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, new_AGEMA_signal_8881, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_8646, new_AGEMA_signal_8645, new_AGEMA_signal_8644, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M25}), .c ({new_AGEMA_signal_9195, new_AGEMA_signal_9194, new_AGEMA_signal_9193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M25_U1 ( .a ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .b ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .clk (clk), .r ({Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386]}), .c ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M26_U1 ( .a ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, new_AGEMA_signal_8899, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M28_U1 ( .a ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, new_AGEMA_signal_8902, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M31_U1 ( .a ({new_AGEMA_signal_8418, new_AGEMA_signal_8417, new_AGEMA_signal_8416, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M20}), .b ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .clk (clk), .r ({Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392]}), .c ({new_AGEMA_signal_8907, new_AGEMA_signal_8906, new_AGEMA_signal_8905, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M33_U1 ( .a ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, new_AGEMA_signal_8659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, new_AGEMA_signal_8908, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M34_U1 ( .a ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_8424, new_AGEMA_signal_8423, new_AGEMA_signal_8422, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M22}), .clk (clk), .r ({Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398]}), .c ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, new_AGEMA_signal_8662, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M36_U1 ( .a ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, new_AGEMA_signal_8896, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_8658, new_AGEMA_signal_8657, new_AGEMA_signal_8656, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M25}), .c ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, new_AGEMA_signal_9208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M25_U1 ( .a ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .b ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .clk (clk), .r ({Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404]}), .c ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M26_U1 ( .a ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, new_AGEMA_signal_8914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M28_U1 ( .a ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8919, new_AGEMA_signal_8918, new_AGEMA_signal_8917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M31_U1 ( .a ({new_AGEMA_signal_8430, new_AGEMA_signal_8429, new_AGEMA_signal_8428, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M20}), .b ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .clk (clk), .r ({Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410]}), .c ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, new_AGEMA_signal_8920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M33_U1 ( .a ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, new_AGEMA_signal_8671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_8925, new_AGEMA_signal_8924, new_AGEMA_signal_8923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M34_U1 ( .a ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_8436, new_AGEMA_signal_8435, new_AGEMA_signal_8434, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M22}), .clk (clk), .r ({Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416]}), .c ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, new_AGEMA_signal_8674, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M36_U1 ( .a ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, new_AGEMA_signal_8911, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_8670, new_AGEMA_signal_8669, new_AGEMA_signal_8668, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M25}), .c ({new_AGEMA_signal_9225, new_AGEMA_signal_9224, new_AGEMA_signal_9223, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M25_U1 ( .a ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .b ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .clk (clk), .r ({Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422]}), .c ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M26_U1 ( .a ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8931, new_AGEMA_signal_8930, new_AGEMA_signal_8929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M28_U1 ( .a ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, new_AGEMA_signal_8932, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M31_U1 ( .a ({new_AGEMA_signal_8442, new_AGEMA_signal_8441, new_AGEMA_signal_8440, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M20}), .b ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .clk (clk), .r ({Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428]}), .c ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, new_AGEMA_signal_8935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M33_U1 ( .a ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, new_AGEMA_signal_8683, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, new_AGEMA_signal_8938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M34_U1 ( .a ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_8448, new_AGEMA_signal_8447, new_AGEMA_signal_8446, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M22}), .clk (clk), .r ({Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434]}), .c ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, new_AGEMA_signal_8686, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M36_U1 ( .a ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, new_AGEMA_signal_8926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_8682, new_AGEMA_signal_8681, new_AGEMA_signal_8680, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M25}), .c ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, new_AGEMA_signal_9238, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_8949, new_AGEMA_signal_8948, new_AGEMA_signal_8947, SubBytesIns_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_0_M27}), .clk (clk), .r ({Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440]}), .c ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_8946, new_AGEMA_signal_8945, new_AGEMA_signal_8944, SubBytesIns_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_0_M24}), .clk (clk), .r ({Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446]}), .c ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, new_AGEMA_signal_9244, SubBytesIns_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_8697, new_AGEMA_signal_8696, new_AGEMA_signal_8695, SubBytesIns_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_8952, new_AGEMA_signal_8951, new_AGEMA_signal_8950, SubBytesIns_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452]}), .c ({new_AGEMA_signal_9249, new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_8943, new_AGEMA_signal_8942, new_AGEMA_signal_8941, SubBytesIns_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_8700, new_AGEMA_signal_8699, new_AGEMA_signal_8698, SubBytesIns_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458]}), .c ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, new_AGEMA_signal_9250, SubBytesIns_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_8457, new_AGEMA_signal_8456, new_AGEMA_signal_8455, SubBytesIns_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_9243, new_AGEMA_signal_9242, new_AGEMA_signal_9241, SubBytesIns_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_9249, new_AGEMA_signal_9248, new_AGEMA_signal_9247, SubBytesIns_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_8955, new_AGEMA_signal_8954, new_AGEMA_signal_8953, SubBytesIns_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_8691, new_AGEMA_signal_8690, new_AGEMA_signal_8689, SubBytesIns_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_9246, new_AGEMA_signal_9245, new_AGEMA_signal_9244, SubBytesIns_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_9252, new_AGEMA_signal_9251, new_AGEMA_signal_9250, SubBytesIns_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_9255, new_AGEMA_signal_9254, new_AGEMA_signal_9253, SubBytesIns_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, new_AGEMA_signal_9874, SubBytesIns_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, new_AGEMA_signal_10585, SubBytesIns_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_8964, new_AGEMA_signal_8963, new_AGEMA_signal_8962, SubBytesIns_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_1_M27}), .clk (clk), .r ({Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464]}), .c ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, new_AGEMA_signal_9256, SubBytesIns_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_8961, new_AGEMA_signal_8960, new_AGEMA_signal_8959, SubBytesIns_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, new_AGEMA_signal_8956, SubBytesIns_Inst_Sbox_1_M24}), .clk (clk), .r ({Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470]}), .c ({new_AGEMA_signal_9261, new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_8709, new_AGEMA_signal_8708, new_AGEMA_signal_8707, SubBytesIns_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_8967, new_AGEMA_signal_8966, new_AGEMA_signal_8965, SubBytesIns_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476]}), .c ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, new_AGEMA_signal_9262, SubBytesIns_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_8958, new_AGEMA_signal_8957, new_AGEMA_signal_8956, SubBytesIns_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_8712, new_AGEMA_signal_8711, new_AGEMA_signal_8710, SubBytesIns_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482]}), .c ({new_AGEMA_signal_9267, new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_8469, new_AGEMA_signal_8468, new_AGEMA_signal_8467, SubBytesIns_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_9258, new_AGEMA_signal_9257, new_AGEMA_signal_9256, SubBytesIns_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_9264, new_AGEMA_signal_9263, new_AGEMA_signal_9262, SubBytesIns_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_8970, new_AGEMA_signal_8969, new_AGEMA_signal_8968, SubBytesIns_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_8703, new_AGEMA_signal_8702, new_AGEMA_signal_8701, SubBytesIns_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_9261, new_AGEMA_signal_9260, new_AGEMA_signal_9259, SubBytesIns_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_9267, new_AGEMA_signal_9266, new_AGEMA_signal_9265, SubBytesIns_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_9270, new_AGEMA_signal_9269, new_AGEMA_signal_9268, SubBytesIns_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910, SubBytesIns_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, new_AGEMA_signal_10621, SubBytesIns_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_8979, new_AGEMA_signal_8978, new_AGEMA_signal_8977, SubBytesIns_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_2_M27}), .clk (clk), .r ({Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488]}), .c ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_8976, new_AGEMA_signal_8975, new_AGEMA_signal_8974, SubBytesIns_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, new_AGEMA_signal_8971, SubBytesIns_Inst_Sbox_2_M24}), .clk (clk), .r ({Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494]}), .c ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, new_AGEMA_signal_9274, SubBytesIns_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_8721, new_AGEMA_signal_8720, new_AGEMA_signal_8719, SubBytesIns_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_8982, new_AGEMA_signal_8981, new_AGEMA_signal_8980, SubBytesIns_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500]}), .c ({new_AGEMA_signal_9279, new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_8973, new_AGEMA_signal_8972, new_AGEMA_signal_8971, SubBytesIns_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_8724, new_AGEMA_signal_8723, new_AGEMA_signal_8722, SubBytesIns_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506]}), .c ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, new_AGEMA_signal_9280, SubBytesIns_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_8481, new_AGEMA_signal_8480, new_AGEMA_signal_8479, SubBytesIns_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_9273, new_AGEMA_signal_9272, new_AGEMA_signal_9271, SubBytesIns_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_9279, new_AGEMA_signal_9278, new_AGEMA_signal_9277, SubBytesIns_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_8985, new_AGEMA_signal_8984, new_AGEMA_signal_8983, SubBytesIns_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_8715, new_AGEMA_signal_8714, new_AGEMA_signal_8713, SubBytesIns_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_9276, new_AGEMA_signal_9275, new_AGEMA_signal_9274, SubBytesIns_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_9282, new_AGEMA_signal_9281, new_AGEMA_signal_9280, SubBytesIns_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_9285, new_AGEMA_signal_9284, new_AGEMA_signal_9283, SubBytesIns_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946, SubBytesIns_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, new_AGEMA_signal_10657, SubBytesIns_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_8994, new_AGEMA_signal_8993, new_AGEMA_signal_8992, SubBytesIns_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_3_M27}), .clk (clk), .r ({Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512]}), .c ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, new_AGEMA_signal_9286, SubBytesIns_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_8991, new_AGEMA_signal_8990, new_AGEMA_signal_8989, SubBytesIns_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, new_AGEMA_signal_8986, SubBytesIns_Inst_Sbox_3_M24}), .clk (clk), .r ({Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518]}), .c ({new_AGEMA_signal_9291, new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_8733, new_AGEMA_signal_8732, new_AGEMA_signal_8731, SubBytesIns_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_8997, new_AGEMA_signal_8996, new_AGEMA_signal_8995, SubBytesIns_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524]}), .c ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, new_AGEMA_signal_9292, SubBytesIns_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_8988, new_AGEMA_signal_8987, new_AGEMA_signal_8986, SubBytesIns_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_8736, new_AGEMA_signal_8735, new_AGEMA_signal_8734, SubBytesIns_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530]}), .c ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_8493, new_AGEMA_signal_8492, new_AGEMA_signal_8491, SubBytesIns_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_9288, new_AGEMA_signal_9287, new_AGEMA_signal_9286, SubBytesIns_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_9294, new_AGEMA_signal_9293, new_AGEMA_signal_9292, SubBytesIns_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_9000, new_AGEMA_signal_8999, new_AGEMA_signal_8998, SubBytesIns_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_8727, new_AGEMA_signal_8726, new_AGEMA_signal_8725, SubBytesIns_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_9291, new_AGEMA_signal_9290, new_AGEMA_signal_9289, SubBytesIns_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_9297, new_AGEMA_signal_9296, new_AGEMA_signal_9295, SubBytesIns_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_9300, new_AGEMA_signal_9299, new_AGEMA_signal_9298, SubBytesIns_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, SubBytesIns_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982, SubBytesIns_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, new_AGEMA_signal_10693, SubBytesIns_Inst_Sbox_3_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M29_U1 ( .a ({new_AGEMA_signal_9009, new_AGEMA_signal_9008, new_AGEMA_signal_9007, SubBytesIns_Inst_Sbox_4_M28}), .b ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_4_M27}), .clk (clk), .r ({Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536]}), .c ({new_AGEMA_signal_9303, new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_4_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M30_U1 ( .a ({new_AGEMA_signal_9006, new_AGEMA_signal_9005, new_AGEMA_signal_9004, SubBytesIns_Inst_Sbox_4_M26}), .b ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, new_AGEMA_signal_9001, SubBytesIns_Inst_Sbox_4_M24}), .clk (clk), .r ({Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542]}), .c ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, new_AGEMA_signal_9304, SubBytesIns_Inst_Sbox_4_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M32_U1 ( .a ({new_AGEMA_signal_8745, new_AGEMA_signal_8744, new_AGEMA_signal_8743, SubBytesIns_Inst_Sbox_4_M27}), .b ({new_AGEMA_signal_9012, new_AGEMA_signal_9011, new_AGEMA_signal_9010, SubBytesIns_Inst_Sbox_4_M31}), .clk (clk), .r ({Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548]}), .c ({new_AGEMA_signal_9309, new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_4_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M35_U1 ( .a ({new_AGEMA_signal_9003, new_AGEMA_signal_9002, new_AGEMA_signal_9001, SubBytesIns_Inst_Sbox_4_M24}), .b ({new_AGEMA_signal_8748, new_AGEMA_signal_8747, new_AGEMA_signal_8746, SubBytesIns_Inst_Sbox_4_M34}), .clk (clk), .r ({Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554]}), .c ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, new_AGEMA_signal_9310, SubBytesIns_Inst_Sbox_4_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M37_U1 ( .a ({new_AGEMA_signal_8505, new_AGEMA_signal_8504, new_AGEMA_signal_8503, SubBytesIns_Inst_Sbox_4_M21}), .b ({new_AGEMA_signal_9303, new_AGEMA_signal_9302, new_AGEMA_signal_9301, SubBytesIns_Inst_Sbox_4_M29}), .c ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M38_U1 ( .a ({new_AGEMA_signal_9309, new_AGEMA_signal_9308, new_AGEMA_signal_9307, SubBytesIns_Inst_Sbox_4_M32}), .b ({new_AGEMA_signal_9015, new_AGEMA_signal_9014, new_AGEMA_signal_9013, SubBytesIns_Inst_Sbox_4_M33}), .c ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M39_U1 ( .a ({new_AGEMA_signal_8739, new_AGEMA_signal_8738, new_AGEMA_signal_8737, SubBytesIns_Inst_Sbox_4_M23}), .b ({new_AGEMA_signal_9306, new_AGEMA_signal_9305, new_AGEMA_signal_9304, SubBytesIns_Inst_Sbox_4_M30}), .c ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M40_U1 ( .a ({new_AGEMA_signal_9312, new_AGEMA_signal_9311, new_AGEMA_signal_9310, SubBytesIns_Inst_Sbox_4_M35}), .b ({new_AGEMA_signal_9315, new_AGEMA_signal_9314, new_AGEMA_signal_9313, SubBytesIns_Inst_Sbox_4_M36}), .c ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M41_U1 ( .a ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M42_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .c ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M43_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .c ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_4_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M44_U1 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .c ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018, SubBytesIns_Inst_Sbox_4_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_M45_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}), .c ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, new_AGEMA_signal_10729, SubBytesIns_Inst_Sbox_4_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M29_U1 ( .a ({new_AGEMA_signal_9024, new_AGEMA_signal_9023, new_AGEMA_signal_9022, SubBytesIns_Inst_Sbox_5_M28}), .b ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_5_M27}), .clk (clk), .r ({Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560]}), .c ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, new_AGEMA_signal_9316, SubBytesIns_Inst_Sbox_5_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M30_U1 ( .a ({new_AGEMA_signal_9021, new_AGEMA_signal_9020, new_AGEMA_signal_9019, SubBytesIns_Inst_Sbox_5_M26}), .b ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, new_AGEMA_signal_9016, SubBytesIns_Inst_Sbox_5_M24}), .clk (clk), .r ({Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566]}), .c ({new_AGEMA_signal_9321, new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_5_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M32_U1 ( .a ({new_AGEMA_signal_8757, new_AGEMA_signal_8756, new_AGEMA_signal_8755, SubBytesIns_Inst_Sbox_5_M27}), .b ({new_AGEMA_signal_9027, new_AGEMA_signal_9026, new_AGEMA_signal_9025, SubBytesIns_Inst_Sbox_5_M31}), .clk (clk), .r ({Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572]}), .c ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, new_AGEMA_signal_9322, SubBytesIns_Inst_Sbox_5_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M35_U1 ( .a ({new_AGEMA_signal_9018, new_AGEMA_signal_9017, new_AGEMA_signal_9016, SubBytesIns_Inst_Sbox_5_M24}), .b ({new_AGEMA_signal_8760, new_AGEMA_signal_8759, new_AGEMA_signal_8758, SubBytesIns_Inst_Sbox_5_M34}), .clk (clk), .r ({Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578]}), .c ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_5_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M37_U1 ( .a ({new_AGEMA_signal_8517, new_AGEMA_signal_8516, new_AGEMA_signal_8515, SubBytesIns_Inst_Sbox_5_M21}), .b ({new_AGEMA_signal_9318, new_AGEMA_signal_9317, new_AGEMA_signal_9316, SubBytesIns_Inst_Sbox_5_M29}), .c ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M38_U1 ( .a ({new_AGEMA_signal_9324, new_AGEMA_signal_9323, new_AGEMA_signal_9322, SubBytesIns_Inst_Sbox_5_M32}), .b ({new_AGEMA_signal_9030, new_AGEMA_signal_9029, new_AGEMA_signal_9028, SubBytesIns_Inst_Sbox_5_M33}), .c ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M39_U1 ( .a ({new_AGEMA_signal_8751, new_AGEMA_signal_8750, new_AGEMA_signal_8749, SubBytesIns_Inst_Sbox_5_M23}), .b ({new_AGEMA_signal_9321, new_AGEMA_signal_9320, new_AGEMA_signal_9319, SubBytesIns_Inst_Sbox_5_M30}), .c ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M40_U1 ( .a ({new_AGEMA_signal_9327, new_AGEMA_signal_9326, new_AGEMA_signal_9325, SubBytesIns_Inst_Sbox_5_M35}), .b ({new_AGEMA_signal_9330, new_AGEMA_signal_9329, new_AGEMA_signal_9328, SubBytesIns_Inst_Sbox_5_M36}), .c ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M41_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M42_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .c ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M43_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .c ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_5_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M44_U1 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .c ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054, SubBytesIns_Inst_Sbox_5_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_M45_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}), .c ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, new_AGEMA_signal_10765, SubBytesIns_Inst_Sbox_5_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M29_U1 ( .a ({new_AGEMA_signal_9039, new_AGEMA_signal_9038, new_AGEMA_signal_9037, SubBytesIns_Inst_Sbox_6_M28}), .b ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_6_M27}), .clk (clk), .r ({Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584]}), .c ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_6_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M30_U1 ( .a ({new_AGEMA_signal_9036, new_AGEMA_signal_9035, new_AGEMA_signal_9034, SubBytesIns_Inst_Sbox_6_M26}), .b ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, new_AGEMA_signal_9031, SubBytesIns_Inst_Sbox_6_M24}), .clk (clk), .r ({Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590]}), .c ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, new_AGEMA_signal_9334, SubBytesIns_Inst_Sbox_6_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M32_U1 ( .a ({new_AGEMA_signal_8769, new_AGEMA_signal_8768, new_AGEMA_signal_8767, SubBytesIns_Inst_Sbox_6_M27}), .b ({new_AGEMA_signal_9042, new_AGEMA_signal_9041, new_AGEMA_signal_9040, SubBytesIns_Inst_Sbox_6_M31}), .clk (clk), .r ({Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596]}), .c ({new_AGEMA_signal_9339, new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_6_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M35_U1 ( .a ({new_AGEMA_signal_9033, new_AGEMA_signal_9032, new_AGEMA_signal_9031, SubBytesIns_Inst_Sbox_6_M24}), .b ({new_AGEMA_signal_8772, new_AGEMA_signal_8771, new_AGEMA_signal_8770, SubBytesIns_Inst_Sbox_6_M34}), .clk (clk), .r ({Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602]}), .c ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, new_AGEMA_signal_9340, SubBytesIns_Inst_Sbox_6_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M37_U1 ( .a ({new_AGEMA_signal_8529, new_AGEMA_signal_8528, new_AGEMA_signal_8527, SubBytesIns_Inst_Sbox_6_M21}), .b ({new_AGEMA_signal_9333, new_AGEMA_signal_9332, new_AGEMA_signal_9331, SubBytesIns_Inst_Sbox_6_M29}), .c ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M38_U1 ( .a ({new_AGEMA_signal_9339, new_AGEMA_signal_9338, new_AGEMA_signal_9337, SubBytesIns_Inst_Sbox_6_M32}), .b ({new_AGEMA_signal_9045, new_AGEMA_signal_9044, new_AGEMA_signal_9043, SubBytesIns_Inst_Sbox_6_M33}), .c ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M39_U1 ( .a ({new_AGEMA_signal_8763, new_AGEMA_signal_8762, new_AGEMA_signal_8761, SubBytesIns_Inst_Sbox_6_M23}), .b ({new_AGEMA_signal_9336, new_AGEMA_signal_9335, new_AGEMA_signal_9334, SubBytesIns_Inst_Sbox_6_M30}), .c ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M40_U1 ( .a ({new_AGEMA_signal_9342, new_AGEMA_signal_9341, new_AGEMA_signal_9340, SubBytesIns_Inst_Sbox_6_M35}), .b ({new_AGEMA_signal_9345, new_AGEMA_signal_9344, new_AGEMA_signal_9343, SubBytesIns_Inst_Sbox_6_M36}), .c ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M41_U1 ( .a ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M42_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .c ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M43_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .c ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_6_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M44_U1 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .c ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, new_AGEMA_signal_10090, SubBytesIns_Inst_Sbox_6_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_M45_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}), .c ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, new_AGEMA_signal_10801, SubBytesIns_Inst_Sbox_6_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M29_U1 ( .a ({new_AGEMA_signal_9054, new_AGEMA_signal_9053, new_AGEMA_signal_9052, SubBytesIns_Inst_Sbox_7_M28}), .b ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_7_M27}), .clk (clk), .r ({Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608]}), .c ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, new_AGEMA_signal_9346, SubBytesIns_Inst_Sbox_7_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M30_U1 ( .a ({new_AGEMA_signal_9051, new_AGEMA_signal_9050, new_AGEMA_signal_9049, SubBytesIns_Inst_Sbox_7_M26}), .b ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, new_AGEMA_signal_9046, SubBytesIns_Inst_Sbox_7_M24}), .clk (clk), .r ({Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614]}), .c ({new_AGEMA_signal_9351, new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_7_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M32_U1 ( .a ({new_AGEMA_signal_8781, new_AGEMA_signal_8780, new_AGEMA_signal_8779, SubBytesIns_Inst_Sbox_7_M27}), .b ({new_AGEMA_signal_9057, new_AGEMA_signal_9056, new_AGEMA_signal_9055, SubBytesIns_Inst_Sbox_7_M31}), .clk (clk), .r ({Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620]}), .c ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, new_AGEMA_signal_9352, SubBytesIns_Inst_Sbox_7_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M35_U1 ( .a ({new_AGEMA_signal_9048, new_AGEMA_signal_9047, new_AGEMA_signal_9046, SubBytesIns_Inst_Sbox_7_M24}), .b ({new_AGEMA_signal_8784, new_AGEMA_signal_8783, new_AGEMA_signal_8782, SubBytesIns_Inst_Sbox_7_M34}), .clk (clk), .r ({Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626]}), .c ({new_AGEMA_signal_9357, new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_7_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M37_U1 ( .a ({new_AGEMA_signal_8541, new_AGEMA_signal_8540, new_AGEMA_signal_8539, SubBytesIns_Inst_Sbox_7_M21}), .b ({new_AGEMA_signal_9348, new_AGEMA_signal_9347, new_AGEMA_signal_9346, SubBytesIns_Inst_Sbox_7_M29}), .c ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M38_U1 ( .a ({new_AGEMA_signal_9354, new_AGEMA_signal_9353, new_AGEMA_signal_9352, SubBytesIns_Inst_Sbox_7_M32}), .b ({new_AGEMA_signal_9060, new_AGEMA_signal_9059, new_AGEMA_signal_9058, SubBytesIns_Inst_Sbox_7_M33}), .c ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M39_U1 ( .a ({new_AGEMA_signal_8775, new_AGEMA_signal_8774, new_AGEMA_signal_8773, SubBytesIns_Inst_Sbox_7_M23}), .b ({new_AGEMA_signal_9351, new_AGEMA_signal_9350, new_AGEMA_signal_9349, SubBytesIns_Inst_Sbox_7_M30}), .c ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M40_U1 ( .a ({new_AGEMA_signal_9357, new_AGEMA_signal_9356, new_AGEMA_signal_9355, SubBytesIns_Inst_Sbox_7_M35}), .b ({new_AGEMA_signal_9360, new_AGEMA_signal_9359, new_AGEMA_signal_9358, SubBytesIns_Inst_Sbox_7_M36}), .c ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M41_U1 ( .a ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M42_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .c ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M43_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .c ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_7_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M44_U1 ( .a ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .c ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, new_AGEMA_signal_10126, SubBytesIns_Inst_Sbox_7_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_M45_U1 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}), .c ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, new_AGEMA_signal_10837, SubBytesIns_Inst_Sbox_7_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M29_U1 ( .a ({new_AGEMA_signal_9069, new_AGEMA_signal_9068, new_AGEMA_signal_9067, SubBytesIns_Inst_Sbox_8_M28}), .b ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_8_M27}), .clk (clk), .r ({Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632]}), .c ({new_AGEMA_signal_9363, new_AGEMA_signal_9362, new_AGEMA_signal_9361, SubBytesIns_Inst_Sbox_8_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M30_U1 ( .a ({new_AGEMA_signal_9066, new_AGEMA_signal_9065, new_AGEMA_signal_9064, SubBytesIns_Inst_Sbox_8_M26}), .b ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_8_M24}), .clk (clk), .r ({Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638]}), .c ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, new_AGEMA_signal_9364, SubBytesIns_Inst_Sbox_8_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M32_U1 ( .a ({new_AGEMA_signal_8793, new_AGEMA_signal_8792, new_AGEMA_signal_8791, SubBytesIns_Inst_Sbox_8_M27}), .b ({new_AGEMA_signal_9072, new_AGEMA_signal_9071, new_AGEMA_signal_9070, SubBytesIns_Inst_Sbox_8_M31}), .clk (clk), .r ({Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644]}), .c ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, new_AGEMA_signal_9367, SubBytesIns_Inst_Sbox_8_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M35_U1 ( .a ({new_AGEMA_signal_9063, new_AGEMA_signal_9062, new_AGEMA_signal_9061, SubBytesIns_Inst_Sbox_8_M24}), .b ({new_AGEMA_signal_8796, new_AGEMA_signal_8795, new_AGEMA_signal_8794, SubBytesIns_Inst_Sbox_8_M34}), .clk (clk), .r ({Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650]}), .c ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, new_AGEMA_signal_9370, SubBytesIns_Inst_Sbox_8_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M37_U1 ( .a ({new_AGEMA_signal_8553, new_AGEMA_signal_8552, new_AGEMA_signal_8551, SubBytesIns_Inst_Sbox_8_M21}), .b ({new_AGEMA_signal_9363, new_AGEMA_signal_9362, new_AGEMA_signal_9361, SubBytesIns_Inst_Sbox_8_M29}), .c ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M38_U1 ( .a ({new_AGEMA_signal_9369, new_AGEMA_signal_9368, new_AGEMA_signal_9367, SubBytesIns_Inst_Sbox_8_M32}), .b ({new_AGEMA_signal_9075, new_AGEMA_signal_9074, new_AGEMA_signal_9073, SubBytesIns_Inst_Sbox_8_M33}), .c ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M39_U1 ( .a ({new_AGEMA_signal_8787, new_AGEMA_signal_8786, new_AGEMA_signal_8785, SubBytesIns_Inst_Sbox_8_M23}), .b ({new_AGEMA_signal_9366, new_AGEMA_signal_9365, new_AGEMA_signal_9364, SubBytesIns_Inst_Sbox_8_M30}), .c ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M40_U1 ( .a ({new_AGEMA_signal_9372, new_AGEMA_signal_9371, new_AGEMA_signal_9370, SubBytesIns_Inst_Sbox_8_M35}), .b ({new_AGEMA_signal_9375, new_AGEMA_signal_9374, new_AGEMA_signal_9373, SubBytesIns_Inst_Sbox_8_M36}), .c ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M41_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M42_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .c ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M43_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .c ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, new_AGEMA_signal_10159, SubBytesIns_Inst_Sbox_8_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M44_U1 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .c ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, new_AGEMA_signal_10162, SubBytesIns_Inst_Sbox_8_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_M45_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}), .c ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, new_AGEMA_signal_10873, SubBytesIns_Inst_Sbox_8_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M29_U1 ( .a ({new_AGEMA_signal_9084, new_AGEMA_signal_9083, new_AGEMA_signal_9082, SubBytesIns_Inst_Sbox_9_M28}), .b ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M27}), .clk (clk), .r ({Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656]}), .c ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, new_AGEMA_signal_9376, SubBytesIns_Inst_Sbox_9_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M30_U1 ( .a ({new_AGEMA_signal_9081, new_AGEMA_signal_9080, new_AGEMA_signal_9079, SubBytesIns_Inst_Sbox_9_M26}), .b ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, new_AGEMA_signal_9076, SubBytesIns_Inst_Sbox_9_M24}), .clk (clk), .r ({Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662]}), .c ({new_AGEMA_signal_9381, new_AGEMA_signal_9380, new_AGEMA_signal_9379, SubBytesIns_Inst_Sbox_9_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M32_U1 ( .a ({new_AGEMA_signal_8805, new_AGEMA_signal_8804, new_AGEMA_signal_8803, SubBytesIns_Inst_Sbox_9_M27}), .b ({new_AGEMA_signal_9087, new_AGEMA_signal_9086, new_AGEMA_signal_9085, SubBytesIns_Inst_Sbox_9_M31}), .clk (clk), .r ({Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668]}), .c ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, new_AGEMA_signal_9382, SubBytesIns_Inst_Sbox_9_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M35_U1 ( .a ({new_AGEMA_signal_9078, new_AGEMA_signal_9077, new_AGEMA_signal_9076, SubBytesIns_Inst_Sbox_9_M24}), .b ({new_AGEMA_signal_8808, new_AGEMA_signal_8807, new_AGEMA_signal_8806, SubBytesIns_Inst_Sbox_9_M34}), .clk (clk), .r ({Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674]}), .c ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, new_AGEMA_signal_9385, SubBytesIns_Inst_Sbox_9_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M37_U1 ( .a ({new_AGEMA_signal_8565, new_AGEMA_signal_8564, new_AGEMA_signal_8563, SubBytesIns_Inst_Sbox_9_M21}), .b ({new_AGEMA_signal_9378, new_AGEMA_signal_9377, new_AGEMA_signal_9376, SubBytesIns_Inst_Sbox_9_M29}), .c ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M38_U1 ( .a ({new_AGEMA_signal_9384, new_AGEMA_signal_9383, new_AGEMA_signal_9382, SubBytesIns_Inst_Sbox_9_M32}), .b ({new_AGEMA_signal_9090, new_AGEMA_signal_9089, new_AGEMA_signal_9088, SubBytesIns_Inst_Sbox_9_M33}), .c ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M39_U1 ( .a ({new_AGEMA_signal_8799, new_AGEMA_signal_8798, new_AGEMA_signal_8797, SubBytesIns_Inst_Sbox_9_M23}), .b ({new_AGEMA_signal_9381, new_AGEMA_signal_9380, new_AGEMA_signal_9379, SubBytesIns_Inst_Sbox_9_M30}), .c ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M40_U1 ( .a ({new_AGEMA_signal_9387, new_AGEMA_signal_9386, new_AGEMA_signal_9385, SubBytesIns_Inst_Sbox_9_M35}), .b ({new_AGEMA_signal_9390, new_AGEMA_signal_9389, new_AGEMA_signal_9388, SubBytesIns_Inst_Sbox_9_M36}), .c ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M41_U1 ( .a ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M42_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .c ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M43_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .c ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, new_AGEMA_signal_10195, SubBytesIns_Inst_Sbox_9_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M44_U1 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .c ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, new_AGEMA_signal_10198, SubBytesIns_Inst_Sbox_9_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_M45_U1 ( .a ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}), .c ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, new_AGEMA_signal_10909, SubBytesIns_Inst_Sbox_9_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M29_U1 ( .a ({new_AGEMA_signal_9099, new_AGEMA_signal_9098, new_AGEMA_signal_9097, SubBytesIns_Inst_Sbox_10_M28}), .b ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M27}), .clk (clk), .r ({Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680]}), .c ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, new_AGEMA_signal_9391, SubBytesIns_Inst_Sbox_10_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M30_U1 ( .a ({new_AGEMA_signal_9096, new_AGEMA_signal_9095, new_AGEMA_signal_9094, SubBytesIns_Inst_Sbox_10_M26}), .b ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_10_M24}), .clk (clk), .r ({Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686]}), .c ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, new_AGEMA_signal_9394, SubBytesIns_Inst_Sbox_10_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M32_U1 ( .a ({new_AGEMA_signal_8817, new_AGEMA_signal_8816, new_AGEMA_signal_8815, SubBytesIns_Inst_Sbox_10_M27}), .b ({new_AGEMA_signal_9102, new_AGEMA_signal_9101, new_AGEMA_signal_9100, SubBytesIns_Inst_Sbox_10_M31}), .clk (clk), .r ({Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692]}), .c ({new_AGEMA_signal_9399, new_AGEMA_signal_9398, new_AGEMA_signal_9397, SubBytesIns_Inst_Sbox_10_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M35_U1 ( .a ({new_AGEMA_signal_9093, new_AGEMA_signal_9092, new_AGEMA_signal_9091, SubBytesIns_Inst_Sbox_10_M24}), .b ({new_AGEMA_signal_8820, new_AGEMA_signal_8819, new_AGEMA_signal_8818, SubBytesIns_Inst_Sbox_10_M34}), .clk (clk), .r ({Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698]}), .c ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, new_AGEMA_signal_9400, SubBytesIns_Inst_Sbox_10_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M37_U1 ( .a ({new_AGEMA_signal_8577, new_AGEMA_signal_8576, new_AGEMA_signal_8575, SubBytesIns_Inst_Sbox_10_M21}), .b ({new_AGEMA_signal_9393, new_AGEMA_signal_9392, new_AGEMA_signal_9391, SubBytesIns_Inst_Sbox_10_M29}), .c ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M38_U1 ( .a ({new_AGEMA_signal_9399, new_AGEMA_signal_9398, new_AGEMA_signal_9397, SubBytesIns_Inst_Sbox_10_M32}), .b ({new_AGEMA_signal_9105, new_AGEMA_signal_9104, new_AGEMA_signal_9103, SubBytesIns_Inst_Sbox_10_M33}), .c ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M39_U1 ( .a ({new_AGEMA_signal_8811, new_AGEMA_signal_8810, new_AGEMA_signal_8809, SubBytesIns_Inst_Sbox_10_M23}), .b ({new_AGEMA_signal_9396, new_AGEMA_signal_9395, new_AGEMA_signal_9394, SubBytesIns_Inst_Sbox_10_M30}), .c ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M40_U1 ( .a ({new_AGEMA_signal_9402, new_AGEMA_signal_9401, new_AGEMA_signal_9400, SubBytesIns_Inst_Sbox_10_M35}), .b ({new_AGEMA_signal_9405, new_AGEMA_signal_9404, new_AGEMA_signal_9403, SubBytesIns_Inst_Sbox_10_M36}), .c ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M41_U1 ( .a ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M42_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .c ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M43_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .c ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, new_AGEMA_signal_10231, SubBytesIns_Inst_Sbox_10_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M44_U1 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .c ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, new_AGEMA_signal_10234, SubBytesIns_Inst_Sbox_10_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_M45_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}), .c ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, new_AGEMA_signal_10945, SubBytesIns_Inst_Sbox_10_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M29_U1 ( .a ({new_AGEMA_signal_9114, new_AGEMA_signal_9113, new_AGEMA_signal_9112, SubBytesIns_Inst_Sbox_11_M28}), .b ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_11_M27}), .clk (clk), .r ({Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704]}), .c ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, new_AGEMA_signal_9406, SubBytesIns_Inst_Sbox_11_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M30_U1 ( .a ({new_AGEMA_signal_9111, new_AGEMA_signal_9110, new_AGEMA_signal_9109, SubBytesIns_Inst_Sbox_11_M26}), .b ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, new_AGEMA_signal_9106, SubBytesIns_Inst_Sbox_11_M24}), .clk (clk), .r ({Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710]}), .c ({new_AGEMA_signal_9411, new_AGEMA_signal_9410, new_AGEMA_signal_9409, SubBytesIns_Inst_Sbox_11_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M32_U1 ( .a ({new_AGEMA_signal_8829, new_AGEMA_signal_8828, new_AGEMA_signal_8827, SubBytesIns_Inst_Sbox_11_M27}), .b ({new_AGEMA_signal_9117, new_AGEMA_signal_9116, new_AGEMA_signal_9115, SubBytesIns_Inst_Sbox_11_M31}), .clk (clk), .r ({Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716]}), .c ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, new_AGEMA_signal_9412, SubBytesIns_Inst_Sbox_11_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M35_U1 ( .a ({new_AGEMA_signal_9108, new_AGEMA_signal_9107, new_AGEMA_signal_9106, SubBytesIns_Inst_Sbox_11_M24}), .b ({new_AGEMA_signal_8832, new_AGEMA_signal_8831, new_AGEMA_signal_8830, SubBytesIns_Inst_Sbox_11_M34}), .clk (clk), .r ({Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722]}), .c ({new_AGEMA_signal_9417, new_AGEMA_signal_9416, new_AGEMA_signal_9415, SubBytesIns_Inst_Sbox_11_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M37_U1 ( .a ({new_AGEMA_signal_8589, new_AGEMA_signal_8588, new_AGEMA_signal_8587, SubBytesIns_Inst_Sbox_11_M21}), .b ({new_AGEMA_signal_9408, new_AGEMA_signal_9407, new_AGEMA_signal_9406, SubBytesIns_Inst_Sbox_11_M29}), .c ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M38_U1 ( .a ({new_AGEMA_signal_9414, new_AGEMA_signal_9413, new_AGEMA_signal_9412, SubBytesIns_Inst_Sbox_11_M32}), .b ({new_AGEMA_signal_9120, new_AGEMA_signal_9119, new_AGEMA_signal_9118, SubBytesIns_Inst_Sbox_11_M33}), .c ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M39_U1 ( .a ({new_AGEMA_signal_8823, new_AGEMA_signal_8822, new_AGEMA_signal_8821, SubBytesIns_Inst_Sbox_11_M23}), .b ({new_AGEMA_signal_9411, new_AGEMA_signal_9410, new_AGEMA_signal_9409, SubBytesIns_Inst_Sbox_11_M30}), .c ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M40_U1 ( .a ({new_AGEMA_signal_9417, new_AGEMA_signal_9416, new_AGEMA_signal_9415, SubBytesIns_Inst_Sbox_11_M35}), .b ({new_AGEMA_signal_9420, new_AGEMA_signal_9419, new_AGEMA_signal_9418, SubBytesIns_Inst_Sbox_11_M36}), .c ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M41_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M42_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .c ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M43_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .c ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, new_AGEMA_signal_10267, SubBytesIns_Inst_Sbox_11_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M44_U1 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .c ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, new_AGEMA_signal_10270, SubBytesIns_Inst_Sbox_11_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_M45_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}), .c ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, new_AGEMA_signal_10981, SubBytesIns_Inst_Sbox_11_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M29_U1 ( .a ({new_AGEMA_signal_9129, new_AGEMA_signal_9128, new_AGEMA_signal_9127, SubBytesIns_Inst_Sbox_12_M28}), .b ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_12_M27}), .clk (clk), .r ({Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728]}), .c ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, new_AGEMA_signal_9421, SubBytesIns_Inst_Sbox_12_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M30_U1 ( .a ({new_AGEMA_signal_9126, new_AGEMA_signal_9125, new_AGEMA_signal_9124, SubBytesIns_Inst_Sbox_12_M26}), .b ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_12_M24}), .clk (clk), .r ({Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734]}), .c ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, new_AGEMA_signal_9424, SubBytesIns_Inst_Sbox_12_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M32_U1 ( .a ({new_AGEMA_signal_8841, new_AGEMA_signal_8840, new_AGEMA_signal_8839, SubBytesIns_Inst_Sbox_12_M27}), .b ({new_AGEMA_signal_9132, new_AGEMA_signal_9131, new_AGEMA_signal_9130, SubBytesIns_Inst_Sbox_12_M31}), .clk (clk), .r ({Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740]}), .c ({new_AGEMA_signal_9429, new_AGEMA_signal_9428, new_AGEMA_signal_9427, SubBytesIns_Inst_Sbox_12_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M35_U1 ( .a ({new_AGEMA_signal_9123, new_AGEMA_signal_9122, new_AGEMA_signal_9121, SubBytesIns_Inst_Sbox_12_M24}), .b ({new_AGEMA_signal_8844, new_AGEMA_signal_8843, new_AGEMA_signal_8842, SubBytesIns_Inst_Sbox_12_M34}), .clk (clk), .r ({Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746]}), .c ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, new_AGEMA_signal_9430, SubBytesIns_Inst_Sbox_12_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M37_U1 ( .a ({new_AGEMA_signal_8601, new_AGEMA_signal_8600, new_AGEMA_signal_8599, SubBytesIns_Inst_Sbox_12_M21}), .b ({new_AGEMA_signal_9423, new_AGEMA_signal_9422, new_AGEMA_signal_9421, SubBytesIns_Inst_Sbox_12_M29}), .c ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M38_U1 ( .a ({new_AGEMA_signal_9429, new_AGEMA_signal_9428, new_AGEMA_signal_9427, SubBytesIns_Inst_Sbox_12_M32}), .b ({new_AGEMA_signal_9135, new_AGEMA_signal_9134, new_AGEMA_signal_9133, SubBytesIns_Inst_Sbox_12_M33}), .c ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M39_U1 ( .a ({new_AGEMA_signal_8835, new_AGEMA_signal_8834, new_AGEMA_signal_8833, SubBytesIns_Inst_Sbox_12_M23}), .b ({new_AGEMA_signal_9426, new_AGEMA_signal_9425, new_AGEMA_signal_9424, SubBytesIns_Inst_Sbox_12_M30}), .c ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M40_U1 ( .a ({new_AGEMA_signal_9432, new_AGEMA_signal_9431, new_AGEMA_signal_9430, SubBytesIns_Inst_Sbox_12_M35}), .b ({new_AGEMA_signal_9435, new_AGEMA_signal_9434, new_AGEMA_signal_9433, SubBytesIns_Inst_Sbox_12_M36}), .c ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M41_U1 ( .a ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M42_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .c ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M43_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .c ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, new_AGEMA_signal_10303, SubBytesIns_Inst_Sbox_12_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M44_U1 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .c ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, new_AGEMA_signal_10306, SubBytesIns_Inst_Sbox_12_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_M45_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}), .c ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, new_AGEMA_signal_11017, SubBytesIns_Inst_Sbox_12_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M29_U1 ( .a ({new_AGEMA_signal_9144, new_AGEMA_signal_9143, new_AGEMA_signal_9142, SubBytesIns_Inst_Sbox_13_M28}), .b ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_13_M27}), .clk (clk), .r ({Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752]}), .c ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, new_AGEMA_signal_9436, SubBytesIns_Inst_Sbox_13_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M30_U1 ( .a ({new_AGEMA_signal_9141, new_AGEMA_signal_9140, new_AGEMA_signal_9139, SubBytesIns_Inst_Sbox_13_M26}), .b ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, new_AGEMA_signal_9136, SubBytesIns_Inst_Sbox_13_M24}), .clk (clk), .r ({Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758]}), .c ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_13_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M32_U1 ( .a ({new_AGEMA_signal_8853, new_AGEMA_signal_8852, new_AGEMA_signal_8851, SubBytesIns_Inst_Sbox_13_M27}), .b ({new_AGEMA_signal_9147, new_AGEMA_signal_9146, new_AGEMA_signal_9145, SubBytesIns_Inst_Sbox_13_M31}), .clk (clk), .r ({Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764]}), .c ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, new_AGEMA_signal_9442, SubBytesIns_Inst_Sbox_13_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M35_U1 ( .a ({new_AGEMA_signal_9138, new_AGEMA_signal_9137, new_AGEMA_signal_9136, SubBytesIns_Inst_Sbox_13_M24}), .b ({new_AGEMA_signal_8856, new_AGEMA_signal_8855, new_AGEMA_signal_8854, SubBytesIns_Inst_Sbox_13_M34}), .clk (clk), .r ({Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770]}), .c ({new_AGEMA_signal_9447, new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_13_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M37_U1 ( .a ({new_AGEMA_signal_8613, new_AGEMA_signal_8612, new_AGEMA_signal_8611, SubBytesIns_Inst_Sbox_13_M21}), .b ({new_AGEMA_signal_9438, new_AGEMA_signal_9437, new_AGEMA_signal_9436, SubBytesIns_Inst_Sbox_13_M29}), .c ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M38_U1 ( .a ({new_AGEMA_signal_9444, new_AGEMA_signal_9443, new_AGEMA_signal_9442, SubBytesIns_Inst_Sbox_13_M32}), .b ({new_AGEMA_signal_9150, new_AGEMA_signal_9149, new_AGEMA_signal_9148, SubBytesIns_Inst_Sbox_13_M33}), .c ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M39_U1 ( .a ({new_AGEMA_signal_8847, new_AGEMA_signal_8846, new_AGEMA_signal_8845, SubBytesIns_Inst_Sbox_13_M23}), .b ({new_AGEMA_signal_9441, new_AGEMA_signal_9440, new_AGEMA_signal_9439, SubBytesIns_Inst_Sbox_13_M30}), .c ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M40_U1 ( .a ({new_AGEMA_signal_9447, new_AGEMA_signal_9446, new_AGEMA_signal_9445, SubBytesIns_Inst_Sbox_13_M35}), .b ({new_AGEMA_signal_9450, new_AGEMA_signal_9449, new_AGEMA_signal_9448, SubBytesIns_Inst_Sbox_13_M36}), .c ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M41_U1 ( .a ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M42_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .c ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M43_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .c ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, new_AGEMA_signal_10339, SubBytesIns_Inst_Sbox_13_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M44_U1 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .c ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, new_AGEMA_signal_10342, SubBytesIns_Inst_Sbox_13_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_M45_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}), .c ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, new_AGEMA_signal_11053, SubBytesIns_Inst_Sbox_13_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M29_U1 ( .a ({new_AGEMA_signal_9159, new_AGEMA_signal_9158, new_AGEMA_signal_9157, SubBytesIns_Inst_Sbox_14_M28}), .b ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_14_M27}), .clk (clk), .r ({Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776]}), .c ({new_AGEMA_signal_9453, new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_14_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M30_U1 ( .a ({new_AGEMA_signal_9156, new_AGEMA_signal_9155, new_AGEMA_signal_9154, SubBytesIns_Inst_Sbox_14_M26}), .b ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_14_M24}), .clk (clk), .r ({Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782]}), .c ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, new_AGEMA_signal_9454, SubBytesIns_Inst_Sbox_14_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M32_U1 ( .a ({new_AGEMA_signal_8865, new_AGEMA_signal_8864, new_AGEMA_signal_8863, SubBytesIns_Inst_Sbox_14_M27}), .b ({new_AGEMA_signal_9162, new_AGEMA_signal_9161, new_AGEMA_signal_9160, SubBytesIns_Inst_Sbox_14_M31}), .clk (clk), .r ({Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788]}), .c ({new_AGEMA_signal_9459, new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_14_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M35_U1 ( .a ({new_AGEMA_signal_9153, new_AGEMA_signal_9152, new_AGEMA_signal_9151, SubBytesIns_Inst_Sbox_14_M24}), .b ({new_AGEMA_signal_8868, new_AGEMA_signal_8867, new_AGEMA_signal_8866, SubBytesIns_Inst_Sbox_14_M34}), .clk (clk), .r ({Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794]}), .c ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, new_AGEMA_signal_9460, SubBytesIns_Inst_Sbox_14_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M37_U1 ( .a ({new_AGEMA_signal_8625, new_AGEMA_signal_8624, new_AGEMA_signal_8623, SubBytesIns_Inst_Sbox_14_M21}), .b ({new_AGEMA_signal_9453, new_AGEMA_signal_9452, new_AGEMA_signal_9451, SubBytesIns_Inst_Sbox_14_M29}), .c ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M38_U1 ( .a ({new_AGEMA_signal_9459, new_AGEMA_signal_9458, new_AGEMA_signal_9457, SubBytesIns_Inst_Sbox_14_M32}), .b ({new_AGEMA_signal_9165, new_AGEMA_signal_9164, new_AGEMA_signal_9163, SubBytesIns_Inst_Sbox_14_M33}), .c ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M39_U1 ( .a ({new_AGEMA_signal_8859, new_AGEMA_signal_8858, new_AGEMA_signal_8857, SubBytesIns_Inst_Sbox_14_M23}), .b ({new_AGEMA_signal_9456, new_AGEMA_signal_9455, new_AGEMA_signal_9454, SubBytesIns_Inst_Sbox_14_M30}), .c ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M40_U1 ( .a ({new_AGEMA_signal_9462, new_AGEMA_signal_9461, new_AGEMA_signal_9460, SubBytesIns_Inst_Sbox_14_M35}), .b ({new_AGEMA_signal_9465, new_AGEMA_signal_9464, new_AGEMA_signal_9463, SubBytesIns_Inst_Sbox_14_M36}), .c ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M41_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M42_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .c ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M43_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .c ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, new_AGEMA_signal_10375, SubBytesIns_Inst_Sbox_14_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M44_U1 ( .a ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .c ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, new_AGEMA_signal_10378, SubBytesIns_Inst_Sbox_14_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_M45_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}), .c ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, new_AGEMA_signal_11089, SubBytesIns_Inst_Sbox_14_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M29_U1 ( .a ({new_AGEMA_signal_9174, new_AGEMA_signal_9173, new_AGEMA_signal_9172, SubBytesIns_Inst_Sbox_15_M28}), .b ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_15_M27}), .clk (clk), .r ({Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800]}), .c ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, new_AGEMA_signal_9466, SubBytesIns_Inst_Sbox_15_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M30_U1 ( .a ({new_AGEMA_signal_9171, new_AGEMA_signal_9170, new_AGEMA_signal_9169, SubBytesIns_Inst_Sbox_15_M26}), .b ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, new_AGEMA_signal_9166, SubBytesIns_Inst_Sbox_15_M24}), .clk (clk), .r ({Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806]}), .c ({new_AGEMA_signal_9471, new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_15_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M32_U1 ( .a ({new_AGEMA_signal_8877, new_AGEMA_signal_8876, new_AGEMA_signal_8875, SubBytesIns_Inst_Sbox_15_M27}), .b ({new_AGEMA_signal_9177, new_AGEMA_signal_9176, new_AGEMA_signal_9175, SubBytesIns_Inst_Sbox_15_M31}), .clk (clk), .r ({Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812]}), .c ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, new_AGEMA_signal_9472, SubBytesIns_Inst_Sbox_15_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M35_U1 ( .a ({new_AGEMA_signal_9168, new_AGEMA_signal_9167, new_AGEMA_signal_9166, SubBytesIns_Inst_Sbox_15_M24}), .b ({new_AGEMA_signal_8880, new_AGEMA_signal_8879, new_AGEMA_signal_8878, SubBytesIns_Inst_Sbox_15_M34}), .clk (clk), .r ({Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818]}), .c ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_15_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M37_U1 ( .a ({new_AGEMA_signal_8637, new_AGEMA_signal_8636, new_AGEMA_signal_8635, SubBytesIns_Inst_Sbox_15_M21}), .b ({new_AGEMA_signal_9468, new_AGEMA_signal_9467, new_AGEMA_signal_9466, SubBytesIns_Inst_Sbox_15_M29}), .c ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M38_U1 ( .a ({new_AGEMA_signal_9474, new_AGEMA_signal_9473, new_AGEMA_signal_9472, SubBytesIns_Inst_Sbox_15_M32}), .b ({new_AGEMA_signal_9180, new_AGEMA_signal_9179, new_AGEMA_signal_9178, SubBytesIns_Inst_Sbox_15_M33}), .c ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M39_U1 ( .a ({new_AGEMA_signal_8871, new_AGEMA_signal_8870, new_AGEMA_signal_8869, SubBytesIns_Inst_Sbox_15_M23}), .b ({new_AGEMA_signal_9471, new_AGEMA_signal_9470, new_AGEMA_signal_9469, SubBytesIns_Inst_Sbox_15_M30}), .c ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M40_U1 ( .a ({new_AGEMA_signal_9477, new_AGEMA_signal_9476, new_AGEMA_signal_9475, SubBytesIns_Inst_Sbox_15_M35}), .b ({new_AGEMA_signal_9480, new_AGEMA_signal_9479, new_AGEMA_signal_9478, SubBytesIns_Inst_Sbox_15_M36}), .c ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M41_U1 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M42_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .c ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M43_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .c ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, new_AGEMA_signal_10411, SubBytesIns_Inst_Sbox_15_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M44_U1 ( .a ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .c ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, new_AGEMA_signal_10414, SubBytesIns_Inst_Sbox_15_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_M45_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}), .c ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, new_AGEMA_signal_11125, SubBytesIns_Inst_Sbox_15_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M29_U1 ( .a ({new_AGEMA_signal_8889, new_AGEMA_signal_8888, new_AGEMA_signal_8887, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M28}), .b ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, new_AGEMA_signal_8647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .clk (clk), .r ({Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824]}), .c ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, new_AGEMA_signal_9181, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M30_U1 ( .a ({new_AGEMA_signal_8886, new_AGEMA_signal_8885, new_AGEMA_signal_8884, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M26}), .b ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, new_AGEMA_signal_8881, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .clk (clk), .r ({Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830]}), .c ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, new_AGEMA_signal_9184, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M32_U1 ( .a ({new_AGEMA_signal_8649, new_AGEMA_signal_8648, new_AGEMA_signal_8647, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M27}), .b ({new_AGEMA_signal_8892, new_AGEMA_signal_8891, new_AGEMA_signal_8890, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M31}), .clk (clk), .r ({Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836]}), .c ({new_AGEMA_signal_9189, new_AGEMA_signal_9188, new_AGEMA_signal_9187, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M35_U1 ( .a ({new_AGEMA_signal_8883, new_AGEMA_signal_8882, new_AGEMA_signal_8881, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M24}), .b ({new_AGEMA_signal_8652, new_AGEMA_signal_8651, new_AGEMA_signal_8650, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M34}), .clk (clk), .r ({Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842]}), .c ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, new_AGEMA_signal_9190, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M37_U1 ( .a ({new_AGEMA_signal_8409, new_AGEMA_signal_8408, new_AGEMA_signal_8407, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M21}), .b ({new_AGEMA_signal_9183, new_AGEMA_signal_9182, new_AGEMA_signal_9181, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M29}), .c ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M38_U1 ( .a ({new_AGEMA_signal_9189, new_AGEMA_signal_9188, new_AGEMA_signal_9187, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M32}), .b ({new_AGEMA_signal_8895, new_AGEMA_signal_8894, new_AGEMA_signal_8893, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M33}), .c ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M39_U1 ( .a ({new_AGEMA_signal_8643, new_AGEMA_signal_8642, new_AGEMA_signal_8641, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M23}), .b ({new_AGEMA_signal_9186, new_AGEMA_signal_9185, new_AGEMA_signal_9184, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M30}), .c ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M40_U1 ( .a ({new_AGEMA_signal_9192, new_AGEMA_signal_9191, new_AGEMA_signal_9190, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M35}), .b ({new_AGEMA_signal_9195, new_AGEMA_signal_9194, new_AGEMA_signal_9193, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M36}), .c ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M41_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M42_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .c ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M43_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .c ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M44_U1 ( .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .c ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, new_AGEMA_signal_9730, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_M45_U1 ( .a ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .c ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, new_AGEMA_signal_10441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M29_U1 ( .a ({new_AGEMA_signal_8904, new_AGEMA_signal_8903, new_AGEMA_signal_8902, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M28}), .b ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, new_AGEMA_signal_8659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .clk (clk), .r ({Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848]}), .c ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, new_AGEMA_signal_9196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M30_U1 ( .a ({new_AGEMA_signal_8901, new_AGEMA_signal_8900, new_AGEMA_signal_8899, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M26}), .b ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, new_AGEMA_signal_8896, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .clk (clk), .r ({Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854]}), .c ({new_AGEMA_signal_9201, new_AGEMA_signal_9200, new_AGEMA_signal_9199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M32_U1 ( .a ({new_AGEMA_signal_8661, new_AGEMA_signal_8660, new_AGEMA_signal_8659, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M27}), .b ({new_AGEMA_signal_8907, new_AGEMA_signal_8906, new_AGEMA_signal_8905, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M31}), .clk (clk), .r ({Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860]}), .c ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, new_AGEMA_signal_9202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M35_U1 ( .a ({new_AGEMA_signal_8898, new_AGEMA_signal_8897, new_AGEMA_signal_8896, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M24}), .b ({new_AGEMA_signal_8664, new_AGEMA_signal_8663, new_AGEMA_signal_8662, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M34}), .clk (clk), .r ({Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866]}), .c ({new_AGEMA_signal_9207, new_AGEMA_signal_9206, new_AGEMA_signal_9205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M37_U1 ( .a ({new_AGEMA_signal_8421, new_AGEMA_signal_8420, new_AGEMA_signal_8419, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M21}), .b ({new_AGEMA_signal_9198, new_AGEMA_signal_9197, new_AGEMA_signal_9196, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M29}), .c ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M38_U1 ( .a ({new_AGEMA_signal_9204, new_AGEMA_signal_9203, new_AGEMA_signal_9202, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M32}), .b ({new_AGEMA_signal_8910, new_AGEMA_signal_8909, new_AGEMA_signal_8908, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M33}), .c ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M39_U1 ( .a ({new_AGEMA_signal_8655, new_AGEMA_signal_8654, new_AGEMA_signal_8653, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M23}), .b ({new_AGEMA_signal_9201, new_AGEMA_signal_9200, new_AGEMA_signal_9199, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M30}), .c ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M40_U1 ( .a ({new_AGEMA_signal_9207, new_AGEMA_signal_9206, new_AGEMA_signal_9205, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M35}), .b ({new_AGEMA_signal_9210, new_AGEMA_signal_9209, new_AGEMA_signal_9208, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M36}), .c ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M41_U1 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M42_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .c ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M43_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .c ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M44_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .c ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, new_AGEMA_signal_9766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_M45_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .c ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M29_U1 ( .a ({new_AGEMA_signal_8919, new_AGEMA_signal_8918, new_AGEMA_signal_8917, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M28}), .b ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, new_AGEMA_signal_8671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .clk (clk), .r ({Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872]}), .c ({new_AGEMA_signal_9213, new_AGEMA_signal_9212, new_AGEMA_signal_9211, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M30_U1 ( .a ({new_AGEMA_signal_8916, new_AGEMA_signal_8915, new_AGEMA_signal_8914, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M26}), .b ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, new_AGEMA_signal_8911, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .clk (clk), .r ({Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878]}), .c ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, new_AGEMA_signal_9214, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M32_U1 ( .a ({new_AGEMA_signal_8673, new_AGEMA_signal_8672, new_AGEMA_signal_8671, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M27}), .b ({new_AGEMA_signal_8922, new_AGEMA_signal_8921, new_AGEMA_signal_8920, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M31}), .clk (clk), .r ({Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884]}), .c ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, new_AGEMA_signal_9217, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M35_U1 ( .a ({new_AGEMA_signal_8913, new_AGEMA_signal_8912, new_AGEMA_signal_8911, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M24}), .b ({new_AGEMA_signal_8676, new_AGEMA_signal_8675, new_AGEMA_signal_8674, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M34}), .clk (clk), .r ({Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890]}), .c ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, new_AGEMA_signal_9220, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M37_U1 ( .a ({new_AGEMA_signal_8433, new_AGEMA_signal_8432, new_AGEMA_signal_8431, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M21}), .b ({new_AGEMA_signal_9213, new_AGEMA_signal_9212, new_AGEMA_signal_9211, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M29}), .c ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M38_U1 ( .a ({new_AGEMA_signal_9219, new_AGEMA_signal_9218, new_AGEMA_signal_9217, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M32}), .b ({new_AGEMA_signal_8925, new_AGEMA_signal_8924, new_AGEMA_signal_8923, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M33}), .c ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M39_U1 ( .a ({new_AGEMA_signal_8667, new_AGEMA_signal_8666, new_AGEMA_signal_8665, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M23}), .b ({new_AGEMA_signal_9216, new_AGEMA_signal_9215, new_AGEMA_signal_9214, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M30}), .c ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M40_U1 ( .a ({new_AGEMA_signal_9222, new_AGEMA_signal_9221, new_AGEMA_signal_9220, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M35}), .b ({new_AGEMA_signal_9225, new_AGEMA_signal_9224, new_AGEMA_signal_9223, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M36}), .c ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M41_U1 ( .a ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M42_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .c ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M43_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .c ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M44_U1 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .c ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, new_AGEMA_signal_9802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_M45_U1 ( .a ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .c ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M29_U1 ( .a ({new_AGEMA_signal_8934, new_AGEMA_signal_8933, new_AGEMA_signal_8932, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M28}), .b ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, new_AGEMA_signal_8683, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .clk (clk), .r ({Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896]}), .c ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, new_AGEMA_signal_9226, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M30_U1 ( .a ({new_AGEMA_signal_8931, new_AGEMA_signal_8930, new_AGEMA_signal_8929, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M26}), .b ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, new_AGEMA_signal_8926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .clk (clk), .r ({Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902]}), .c ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, new_AGEMA_signal_9229, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M32_U1 ( .a ({new_AGEMA_signal_8685, new_AGEMA_signal_8684, new_AGEMA_signal_8683, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M27}), .b ({new_AGEMA_signal_8937, new_AGEMA_signal_8936, new_AGEMA_signal_8935, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M31}), .clk (clk), .r ({Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908]}), .c ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, new_AGEMA_signal_9232, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M35_U1 ( .a ({new_AGEMA_signal_8928, new_AGEMA_signal_8927, new_AGEMA_signal_8926, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M24}), .b ({new_AGEMA_signal_8688, new_AGEMA_signal_8687, new_AGEMA_signal_8686, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M34}), .clk (clk), .r ({Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914]}), .c ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, new_AGEMA_signal_9235, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M37_U1 ( .a ({new_AGEMA_signal_8445, new_AGEMA_signal_8444, new_AGEMA_signal_8443, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M21}), .b ({new_AGEMA_signal_9228, new_AGEMA_signal_9227, new_AGEMA_signal_9226, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M29}), .c ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M38_U1 ( .a ({new_AGEMA_signal_9234, new_AGEMA_signal_9233, new_AGEMA_signal_9232, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M32}), .b ({new_AGEMA_signal_8940, new_AGEMA_signal_8939, new_AGEMA_signal_8938, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M33}), .c ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M39_U1 ( .a ({new_AGEMA_signal_8679, new_AGEMA_signal_8678, new_AGEMA_signal_8677, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M23}), .b ({new_AGEMA_signal_9231, new_AGEMA_signal_9230, new_AGEMA_signal_9229, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M30}), .c ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M40_U1 ( .a ({new_AGEMA_signal_9237, new_AGEMA_signal_9236, new_AGEMA_signal_9235, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M35}), .b ({new_AGEMA_signal_9240, new_AGEMA_signal_9239, new_AGEMA_signal_9238, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M36}), .c ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M41_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M42_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .c ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M43_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .c ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, new_AGEMA_signal_9835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M44_U1 ( .a ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .c ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, new_AGEMA_signal_9838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_M45_U1 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .c ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, new_AGEMA_signal_10549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    mux2_masked #(.security_order(3), .pipeline(0)) U858 ( .s (n321), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .a ({new_AGEMA_signal_15192, new_AGEMA_signal_15191, new_AGEMA_signal_15190, MixColumnsOutput[0]}), .c ({new_AGEMA_signal_15474, new_AGEMA_signal_15473, new_AGEMA_signal_15472, RoundOutput[0]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U859 ( .s (n321), .b ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .a ({new_AGEMA_signal_15717, new_AGEMA_signal_15716, new_AGEMA_signal_15715, MixColumnsOutput[100]}), .c ({new_AGEMA_signal_16053, new_AGEMA_signal_16052, new_AGEMA_signal_16051, RoundOutput[100]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U860 ( .s (n321), .b ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .a ({new_AGEMA_signal_14823, new_AGEMA_signal_14822, new_AGEMA_signal_14821, MixColumnsOutput[101]}), .c ({new_AGEMA_signal_15477, new_AGEMA_signal_15476, new_AGEMA_signal_15475, RoundOutput[101]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U861 ( .s (n321), .b ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .a ({new_AGEMA_signal_14820, new_AGEMA_signal_14819, new_AGEMA_signal_14818, MixColumnsOutput[102]}), .c ({new_AGEMA_signal_15480, new_AGEMA_signal_15479, new_AGEMA_signal_15478, RoundOutput[102]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U862 ( .s (n321), .b ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .a ({new_AGEMA_signal_14817, new_AGEMA_signal_14816, new_AGEMA_signal_14815, MixColumnsOutput[103]}), .c ({new_AGEMA_signal_15483, new_AGEMA_signal_15482, new_AGEMA_signal_15481, RoundOutput[103]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U863 ( .s (n321), .b ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .a ({new_AGEMA_signal_14814, new_AGEMA_signal_14813, new_AGEMA_signal_14812, MixColumnsOutput[104]}), .c ({new_AGEMA_signal_15486, new_AGEMA_signal_15485, new_AGEMA_signal_15484, RoundOutput[104]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U864 ( .s (n321), .b ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .a ({new_AGEMA_signal_15714, new_AGEMA_signal_15713, new_AGEMA_signal_15712, MixColumnsOutput[105]}), .c ({new_AGEMA_signal_16056, new_AGEMA_signal_16055, new_AGEMA_signal_16054, RoundOutput[105]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U865 ( .s (n321), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .a ({new_AGEMA_signal_14901, new_AGEMA_signal_14900, new_AGEMA_signal_14899, MixColumnsOutput[106]}), .c ({new_AGEMA_signal_15489, new_AGEMA_signal_15488, new_AGEMA_signal_15487, RoundOutput[106]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U866 ( .s (n315), .b ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .a ({new_AGEMA_signal_15747, new_AGEMA_signal_15746, new_AGEMA_signal_15745, MixColumnsOutput[107]}), .c ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, new_AGEMA_signal_16057, RoundOutput[107]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U867 ( .s (n316), .b ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .a ({new_AGEMA_signal_15744, new_AGEMA_signal_15743, new_AGEMA_signal_15742, MixColumnsOutput[108]}), .c ({new_AGEMA_signal_16062, new_AGEMA_signal_16061, new_AGEMA_signal_16060, RoundOutput[108]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U868 ( .s (n317), .b ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .a ({new_AGEMA_signal_14892, new_AGEMA_signal_14891, new_AGEMA_signal_14890, MixColumnsOutput[109]}), .c ({new_AGEMA_signal_15492, new_AGEMA_signal_15491, new_AGEMA_signal_15490, RoundOutput[109]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U869 ( .s (n318), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .a ({new_AGEMA_signal_15189, new_AGEMA_signal_15188, new_AGEMA_signal_15187, MixColumnsOutput[10]}), .c ({new_AGEMA_signal_15495, new_AGEMA_signal_15494, new_AGEMA_signal_15493, RoundOutput[10]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U870 ( .s (n319), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .a ({new_AGEMA_signal_14889, new_AGEMA_signal_14888, new_AGEMA_signal_14887, MixColumnsOutput[110]}), .c ({new_AGEMA_signal_15498, new_AGEMA_signal_15497, new_AGEMA_signal_15496, RoundOutput[110]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U871 ( .s (n320), .b ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .a ({new_AGEMA_signal_14886, new_AGEMA_signal_14885, new_AGEMA_signal_14884, MixColumnsOutput[111]}), .c ({new_AGEMA_signal_15501, new_AGEMA_signal_15500, new_AGEMA_signal_15499, RoundOutput[111]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U872 ( .s (n319), .b ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .a ({new_AGEMA_signal_14883, new_AGEMA_signal_14882, new_AGEMA_signal_14881, MixColumnsOutput[112]}), .c ({new_AGEMA_signal_15504, new_AGEMA_signal_15503, new_AGEMA_signal_15502, RoundOutput[112]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U873 ( .s (n318), .b ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .a ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, new_AGEMA_signal_15739, MixColumnsOutput[113]}), .c ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, new_AGEMA_signal_16063, RoundOutput[113]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U874 ( .s (n318), .b ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .a ({new_AGEMA_signal_14877, new_AGEMA_signal_14876, new_AGEMA_signal_14875, MixColumnsOutput[114]}), .c ({new_AGEMA_signal_15507, new_AGEMA_signal_15506, new_AGEMA_signal_15505, RoundOutput[114]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U875 ( .s (n315), .b ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .a ({new_AGEMA_signal_15738, new_AGEMA_signal_15737, new_AGEMA_signal_15736, MixColumnsOutput[115]}), .c ({new_AGEMA_signal_16068, new_AGEMA_signal_16067, new_AGEMA_signal_16066, RoundOutput[115]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U876 ( .s (n316), .b ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .a ({new_AGEMA_signal_15732, new_AGEMA_signal_15731, new_AGEMA_signal_15730, MixColumnsOutput[116]}), .c ({new_AGEMA_signal_16071, new_AGEMA_signal_16070, new_AGEMA_signal_16069, RoundOutput[116]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U877 ( .s (n317), .b ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .a ({new_AGEMA_signal_14865, new_AGEMA_signal_14864, new_AGEMA_signal_14863, MixColumnsOutput[117]}), .c ({new_AGEMA_signal_15510, new_AGEMA_signal_15509, new_AGEMA_signal_15508, RoundOutput[117]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U878 ( .s (n319), .b ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .a ({new_AGEMA_signal_14862, new_AGEMA_signal_14861, new_AGEMA_signal_14860, MixColumnsOutput[118]}), .c ({new_AGEMA_signal_15513, new_AGEMA_signal_15512, new_AGEMA_signal_15511, RoundOutput[118]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U879 ( .s (n320), .b ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .a ({new_AGEMA_signal_14859, new_AGEMA_signal_14858, new_AGEMA_signal_14857, MixColumnsOutput[119]}), .c ({new_AGEMA_signal_15516, new_AGEMA_signal_15515, new_AGEMA_signal_15514, RoundOutput[119]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U880 ( .s (n320), .b ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .a ({new_AGEMA_signal_15855, new_AGEMA_signal_15854, new_AGEMA_signal_15853, MixColumnsOutput[11]}), .c ({new_AGEMA_signal_16074, new_AGEMA_signal_16073, new_AGEMA_signal_16072, RoundOutput[11]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U881 ( .s (n319), .b ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .a ({new_AGEMA_signal_14856, new_AGEMA_signal_14855, new_AGEMA_signal_14854, MixColumnsOutput[120]}), .c ({new_AGEMA_signal_15519, new_AGEMA_signal_15518, new_AGEMA_signal_15517, RoundOutput[120]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U882 ( .s (n318), .b ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .a ({new_AGEMA_signal_15729, new_AGEMA_signal_15728, new_AGEMA_signal_15727, MixColumnsOutput[121]}), .c ({new_AGEMA_signal_16077, new_AGEMA_signal_16076, new_AGEMA_signal_16075, RoundOutput[121]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U883 ( .s (n319), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .a ({new_AGEMA_signal_14850, new_AGEMA_signal_14849, new_AGEMA_signal_14848, MixColumnsOutput[122]}), .c ({new_AGEMA_signal_15522, new_AGEMA_signal_15521, new_AGEMA_signal_15520, RoundOutput[122]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U884 ( .s (n320), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .a ({new_AGEMA_signal_15726, new_AGEMA_signal_15725, new_AGEMA_signal_15724, MixColumnsOutput[123]}), .c ({new_AGEMA_signal_16080, new_AGEMA_signal_16079, new_AGEMA_signal_16078, RoundOutput[123]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U885 ( .s (n316), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .a ({new_AGEMA_signal_15723, new_AGEMA_signal_15722, new_AGEMA_signal_15721, MixColumnsOutput[124]}), .c ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, new_AGEMA_signal_16081, RoundOutput[124]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U886 ( .s (n320), .b ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .a ({new_AGEMA_signal_14841, new_AGEMA_signal_14840, new_AGEMA_signal_14839, MixColumnsOutput[125]}), .c ({new_AGEMA_signal_15525, new_AGEMA_signal_15524, new_AGEMA_signal_15523, RoundOutput[125]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U887 ( .s (n316), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .a ({new_AGEMA_signal_14835, new_AGEMA_signal_14834, new_AGEMA_signal_14833, MixColumnsOutput[126]}), .c ({new_AGEMA_signal_15528, new_AGEMA_signal_15527, new_AGEMA_signal_15526, RoundOutput[126]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U888 ( .s (n317), .b ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .a ({new_AGEMA_signal_14832, new_AGEMA_signal_14831, new_AGEMA_signal_14830, MixColumnsOutput[127]}), .c ({new_AGEMA_signal_15531, new_AGEMA_signal_15530, new_AGEMA_signal_15529, RoundOutput[127]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U889 ( .s (n315), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .a ({new_AGEMA_signal_15852, new_AGEMA_signal_15851, new_AGEMA_signal_15850, MixColumnsOutput[12]}), .c ({new_AGEMA_signal_16086, new_AGEMA_signal_16085, new_AGEMA_signal_16084, RoundOutput[12]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U890 ( .s (n317), .b ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .a ({new_AGEMA_signal_15180, new_AGEMA_signal_15179, new_AGEMA_signal_15178, MixColumnsOutput[13]}), .c ({new_AGEMA_signal_15534, new_AGEMA_signal_15533, new_AGEMA_signal_15532, RoundOutput[13]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U891 ( .s (n316), .b ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .a ({new_AGEMA_signal_15177, new_AGEMA_signal_15176, new_AGEMA_signal_15175, MixColumnsOutput[14]}), .c ({new_AGEMA_signal_15537, new_AGEMA_signal_15536, new_AGEMA_signal_15535, RoundOutput[14]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U892 ( .s (n317), .b ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .a ({new_AGEMA_signal_15174, new_AGEMA_signal_15173, new_AGEMA_signal_15172, MixColumnsOutput[15]}), .c ({new_AGEMA_signal_15540, new_AGEMA_signal_15539, new_AGEMA_signal_15538, RoundOutput[15]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U893 ( .s (n315), .b ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .a ({new_AGEMA_signal_15171, new_AGEMA_signal_15170, new_AGEMA_signal_15169, MixColumnsOutput[16]}), .c ({new_AGEMA_signal_15543, new_AGEMA_signal_15542, new_AGEMA_signal_15541, RoundOutput[16]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U894 ( .s (n318), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .a ({new_AGEMA_signal_15849, new_AGEMA_signal_15848, new_AGEMA_signal_15847, MixColumnsOutput[17]}), .c ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, new_AGEMA_signal_16087, RoundOutput[17]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U895 ( .s (n319), .b ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .a ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, new_AGEMA_signal_15163, MixColumnsOutput[18]}), .c ({new_AGEMA_signal_15546, new_AGEMA_signal_15545, new_AGEMA_signal_15544, RoundOutput[18]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U896 ( .s (n320), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .a ({new_AGEMA_signal_15846, new_AGEMA_signal_15845, new_AGEMA_signal_15844, MixColumnsOutput[19]}), .c ({new_AGEMA_signal_16092, new_AGEMA_signal_16091, new_AGEMA_signal_16090, RoundOutput[19]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U897 ( .s (n318), .b ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .a ({new_AGEMA_signal_15843, new_AGEMA_signal_15842, new_AGEMA_signal_15841, MixColumnsOutput[1]}), .c ({new_AGEMA_signal_16095, new_AGEMA_signal_16094, new_AGEMA_signal_16093, RoundOutput[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U898 ( .s (n319), .b ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .a ({new_AGEMA_signal_15840, new_AGEMA_signal_15839, new_AGEMA_signal_15838, MixColumnsOutput[20]}), .c ({new_AGEMA_signal_16098, new_AGEMA_signal_16097, new_AGEMA_signal_16096, RoundOutput[20]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U899 ( .s (n316), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .a ({new_AGEMA_signal_15153, new_AGEMA_signal_15152, new_AGEMA_signal_15151, MixColumnsOutput[21]}), .c ({new_AGEMA_signal_15549, new_AGEMA_signal_15548, new_AGEMA_signal_15547, RoundOutput[21]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U900 ( .s (n317), .b ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .a ({new_AGEMA_signal_15150, new_AGEMA_signal_15149, new_AGEMA_signal_15148, MixColumnsOutput[22]}), .c ({new_AGEMA_signal_15552, new_AGEMA_signal_15551, new_AGEMA_signal_15550, RoundOutput[22]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U901 ( .s (n315), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .a ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, new_AGEMA_signal_15145, MixColumnsOutput[23]}), .c ({new_AGEMA_signal_15555, new_AGEMA_signal_15554, new_AGEMA_signal_15553, RoundOutput[23]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U902 ( .s (n320), .b ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .a ({new_AGEMA_signal_15144, new_AGEMA_signal_15143, new_AGEMA_signal_15142, MixColumnsOutput[24]}), .c ({new_AGEMA_signal_15558, new_AGEMA_signal_15557, new_AGEMA_signal_15556, RoundOutput[24]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U903 ( .s (n318), .b ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .a ({new_AGEMA_signal_15837, new_AGEMA_signal_15836, new_AGEMA_signal_15835, MixColumnsOutput[25]}), .c ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, new_AGEMA_signal_16099, RoundOutput[25]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U904 ( .s (n316), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .a ({new_AGEMA_signal_15138, new_AGEMA_signal_15137, new_AGEMA_signal_15136, MixColumnsOutput[26]}), .c ({new_AGEMA_signal_15561, new_AGEMA_signal_15560, new_AGEMA_signal_15559, RoundOutput[26]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U905 ( .s (n317), .b ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .a ({new_AGEMA_signal_15834, new_AGEMA_signal_15833, new_AGEMA_signal_15832, MixColumnsOutput[27]}), .c ({new_AGEMA_signal_16104, new_AGEMA_signal_16103, new_AGEMA_signal_16102, RoundOutput[27]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U906 ( .s (n315), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .a ({new_AGEMA_signal_15831, new_AGEMA_signal_15830, new_AGEMA_signal_15829, MixColumnsOutput[28]}), .c ({new_AGEMA_signal_16107, new_AGEMA_signal_16106, new_AGEMA_signal_16105, RoundOutput[28]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U907 ( .s (n319), .b ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .a ({new_AGEMA_signal_15129, new_AGEMA_signal_15128, new_AGEMA_signal_15127, MixColumnsOutput[29]}), .c ({new_AGEMA_signal_15564, new_AGEMA_signal_15563, new_AGEMA_signal_15562, RoundOutput[29]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U908 ( .s (n315), .b ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .a ({new_AGEMA_signal_15126, new_AGEMA_signal_15125, new_AGEMA_signal_15124, MixColumnsOutput[2]}), .c ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, new_AGEMA_signal_15565, RoundOutput[2]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U909 ( .s (n320), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .a ({new_AGEMA_signal_15123, new_AGEMA_signal_15122, new_AGEMA_signal_15121, MixColumnsOutput[30]}), .c ({new_AGEMA_signal_15570, new_AGEMA_signal_15569, new_AGEMA_signal_15568, RoundOutput[30]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U910 ( .s (n318), .b ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .a ({new_AGEMA_signal_15120, new_AGEMA_signal_15119, new_AGEMA_signal_15118, MixColumnsOutput[31]}), .c ({new_AGEMA_signal_15573, new_AGEMA_signal_15572, new_AGEMA_signal_15571, RoundOutput[31]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U911 ( .s (n316), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .a ({new_AGEMA_signal_15096, new_AGEMA_signal_15095, new_AGEMA_signal_15094, MixColumnsOutput[32]}), .c ({new_AGEMA_signal_15576, new_AGEMA_signal_15575, new_AGEMA_signal_15574, RoundOutput[32]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U912 ( .s (n317), .b ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .a ({new_AGEMA_signal_15807, new_AGEMA_signal_15806, new_AGEMA_signal_15805, MixColumnsOutput[33]}), .c ({new_AGEMA_signal_16110, new_AGEMA_signal_16109, new_AGEMA_signal_16108, RoundOutput[33]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U913 ( .s (n315), .b ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .a ({new_AGEMA_signal_15030, new_AGEMA_signal_15029, new_AGEMA_signal_15028, MixColumnsOutput[34]}), .c ({new_AGEMA_signal_15579, new_AGEMA_signal_15578, new_AGEMA_signal_15577, RoundOutput[34]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U914 ( .s (n320), .b ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .a ({new_AGEMA_signal_15792, new_AGEMA_signal_15791, new_AGEMA_signal_15790, MixColumnsOutput[35]}), .c ({new_AGEMA_signal_16113, new_AGEMA_signal_16112, new_AGEMA_signal_16111, RoundOutput[35]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U915 ( .s (n320), .b ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .a ({new_AGEMA_signal_15789, new_AGEMA_signal_15788, new_AGEMA_signal_15787, MixColumnsOutput[36]}), .c ({new_AGEMA_signal_16116, new_AGEMA_signal_16115, new_AGEMA_signal_16114, RoundOutput[36]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U916 ( .s (n320), .b ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .a ({new_AGEMA_signal_15015, new_AGEMA_signal_15014, new_AGEMA_signal_15013, MixColumnsOutput[37]}), .c ({new_AGEMA_signal_15582, new_AGEMA_signal_15581, new_AGEMA_signal_15580, RoundOutput[37]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U917 ( .s (n320), .b ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .a ({new_AGEMA_signal_15012, new_AGEMA_signal_15011, new_AGEMA_signal_15010, MixColumnsOutput[38]}), .c ({new_AGEMA_signal_15585, new_AGEMA_signal_15584, new_AGEMA_signal_15583, RoundOutput[38]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U918 ( .s (n320), .b ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .a ({new_AGEMA_signal_15009, new_AGEMA_signal_15008, new_AGEMA_signal_15007, MixColumnsOutput[39]}), .c ({new_AGEMA_signal_15588, new_AGEMA_signal_15587, new_AGEMA_signal_15586, RoundOutput[39]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U919 ( .s (n320), .b ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .a ({new_AGEMA_signal_15828, new_AGEMA_signal_15827, new_AGEMA_signal_15826, MixColumnsOutput[3]}), .c ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, new_AGEMA_signal_16117, RoundOutput[3]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U920 ( .s (n320), .b ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .a ({new_AGEMA_signal_15006, new_AGEMA_signal_15005, new_AGEMA_signal_15004, MixColumnsOutput[40]}), .c ({new_AGEMA_signal_15591, new_AGEMA_signal_15590, new_AGEMA_signal_15589, RoundOutput[40]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U921 ( .s (n320), .b ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .a ({new_AGEMA_signal_15786, new_AGEMA_signal_15785, new_AGEMA_signal_15784, MixColumnsOutput[41]}), .c ({new_AGEMA_signal_16122, new_AGEMA_signal_16121, new_AGEMA_signal_16120, RoundOutput[41]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U922 ( .s (n320), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .a ({new_AGEMA_signal_15093, new_AGEMA_signal_15092, new_AGEMA_signal_15091, MixColumnsOutput[42]}), .c ({new_AGEMA_signal_15594, new_AGEMA_signal_15593, new_AGEMA_signal_15592, RoundOutput[42]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U923 ( .s (n320), .b ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .a ({new_AGEMA_signal_15819, new_AGEMA_signal_15818, new_AGEMA_signal_15817, MixColumnsOutput[43]}), .c ({new_AGEMA_signal_16125, new_AGEMA_signal_16124, new_AGEMA_signal_16123, RoundOutput[43]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U924 ( .s (n320), .b ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .a ({new_AGEMA_signal_15816, new_AGEMA_signal_15815, new_AGEMA_signal_15814, MixColumnsOutput[44]}), .c ({new_AGEMA_signal_16128, new_AGEMA_signal_16127, new_AGEMA_signal_16126, RoundOutput[44]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U925 ( .s (n320), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .a ({new_AGEMA_signal_15084, new_AGEMA_signal_15083, new_AGEMA_signal_15082, MixColumnsOutput[45]}), .c ({new_AGEMA_signal_15597, new_AGEMA_signal_15596, new_AGEMA_signal_15595, RoundOutput[45]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U926 ( .s (n319), .b ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .a ({new_AGEMA_signal_15081, new_AGEMA_signal_15080, new_AGEMA_signal_15079, MixColumnsOutput[46]}), .c ({new_AGEMA_signal_15600, new_AGEMA_signal_15599, new_AGEMA_signal_15598, RoundOutput[46]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U927 ( .s (n319), .b ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .a ({new_AGEMA_signal_15078, new_AGEMA_signal_15077, new_AGEMA_signal_15076, MixColumnsOutput[47]}), .c ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, new_AGEMA_signal_15601, RoundOutput[47]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U928 ( .s (n319), .b ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .a ({new_AGEMA_signal_15075, new_AGEMA_signal_15074, new_AGEMA_signal_15073, MixColumnsOutput[48]}), .c ({new_AGEMA_signal_15606, new_AGEMA_signal_15605, new_AGEMA_signal_15604, RoundOutput[48]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U929 ( .s (n319), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .a ({new_AGEMA_signal_15813, new_AGEMA_signal_15812, new_AGEMA_signal_15811, MixColumnsOutput[49]}), .c ({new_AGEMA_signal_16131, new_AGEMA_signal_16130, new_AGEMA_signal_16129, RoundOutput[49]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U930 ( .s (n319), .b ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .a ({new_AGEMA_signal_15825, new_AGEMA_signal_15824, new_AGEMA_signal_15823, MixColumnsOutput[4]}), .c ({new_AGEMA_signal_16134, new_AGEMA_signal_16133, new_AGEMA_signal_16132, RoundOutput[4]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U931 ( .s (n319), .b ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .a ({new_AGEMA_signal_15069, new_AGEMA_signal_15068, new_AGEMA_signal_15067, MixColumnsOutput[50]}), .c ({new_AGEMA_signal_15609, new_AGEMA_signal_15608, new_AGEMA_signal_15607, RoundOutput[50]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U932 ( .s (n319), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .a ({new_AGEMA_signal_15810, new_AGEMA_signal_15809, new_AGEMA_signal_15808, MixColumnsOutput[51]}), .c ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, new_AGEMA_signal_16135, RoundOutput[51]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U933 ( .s (n319), .b ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .a ({new_AGEMA_signal_15804, new_AGEMA_signal_15803, new_AGEMA_signal_15802, MixColumnsOutput[52]}), .c ({new_AGEMA_signal_16140, new_AGEMA_signal_16139, new_AGEMA_signal_16138, RoundOutput[52]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U934 ( .s (n319), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .a ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, new_AGEMA_signal_15055, MixColumnsOutput[53]}), .c ({new_AGEMA_signal_15612, new_AGEMA_signal_15611, new_AGEMA_signal_15610, RoundOutput[53]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U935 ( .s (n319), .b ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .a ({new_AGEMA_signal_15054, new_AGEMA_signal_15053, new_AGEMA_signal_15052, MixColumnsOutput[54]}), .c ({new_AGEMA_signal_15615, new_AGEMA_signal_15614, new_AGEMA_signal_15613, RoundOutput[54]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U936 ( .s (n319), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .a ({new_AGEMA_signal_15051, new_AGEMA_signal_15050, new_AGEMA_signal_15049, MixColumnsOutput[55]}), .c ({new_AGEMA_signal_15618, new_AGEMA_signal_15617, new_AGEMA_signal_15616, RoundOutput[55]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U937 ( .s (n319), .b ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .a ({new_AGEMA_signal_15048, new_AGEMA_signal_15047, new_AGEMA_signal_15046, MixColumnsOutput[56]}), .c ({new_AGEMA_signal_15621, new_AGEMA_signal_15620, new_AGEMA_signal_15619, RoundOutput[56]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U938 ( .s (n318), .b ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .a ({new_AGEMA_signal_15801, new_AGEMA_signal_15800, new_AGEMA_signal_15799, MixColumnsOutput[57]}), .c ({new_AGEMA_signal_16143, new_AGEMA_signal_16142, new_AGEMA_signal_16141, RoundOutput[57]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U939 ( .s (n318), .b ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .a ({new_AGEMA_signal_15042, new_AGEMA_signal_15041, new_AGEMA_signal_15040, MixColumnsOutput[58]}), .c ({new_AGEMA_signal_15624, new_AGEMA_signal_15623, new_AGEMA_signal_15622, RoundOutput[58]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U940 ( .s (n318), .b ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .a ({new_AGEMA_signal_15798, new_AGEMA_signal_15797, new_AGEMA_signal_15796, MixColumnsOutput[59]}), .c ({new_AGEMA_signal_16146, new_AGEMA_signal_16145, new_AGEMA_signal_16144, RoundOutput[59]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U941 ( .s (n318), .b ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .a ({new_AGEMA_signal_15111, new_AGEMA_signal_15110, new_AGEMA_signal_15109, MixColumnsOutput[5]}), .c ({new_AGEMA_signal_15627, new_AGEMA_signal_15626, new_AGEMA_signal_15625, RoundOutput[5]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U942 ( .s (n318), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .a ({new_AGEMA_signal_15795, new_AGEMA_signal_15794, new_AGEMA_signal_15793, MixColumnsOutput[60]}), .c ({new_AGEMA_signal_16149, new_AGEMA_signal_16148, new_AGEMA_signal_16147, RoundOutput[60]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U943 ( .s (n318), .b ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .a ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, new_AGEMA_signal_15031, MixColumnsOutput[61]}), .c ({new_AGEMA_signal_15630, new_AGEMA_signal_15629, new_AGEMA_signal_15628, RoundOutput[61]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U944 ( .s (n318), .b ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .a ({new_AGEMA_signal_15027, new_AGEMA_signal_15026, new_AGEMA_signal_15025, MixColumnsOutput[62]}), .c ({new_AGEMA_signal_15633, new_AGEMA_signal_15632, new_AGEMA_signal_15631, RoundOutput[62]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U945 ( .s (n318), .b ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .a ({new_AGEMA_signal_15024, new_AGEMA_signal_15023, new_AGEMA_signal_15022, MixColumnsOutput[63]}), .c ({new_AGEMA_signal_15636, new_AGEMA_signal_15635, new_AGEMA_signal_15634, RoundOutput[63]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U946 ( .s (n318), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .a ({new_AGEMA_signal_15000, new_AGEMA_signal_14999, new_AGEMA_signal_14998, MixColumnsOutput[64]}), .c ({new_AGEMA_signal_15639, new_AGEMA_signal_15638, new_AGEMA_signal_15637, RoundOutput[64]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U947 ( .s (n318), .b ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .a ({new_AGEMA_signal_15771, new_AGEMA_signal_15770, new_AGEMA_signal_15769, MixColumnsOutput[65]}), .c ({new_AGEMA_signal_16152, new_AGEMA_signal_16151, new_AGEMA_signal_16150, RoundOutput[65]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U948 ( .s (n318), .b ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .a ({new_AGEMA_signal_14934, new_AGEMA_signal_14933, new_AGEMA_signal_14932, MixColumnsOutput[66]}), .c ({new_AGEMA_signal_15642, new_AGEMA_signal_15641, new_AGEMA_signal_15640, RoundOutput[66]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U949 ( .s (n318), .b ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .a ({new_AGEMA_signal_15756, new_AGEMA_signal_15755, new_AGEMA_signal_15754, MixColumnsOutput[67]}), .c ({new_AGEMA_signal_16155, new_AGEMA_signal_16154, new_AGEMA_signal_16153, RoundOutput[67]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U950 ( .s (n317), .b ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .a ({new_AGEMA_signal_15753, new_AGEMA_signal_15752, new_AGEMA_signal_15751, MixColumnsOutput[68]}), .c ({new_AGEMA_signal_16158, new_AGEMA_signal_16157, new_AGEMA_signal_16156, RoundOutput[68]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U951 ( .s (n317), .b ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .a ({new_AGEMA_signal_14919, new_AGEMA_signal_14918, new_AGEMA_signal_14917, MixColumnsOutput[69]}), .c ({new_AGEMA_signal_15645, new_AGEMA_signal_15644, new_AGEMA_signal_15643, RoundOutput[69]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U952 ( .s (n317), .b ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .a ({new_AGEMA_signal_15108, new_AGEMA_signal_15107, new_AGEMA_signal_15106, MixColumnsOutput[6]}), .c ({new_AGEMA_signal_15648, new_AGEMA_signal_15647, new_AGEMA_signal_15646, RoundOutput[6]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U953 ( .s (n317), .b ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .a ({new_AGEMA_signal_14916, new_AGEMA_signal_14915, new_AGEMA_signal_14914, MixColumnsOutput[70]}), .c ({new_AGEMA_signal_15651, new_AGEMA_signal_15650, new_AGEMA_signal_15649, RoundOutput[70]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U954 ( .s (n317), .b ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .a ({new_AGEMA_signal_14913, new_AGEMA_signal_14912, new_AGEMA_signal_14911, MixColumnsOutput[71]}), .c ({new_AGEMA_signal_15654, new_AGEMA_signal_15653, new_AGEMA_signal_15652, RoundOutput[71]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U955 ( .s (n317), .b ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .a ({new_AGEMA_signal_14910, new_AGEMA_signal_14909, new_AGEMA_signal_14908, MixColumnsOutput[72]}), .c ({new_AGEMA_signal_15657, new_AGEMA_signal_15656, new_AGEMA_signal_15655, RoundOutput[72]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U956 ( .s (n317), .b ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .a ({new_AGEMA_signal_15750, new_AGEMA_signal_15749, new_AGEMA_signal_15748, MixColumnsOutput[73]}), .c ({new_AGEMA_signal_16161, new_AGEMA_signal_16160, new_AGEMA_signal_16159, RoundOutput[73]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U957 ( .s (n317), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .a ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, new_AGEMA_signal_14995, MixColumnsOutput[74]}), .c ({new_AGEMA_signal_15660, new_AGEMA_signal_15659, new_AGEMA_signal_15658, RoundOutput[74]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U958 ( .s (n317), .b ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .a ({new_AGEMA_signal_15783, new_AGEMA_signal_15782, new_AGEMA_signal_15781, MixColumnsOutput[75]}), .c ({new_AGEMA_signal_16164, new_AGEMA_signal_16163, new_AGEMA_signal_16162, RoundOutput[75]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U959 ( .s (n317), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .a ({new_AGEMA_signal_15780, new_AGEMA_signal_15779, new_AGEMA_signal_15778, MixColumnsOutput[76]}), .c ({new_AGEMA_signal_16167, new_AGEMA_signal_16166, new_AGEMA_signal_16165, RoundOutput[76]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U960 ( .s (n317), .b ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .a ({new_AGEMA_signal_14988, new_AGEMA_signal_14987, new_AGEMA_signal_14986, MixColumnsOutput[77]}), .c ({new_AGEMA_signal_15663, new_AGEMA_signal_15662, new_AGEMA_signal_15661, RoundOutput[77]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U961 ( .s (n317), .b ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .a ({new_AGEMA_signal_14985, new_AGEMA_signal_14984, new_AGEMA_signal_14983, MixColumnsOutput[78]}), .c ({new_AGEMA_signal_15666, new_AGEMA_signal_15665, new_AGEMA_signal_15664, RoundOutput[78]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U962 ( .s (n316), .b ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .a ({new_AGEMA_signal_14982, new_AGEMA_signal_14981, new_AGEMA_signal_14980, MixColumnsOutput[79]}), .c ({new_AGEMA_signal_15669, new_AGEMA_signal_15668, new_AGEMA_signal_15667, RoundOutput[79]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U963 ( .s (n316), .b ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .a ({new_AGEMA_signal_15105, new_AGEMA_signal_15104, new_AGEMA_signal_15103, MixColumnsOutput[7]}), .c ({new_AGEMA_signal_15672, new_AGEMA_signal_15671, new_AGEMA_signal_15670, RoundOutput[7]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U964 ( .s (n316), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .a ({new_AGEMA_signal_14979, new_AGEMA_signal_14978, new_AGEMA_signal_14977, MixColumnsOutput[80]}), .c ({new_AGEMA_signal_15675, new_AGEMA_signal_15674, new_AGEMA_signal_15673, RoundOutput[80]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U965 ( .s (n316), .b ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .a ({new_AGEMA_signal_15777, new_AGEMA_signal_15776, new_AGEMA_signal_15775, MixColumnsOutput[81]}), .c ({new_AGEMA_signal_16170, new_AGEMA_signal_16169, new_AGEMA_signal_16168, RoundOutput[81]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U966 ( .s (n316), .b ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .a ({new_AGEMA_signal_14973, new_AGEMA_signal_14972, new_AGEMA_signal_14971, MixColumnsOutput[82]}), .c ({new_AGEMA_signal_15678, new_AGEMA_signal_15677, new_AGEMA_signal_15676, RoundOutput[82]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U967 ( .s (n316), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .a ({new_AGEMA_signal_15774, new_AGEMA_signal_15773, new_AGEMA_signal_15772, MixColumnsOutput[83]}), .c ({new_AGEMA_signal_16173, new_AGEMA_signal_16172, new_AGEMA_signal_16171, RoundOutput[83]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U968 ( .s (n316), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .a ({new_AGEMA_signal_15768, new_AGEMA_signal_15767, new_AGEMA_signal_15766, MixColumnsOutput[84]}), .c ({new_AGEMA_signal_16176, new_AGEMA_signal_16175, new_AGEMA_signal_16174, RoundOutput[84]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U969 ( .s (n316), .b ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .a ({new_AGEMA_signal_14961, new_AGEMA_signal_14960, new_AGEMA_signal_14959, MixColumnsOutput[85]}), .c ({new_AGEMA_signal_15681, new_AGEMA_signal_15680, new_AGEMA_signal_15679, RoundOutput[85]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U970 ( .s (n316), .b ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .a ({new_AGEMA_signal_14958, new_AGEMA_signal_14957, new_AGEMA_signal_14956, MixColumnsOutput[86]}), .c ({new_AGEMA_signal_15684, new_AGEMA_signal_15683, new_AGEMA_signal_15682, RoundOutput[86]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U971 ( .s (n316), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .a ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, new_AGEMA_signal_14953, MixColumnsOutput[87]}), .c ({new_AGEMA_signal_15687, new_AGEMA_signal_15686, new_AGEMA_signal_15685, RoundOutput[87]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U972 ( .s (n316), .b ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .a ({new_AGEMA_signal_14952, new_AGEMA_signal_14951, new_AGEMA_signal_14950, MixColumnsOutput[88]}), .c ({new_AGEMA_signal_15690, new_AGEMA_signal_15689, new_AGEMA_signal_15688, RoundOutput[88]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U973 ( .s (n316), .b ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .a ({new_AGEMA_signal_15765, new_AGEMA_signal_15764, new_AGEMA_signal_15763, MixColumnsOutput[89]}), .c ({new_AGEMA_signal_16179, new_AGEMA_signal_16178, new_AGEMA_signal_16177, RoundOutput[89]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U974 ( .s (n315), .b ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .a ({new_AGEMA_signal_15102, new_AGEMA_signal_15101, new_AGEMA_signal_15100, MixColumnsOutput[8]}), .c ({new_AGEMA_signal_15693, new_AGEMA_signal_15692, new_AGEMA_signal_15691, RoundOutput[8]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U975 ( .s (n315), .b ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .a ({new_AGEMA_signal_14946, new_AGEMA_signal_14945, new_AGEMA_signal_14944, MixColumnsOutput[90]}), .c ({new_AGEMA_signal_15696, new_AGEMA_signal_15695, new_AGEMA_signal_15694, RoundOutput[90]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U976 ( .s (n315), .b ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .a ({new_AGEMA_signal_15762, new_AGEMA_signal_15761, new_AGEMA_signal_15760, MixColumnsOutput[91]}), .c ({new_AGEMA_signal_16182, new_AGEMA_signal_16181, new_AGEMA_signal_16180, RoundOutput[91]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U977 ( .s (n315), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .a ({new_AGEMA_signal_15759, new_AGEMA_signal_15758, new_AGEMA_signal_15757, MixColumnsOutput[92]}), .c ({new_AGEMA_signal_16185, new_AGEMA_signal_16184, new_AGEMA_signal_16183, RoundOutput[92]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U978 ( .s (n315), .b ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .a ({new_AGEMA_signal_14937, new_AGEMA_signal_14936, new_AGEMA_signal_14935, MixColumnsOutput[93]}), .c ({new_AGEMA_signal_15699, new_AGEMA_signal_15698, new_AGEMA_signal_15697, RoundOutput[93]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U979 ( .s (n315), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .a ({new_AGEMA_signal_14931, new_AGEMA_signal_14930, new_AGEMA_signal_14929, MixColumnsOutput[94]}), .c ({new_AGEMA_signal_15702, new_AGEMA_signal_15701, new_AGEMA_signal_15700, RoundOutput[94]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U980 ( .s (n315), .b ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .a ({new_AGEMA_signal_14928, new_AGEMA_signal_14927, new_AGEMA_signal_14926, MixColumnsOutput[95]}), .c ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, new_AGEMA_signal_15703, RoundOutput[95]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U981 ( .s (n315), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .a ({new_AGEMA_signal_14904, new_AGEMA_signal_14903, new_AGEMA_signal_14902, MixColumnsOutput[96]}), .c ({new_AGEMA_signal_15708, new_AGEMA_signal_15707, new_AGEMA_signal_15706, RoundOutput[96]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U982 ( .s (n315), .b ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .a ({new_AGEMA_signal_15735, new_AGEMA_signal_15734, new_AGEMA_signal_15733, MixColumnsOutput[97]}), .c ({new_AGEMA_signal_16188, new_AGEMA_signal_16187, new_AGEMA_signal_16186, RoundOutput[97]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U983 ( .s (n315), .b ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .a ({new_AGEMA_signal_14838, new_AGEMA_signal_14837, new_AGEMA_signal_14836, MixColumnsOutput[98]}), .c ({new_AGEMA_signal_15711, new_AGEMA_signal_15710, new_AGEMA_signal_15709, RoundOutput[98]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U984 ( .s (n315), .b ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .a ({new_AGEMA_signal_15720, new_AGEMA_signal_15719, new_AGEMA_signal_15718, MixColumnsOutput[99]}), .c ({new_AGEMA_signal_16191, new_AGEMA_signal_16190, new_AGEMA_signal_16189, RoundOutput[99]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) U985 ( .s (n315), .b ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .a ({new_AGEMA_signal_15822, new_AGEMA_signal_15821, new_AGEMA_signal_15820, MixColumnsOutput[9]}), .c ({new_AGEMA_signal_16194, new_AGEMA_signal_16193, new_AGEMA_signal_16192, RoundOutput[9]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15474, new_AGEMA_signal_15473, new_AGEMA_signal_15472, RoundOutput[0]}), .a ({plaintext_s3[0], plaintext_s2[0], plaintext_s1[0], plaintext_s0[0]}), .c ({new_AGEMA_signal_16200, new_AGEMA_signal_16199, new_AGEMA_signal_16198, RoundReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16095, new_AGEMA_signal_16094, new_AGEMA_signal_16093, RoundOutput[1]}), .a ({plaintext_s3[1], plaintext_s2[1], plaintext_s1[1], plaintext_s0[1]}), .c ({new_AGEMA_signal_16722, new_AGEMA_signal_16721, new_AGEMA_signal_16720, RoundReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15567, new_AGEMA_signal_15566, new_AGEMA_signal_15565, RoundOutput[2]}), .a ({plaintext_s3[2], plaintext_s2[2], plaintext_s1[2], plaintext_s0[2]}), .c ({new_AGEMA_signal_16206, new_AGEMA_signal_16205, new_AGEMA_signal_16204, RoundReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16119, new_AGEMA_signal_16118, new_AGEMA_signal_16117, RoundOutput[3]}), .a ({plaintext_s3[3], plaintext_s2[3], plaintext_s1[3], plaintext_s0[3]}), .c ({new_AGEMA_signal_16728, new_AGEMA_signal_16727, new_AGEMA_signal_16726, RoundReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16134, new_AGEMA_signal_16133, new_AGEMA_signal_16132, RoundOutput[4]}), .a ({plaintext_s3[4], plaintext_s2[4], plaintext_s1[4], plaintext_s0[4]}), .c ({new_AGEMA_signal_16734, new_AGEMA_signal_16733, new_AGEMA_signal_16732, RoundReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15627, new_AGEMA_signal_15626, new_AGEMA_signal_15625, RoundOutput[5]}), .a ({plaintext_s3[5], plaintext_s2[5], plaintext_s1[5], plaintext_s0[5]}), .c ({new_AGEMA_signal_16212, new_AGEMA_signal_16211, new_AGEMA_signal_16210, RoundReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15648, new_AGEMA_signal_15647, new_AGEMA_signal_15646, RoundOutput[6]}), .a ({plaintext_s3[6], plaintext_s2[6], plaintext_s1[6], plaintext_s0[6]}), .c ({new_AGEMA_signal_16218, new_AGEMA_signal_16217, new_AGEMA_signal_16216, RoundReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15672, new_AGEMA_signal_15671, new_AGEMA_signal_15670, RoundOutput[7]}), .a ({plaintext_s3[7], plaintext_s2[7], plaintext_s1[7], plaintext_s0[7]}), .c ({new_AGEMA_signal_16224, new_AGEMA_signal_16223, new_AGEMA_signal_16222, RoundReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15693, new_AGEMA_signal_15692, new_AGEMA_signal_15691, RoundOutput[8]}), .a ({plaintext_s3[8], plaintext_s2[8], plaintext_s1[8], plaintext_s0[8]}), .c ({new_AGEMA_signal_16230, new_AGEMA_signal_16229, new_AGEMA_signal_16228, RoundReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16194, new_AGEMA_signal_16193, new_AGEMA_signal_16192, RoundOutput[9]}), .a ({plaintext_s3[9], plaintext_s2[9], plaintext_s1[9], plaintext_s0[9]}), .c ({new_AGEMA_signal_16740, new_AGEMA_signal_16739, new_AGEMA_signal_16738, RoundReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15495, new_AGEMA_signal_15494, new_AGEMA_signal_15493, RoundOutput[10]}), .a ({plaintext_s3[10], plaintext_s2[10], plaintext_s1[10], plaintext_s0[10]}), .c ({new_AGEMA_signal_16236, new_AGEMA_signal_16235, new_AGEMA_signal_16234, RoundReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16074, new_AGEMA_signal_16073, new_AGEMA_signal_16072, RoundOutput[11]}), .a ({plaintext_s3[11], plaintext_s2[11], plaintext_s1[11], plaintext_s0[11]}), .c ({new_AGEMA_signal_16746, new_AGEMA_signal_16745, new_AGEMA_signal_16744, RoundReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16086, new_AGEMA_signal_16085, new_AGEMA_signal_16084, RoundOutput[12]}), .a ({plaintext_s3[12], plaintext_s2[12], plaintext_s1[12], plaintext_s0[12]}), .c ({new_AGEMA_signal_16752, new_AGEMA_signal_16751, new_AGEMA_signal_16750, RoundReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15534, new_AGEMA_signal_15533, new_AGEMA_signal_15532, RoundOutput[13]}), .a ({plaintext_s3[13], plaintext_s2[13], plaintext_s1[13], plaintext_s0[13]}), .c ({new_AGEMA_signal_16242, new_AGEMA_signal_16241, new_AGEMA_signal_16240, RoundReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15537, new_AGEMA_signal_15536, new_AGEMA_signal_15535, RoundOutput[14]}), .a ({plaintext_s3[14], plaintext_s2[14], plaintext_s1[14], plaintext_s0[14]}), .c ({new_AGEMA_signal_16248, new_AGEMA_signal_16247, new_AGEMA_signal_16246, RoundReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15540, new_AGEMA_signal_15539, new_AGEMA_signal_15538, RoundOutput[15]}), .a ({plaintext_s3[15], plaintext_s2[15], plaintext_s1[15], plaintext_s0[15]}), .c ({new_AGEMA_signal_16254, new_AGEMA_signal_16253, new_AGEMA_signal_16252, RoundReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15543, new_AGEMA_signal_15542, new_AGEMA_signal_15541, RoundOutput[16]}), .a ({plaintext_s3[16], plaintext_s2[16], plaintext_s1[16], plaintext_s0[16]}), .c ({new_AGEMA_signal_16260, new_AGEMA_signal_16259, new_AGEMA_signal_16258, RoundReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16089, new_AGEMA_signal_16088, new_AGEMA_signal_16087, RoundOutput[17]}), .a ({plaintext_s3[17], plaintext_s2[17], plaintext_s1[17], plaintext_s0[17]}), .c ({new_AGEMA_signal_16758, new_AGEMA_signal_16757, new_AGEMA_signal_16756, RoundReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15546, new_AGEMA_signal_15545, new_AGEMA_signal_15544, RoundOutput[18]}), .a ({plaintext_s3[18], plaintext_s2[18], plaintext_s1[18], plaintext_s0[18]}), .c ({new_AGEMA_signal_16266, new_AGEMA_signal_16265, new_AGEMA_signal_16264, RoundReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16092, new_AGEMA_signal_16091, new_AGEMA_signal_16090, RoundOutput[19]}), .a ({plaintext_s3[19], plaintext_s2[19], plaintext_s1[19], plaintext_s0[19]}), .c ({new_AGEMA_signal_16764, new_AGEMA_signal_16763, new_AGEMA_signal_16762, RoundReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16098, new_AGEMA_signal_16097, new_AGEMA_signal_16096, RoundOutput[20]}), .a ({plaintext_s3[20], plaintext_s2[20], plaintext_s1[20], plaintext_s0[20]}), .c ({new_AGEMA_signal_16770, new_AGEMA_signal_16769, new_AGEMA_signal_16768, RoundReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15549, new_AGEMA_signal_15548, new_AGEMA_signal_15547, RoundOutput[21]}), .a ({plaintext_s3[21], plaintext_s2[21], plaintext_s1[21], plaintext_s0[21]}), .c ({new_AGEMA_signal_16272, new_AGEMA_signal_16271, new_AGEMA_signal_16270, RoundReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15552, new_AGEMA_signal_15551, new_AGEMA_signal_15550, RoundOutput[22]}), .a ({plaintext_s3[22], plaintext_s2[22], plaintext_s1[22], plaintext_s0[22]}), .c ({new_AGEMA_signal_16278, new_AGEMA_signal_16277, new_AGEMA_signal_16276, RoundReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15555, new_AGEMA_signal_15554, new_AGEMA_signal_15553, RoundOutput[23]}), .a ({plaintext_s3[23], plaintext_s2[23], plaintext_s1[23], plaintext_s0[23]}), .c ({new_AGEMA_signal_16284, new_AGEMA_signal_16283, new_AGEMA_signal_16282, RoundReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15558, new_AGEMA_signal_15557, new_AGEMA_signal_15556, RoundOutput[24]}), .a ({plaintext_s3[24], plaintext_s2[24], plaintext_s1[24], plaintext_s0[24]}), .c ({new_AGEMA_signal_16290, new_AGEMA_signal_16289, new_AGEMA_signal_16288, RoundReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16101, new_AGEMA_signal_16100, new_AGEMA_signal_16099, RoundOutput[25]}), .a ({plaintext_s3[25], plaintext_s2[25], plaintext_s1[25], plaintext_s0[25]}), .c ({new_AGEMA_signal_16776, new_AGEMA_signal_16775, new_AGEMA_signal_16774, RoundReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15561, new_AGEMA_signal_15560, new_AGEMA_signal_15559, RoundOutput[26]}), .a ({plaintext_s3[26], plaintext_s2[26], plaintext_s1[26], plaintext_s0[26]}), .c ({new_AGEMA_signal_16296, new_AGEMA_signal_16295, new_AGEMA_signal_16294, RoundReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16104, new_AGEMA_signal_16103, new_AGEMA_signal_16102, RoundOutput[27]}), .a ({plaintext_s3[27], plaintext_s2[27], plaintext_s1[27], plaintext_s0[27]}), .c ({new_AGEMA_signal_16782, new_AGEMA_signal_16781, new_AGEMA_signal_16780, RoundReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16107, new_AGEMA_signal_16106, new_AGEMA_signal_16105, RoundOutput[28]}), .a ({plaintext_s3[28], plaintext_s2[28], plaintext_s1[28], plaintext_s0[28]}), .c ({new_AGEMA_signal_16788, new_AGEMA_signal_16787, new_AGEMA_signal_16786, RoundReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15564, new_AGEMA_signal_15563, new_AGEMA_signal_15562, RoundOutput[29]}), .a ({plaintext_s3[29], plaintext_s2[29], plaintext_s1[29], plaintext_s0[29]}), .c ({new_AGEMA_signal_16302, new_AGEMA_signal_16301, new_AGEMA_signal_16300, RoundReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15570, new_AGEMA_signal_15569, new_AGEMA_signal_15568, RoundOutput[30]}), .a ({plaintext_s3[30], plaintext_s2[30], plaintext_s1[30], plaintext_s0[30]}), .c ({new_AGEMA_signal_16308, new_AGEMA_signal_16307, new_AGEMA_signal_16306, RoundReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15573, new_AGEMA_signal_15572, new_AGEMA_signal_15571, RoundOutput[31]}), .a ({plaintext_s3[31], plaintext_s2[31], plaintext_s1[31], plaintext_s0[31]}), .c ({new_AGEMA_signal_16314, new_AGEMA_signal_16313, new_AGEMA_signal_16312, RoundReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15576, new_AGEMA_signal_15575, new_AGEMA_signal_15574, RoundOutput[32]}), .a ({plaintext_s3[32], plaintext_s2[32], plaintext_s1[32], plaintext_s0[32]}), .c ({new_AGEMA_signal_16320, new_AGEMA_signal_16319, new_AGEMA_signal_16318, RoundReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16110, new_AGEMA_signal_16109, new_AGEMA_signal_16108, RoundOutput[33]}), .a ({plaintext_s3[33], plaintext_s2[33], plaintext_s1[33], plaintext_s0[33]}), .c ({new_AGEMA_signal_16794, new_AGEMA_signal_16793, new_AGEMA_signal_16792, RoundReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15579, new_AGEMA_signal_15578, new_AGEMA_signal_15577, RoundOutput[34]}), .a ({plaintext_s3[34], plaintext_s2[34], plaintext_s1[34], plaintext_s0[34]}), .c ({new_AGEMA_signal_16326, new_AGEMA_signal_16325, new_AGEMA_signal_16324, RoundReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16113, new_AGEMA_signal_16112, new_AGEMA_signal_16111, RoundOutput[35]}), .a ({plaintext_s3[35], plaintext_s2[35], plaintext_s1[35], plaintext_s0[35]}), .c ({new_AGEMA_signal_16800, new_AGEMA_signal_16799, new_AGEMA_signal_16798, RoundReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16116, new_AGEMA_signal_16115, new_AGEMA_signal_16114, RoundOutput[36]}), .a ({plaintext_s3[36], plaintext_s2[36], plaintext_s1[36], plaintext_s0[36]}), .c ({new_AGEMA_signal_16806, new_AGEMA_signal_16805, new_AGEMA_signal_16804, RoundReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15582, new_AGEMA_signal_15581, new_AGEMA_signal_15580, RoundOutput[37]}), .a ({plaintext_s3[37], plaintext_s2[37], plaintext_s1[37], plaintext_s0[37]}), .c ({new_AGEMA_signal_16332, new_AGEMA_signal_16331, new_AGEMA_signal_16330, RoundReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15585, new_AGEMA_signal_15584, new_AGEMA_signal_15583, RoundOutput[38]}), .a ({plaintext_s3[38], plaintext_s2[38], plaintext_s1[38], plaintext_s0[38]}), .c ({new_AGEMA_signal_16338, new_AGEMA_signal_16337, new_AGEMA_signal_16336, RoundReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15588, new_AGEMA_signal_15587, new_AGEMA_signal_15586, RoundOutput[39]}), .a ({plaintext_s3[39], plaintext_s2[39], plaintext_s1[39], plaintext_s0[39]}), .c ({new_AGEMA_signal_16344, new_AGEMA_signal_16343, new_AGEMA_signal_16342, RoundReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15591, new_AGEMA_signal_15590, new_AGEMA_signal_15589, RoundOutput[40]}), .a ({plaintext_s3[40], plaintext_s2[40], plaintext_s1[40], plaintext_s0[40]}), .c ({new_AGEMA_signal_16350, new_AGEMA_signal_16349, new_AGEMA_signal_16348, RoundReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16122, new_AGEMA_signal_16121, new_AGEMA_signal_16120, RoundOutput[41]}), .a ({plaintext_s3[41], plaintext_s2[41], plaintext_s1[41], plaintext_s0[41]}), .c ({new_AGEMA_signal_16812, new_AGEMA_signal_16811, new_AGEMA_signal_16810, RoundReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15594, new_AGEMA_signal_15593, new_AGEMA_signal_15592, RoundOutput[42]}), .a ({plaintext_s3[42], plaintext_s2[42], plaintext_s1[42], plaintext_s0[42]}), .c ({new_AGEMA_signal_16356, new_AGEMA_signal_16355, new_AGEMA_signal_16354, RoundReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16125, new_AGEMA_signal_16124, new_AGEMA_signal_16123, RoundOutput[43]}), .a ({plaintext_s3[43], plaintext_s2[43], plaintext_s1[43], plaintext_s0[43]}), .c ({new_AGEMA_signal_16818, new_AGEMA_signal_16817, new_AGEMA_signal_16816, RoundReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16128, new_AGEMA_signal_16127, new_AGEMA_signal_16126, RoundOutput[44]}), .a ({plaintext_s3[44], plaintext_s2[44], plaintext_s1[44], plaintext_s0[44]}), .c ({new_AGEMA_signal_16824, new_AGEMA_signal_16823, new_AGEMA_signal_16822, RoundReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15597, new_AGEMA_signal_15596, new_AGEMA_signal_15595, RoundOutput[45]}), .a ({plaintext_s3[45], plaintext_s2[45], plaintext_s1[45], plaintext_s0[45]}), .c ({new_AGEMA_signal_16362, new_AGEMA_signal_16361, new_AGEMA_signal_16360, RoundReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15600, new_AGEMA_signal_15599, new_AGEMA_signal_15598, RoundOutput[46]}), .a ({plaintext_s3[46], plaintext_s2[46], plaintext_s1[46], plaintext_s0[46]}), .c ({new_AGEMA_signal_16368, new_AGEMA_signal_16367, new_AGEMA_signal_16366, RoundReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15603, new_AGEMA_signal_15602, new_AGEMA_signal_15601, RoundOutput[47]}), .a ({plaintext_s3[47], plaintext_s2[47], plaintext_s1[47], plaintext_s0[47]}), .c ({new_AGEMA_signal_16374, new_AGEMA_signal_16373, new_AGEMA_signal_16372, RoundReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15606, new_AGEMA_signal_15605, new_AGEMA_signal_15604, RoundOutput[48]}), .a ({plaintext_s3[48], plaintext_s2[48], plaintext_s1[48], plaintext_s0[48]}), .c ({new_AGEMA_signal_16380, new_AGEMA_signal_16379, new_AGEMA_signal_16378, RoundReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16131, new_AGEMA_signal_16130, new_AGEMA_signal_16129, RoundOutput[49]}), .a ({plaintext_s3[49], plaintext_s2[49], plaintext_s1[49], plaintext_s0[49]}), .c ({new_AGEMA_signal_16830, new_AGEMA_signal_16829, new_AGEMA_signal_16828, RoundReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15609, new_AGEMA_signal_15608, new_AGEMA_signal_15607, RoundOutput[50]}), .a ({plaintext_s3[50], plaintext_s2[50], plaintext_s1[50], plaintext_s0[50]}), .c ({new_AGEMA_signal_16386, new_AGEMA_signal_16385, new_AGEMA_signal_16384, RoundReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16137, new_AGEMA_signal_16136, new_AGEMA_signal_16135, RoundOutput[51]}), .a ({plaintext_s3[51], plaintext_s2[51], plaintext_s1[51], plaintext_s0[51]}), .c ({new_AGEMA_signal_16836, new_AGEMA_signal_16835, new_AGEMA_signal_16834, RoundReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16140, new_AGEMA_signal_16139, new_AGEMA_signal_16138, RoundOutput[52]}), .a ({plaintext_s3[52], plaintext_s2[52], plaintext_s1[52], plaintext_s0[52]}), .c ({new_AGEMA_signal_16842, new_AGEMA_signal_16841, new_AGEMA_signal_16840, RoundReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15612, new_AGEMA_signal_15611, new_AGEMA_signal_15610, RoundOutput[53]}), .a ({plaintext_s3[53], plaintext_s2[53], plaintext_s1[53], plaintext_s0[53]}), .c ({new_AGEMA_signal_16392, new_AGEMA_signal_16391, new_AGEMA_signal_16390, RoundReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15615, new_AGEMA_signal_15614, new_AGEMA_signal_15613, RoundOutput[54]}), .a ({plaintext_s3[54], plaintext_s2[54], plaintext_s1[54], plaintext_s0[54]}), .c ({new_AGEMA_signal_16398, new_AGEMA_signal_16397, new_AGEMA_signal_16396, RoundReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15618, new_AGEMA_signal_15617, new_AGEMA_signal_15616, RoundOutput[55]}), .a ({plaintext_s3[55], plaintext_s2[55], plaintext_s1[55], plaintext_s0[55]}), .c ({new_AGEMA_signal_16404, new_AGEMA_signal_16403, new_AGEMA_signal_16402, RoundReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15621, new_AGEMA_signal_15620, new_AGEMA_signal_15619, RoundOutput[56]}), .a ({plaintext_s3[56], plaintext_s2[56], plaintext_s1[56], plaintext_s0[56]}), .c ({new_AGEMA_signal_16410, new_AGEMA_signal_16409, new_AGEMA_signal_16408, RoundReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16143, new_AGEMA_signal_16142, new_AGEMA_signal_16141, RoundOutput[57]}), .a ({plaintext_s3[57], plaintext_s2[57], plaintext_s1[57], plaintext_s0[57]}), .c ({new_AGEMA_signal_16848, new_AGEMA_signal_16847, new_AGEMA_signal_16846, RoundReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15624, new_AGEMA_signal_15623, new_AGEMA_signal_15622, RoundOutput[58]}), .a ({plaintext_s3[58], plaintext_s2[58], plaintext_s1[58], plaintext_s0[58]}), .c ({new_AGEMA_signal_16416, new_AGEMA_signal_16415, new_AGEMA_signal_16414, RoundReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16146, new_AGEMA_signal_16145, new_AGEMA_signal_16144, RoundOutput[59]}), .a ({plaintext_s3[59], plaintext_s2[59], plaintext_s1[59], plaintext_s0[59]}), .c ({new_AGEMA_signal_16854, new_AGEMA_signal_16853, new_AGEMA_signal_16852, RoundReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16149, new_AGEMA_signal_16148, new_AGEMA_signal_16147, RoundOutput[60]}), .a ({plaintext_s3[60], plaintext_s2[60], plaintext_s1[60], plaintext_s0[60]}), .c ({new_AGEMA_signal_16860, new_AGEMA_signal_16859, new_AGEMA_signal_16858, RoundReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15630, new_AGEMA_signal_15629, new_AGEMA_signal_15628, RoundOutput[61]}), .a ({plaintext_s3[61], plaintext_s2[61], plaintext_s1[61], plaintext_s0[61]}), .c ({new_AGEMA_signal_16422, new_AGEMA_signal_16421, new_AGEMA_signal_16420, RoundReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15633, new_AGEMA_signal_15632, new_AGEMA_signal_15631, RoundOutput[62]}), .a ({plaintext_s3[62], plaintext_s2[62], plaintext_s1[62], plaintext_s0[62]}), .c ({new_AGEMA_signal_16428, new_AGEMA_signal_16427, new_AGEMA_signal_16426, RoundReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15636, new_AGEMA_signal_15635, new_AGEMA_signal_15634, RoundOutput[63]}), .a ({plaintext_s3[63], plaintext_s2[63], plaintext_s1[63], plaintext_s0[63]}), .c ({new_AGEMA_signal_16434, new_AGEMA_signal_16433, new_AGEMA_signal_16432, RoundReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15639, new_AGEMA_signal_15638, new_AGEMA_signal_15637, RoundOutput[64]}), .a ({plaintext_s3[64], plaintext_s2[64], plaintext_s1[64], plaintext_s0[64]}), .c ({new_AGEMA_signal_16440, new_AGEMA_signal_16439, new_AGEMA_signal_16438, RoundReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16152, new_AGEMA_signal_16151, new_AGEMA_signal_16150, RoundOutput[65]}), .a ({plaintext_s3[65], plaintext_s2[65], plaintext_s1[65], plaintext_s0[65]}), .c ({new_AGEMA_signal_16866, new_AGEMA_signal_16865, new_AGEMA_signal_16864, RoundReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15642, new_AGEMA_signal_15641, new_AGEMA_signal_15640, RoundOutput[66]}), .a ({plaintext_s3[66], plaintext_s2[66], plaintext_s1[66], plaintext_s0[66]}), .c ({new_AGEMA_signal_16446, new_AGEMA_signal_16445, new_AGEMA_signal_16444, RoundReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16155, new_AGEMA_signal_16154, new_AGEMA_signal_16153, RoundOutput[67]}), .a ({plaintext_s3[67], plaintext_s2[67], plaintext_s1[67], plaintext_s0[67]}), .c ({new_AGEMA_signal_16872, new_AGEMA_signal_16871, new_AGEMA_signal_16870, RoundReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16158, new_AGEMA_signal_16157, new_AGEMA_signal_16156, RoundOutput[68]}), .a ({plaintext_s3[68], plaintext_s2[68], plaintext_s1[68], plaintext_s0[68]}), .c ({new_AGEMA_signal_16878, new_AGEMA_signal_16877, new_AGEMA_signal_16876, RoundReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15645, new_AGEMA_signal_15644, new_AGEMA_signal_15643, RoundOutput[69]}), .a ({plaintext_s3[69], plaintext_s2[69], plaintext_s1[69], plaintext_s0[69]}), .c ({new_AGEMA_signal_16452, new_AGEMA_signal_16451, new_AGEMA_signal_16450, RoundReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15651, new_AGEMA_signal_15650, new_AGEMA_signal_15649, RoundOutput[70]}), .a ({plaintext_s3[70], plaintext_s2[70], plaintext_s1[70], plaintext_s0[70]}), .c ({new_AGEMA_signal_16458, new_AGEMA_signal_16457, new_AGEMA_signal_16456, RoundReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15654, new_AGEMA_signal_15653, new_AGEMA_signal_15652, RoundOutput[71]}), .a ({plaintext_s3[71], plaintext_s2[71], plaintext_s1[71], plaintext_s0[71]}), .c ({new_AGEMA_signal_16464, new_AGEMA_signal_16463, new_AGEMA_signal_16462, RoundReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15657, new_AGEMA_signal_15656, new_AGEMA_signal_15655, RoundOutput[72]}), .a ({plaintext_s3[72], plaintext_s2[72], plaintext_s1[72], plaintext_s0[72]}), .c ({new_AGEMA_signal_16470, new_AGEMA_signal_16469, new_AGEMA_signal_16468, RoundReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16161, new_AGEMA_signal_16160, new_AGEMA_signal_16159, RoundOutput[73]}), .a ({plaintext_s3[73], plaintext_s2[73], plaintext_s1[73], plaintext_s0[73]}), .c ({new_AGEMA_signal_16884, new_AGEMA_signal_16883, new_AGEMA_signal_16882, RoundReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15660, new_AGEMA_signal_15659, new_AGEMA_signal_15658, RoundOutput[74]}), .a ({plaintext_s3[74], plaintext_s2[74], plaintext_s1[74], plaintext_s0[74]}), .c ({new_AGEMA_signal_16476, new_AGEMA_signal_16475, new_AGEMA_signal_16474, RoundReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16164, new_AGEMA_signal_16163, new_AGEMA_signal_16162, RoundOutput[75]}), .a ({plaintext_s3[75], plaintext_s2[75], plaintext_s1[75], plaintext_s0[75]}), .c ({new_AGEMA_signal_16890, new_AGEMA_signal_16889, new_AGEMA_signal_16888, RoundReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16167, new_AGEMA_signal_16166, new_AGEMA_signal_16165, RoundOutput[76]}), .a ({plaintext_s3[76], plaintext_s2[76], plaintext_s1[76], plaintext_s0[76]}), .c ({new_AGEMA_signal_16896, new_AGEMA_signal_16895, new_AGEMA_signal_16894, RoundReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15663, new_AGEMA_signal_15662, new_AGEMA_signal_15661, RoundOutput[77]}), .a ({plaintext_s3[77], plaintext_s2[77], plaintext_s1[77], plaintext_s0[77]}), .c ({new_AGEMA_signal_16482, new_AGEMA_signal_16481, new_AGEMA_signal_16480, RoundReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15666, new_AGEMA_signal_15665, new_AGEMA_signal_15664, RoundOutput[78]}), .a ({plaintext_s3[78], plaintext_s2[78], plaintext_s1[78], plaintext_s0[78]}), .c ({new_AGEMA_signal_16488, new_AGEMA_signal_16487, new_AGEMA_signal_16486, RoundReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15669, new_AGEMA_signal_15668, new_AGEMA_signal_15667, RoundOutput[79]}), .a ({plaintext_s3[79], plaintext_s2[79], plaintext_s1[79], plaintext_s0[79]}), .c ({new_AGEMA_signal_16494, new_AGEMA_signal_16493, new_AGEMA_signal_16492, RoundReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15675, new_AGEMA_signal_15674, new_AGEMA_signal_15673, RoundOutput[80]}), .a ({plaintext_s3[80], plaintext_s2[80], plaintext_s1[80], plaintext_s0[80]}), .c ({new_AGEMA_signal_16500, new_AGEMA_signal_16499, new_AGEMA_signal_16498, RoundReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16170, new_AGEMA_signal_16169, new_AGEMA_signal_16168, RoundOutput[81]}), .a ({plaintext_s3[81], plaintext_s2[81], plaintext_s1[81], plaintext_s0[81]}), .c ({new_AGEMA_signal_16902, new_AGEMA_signal_16901, new_AGEMA_signal_16900, RoundReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15678, new_AGEMA_signal_15677, new_AGEMA_signal_15676, RoundOutput[82]}), .a ({plaintext_s3[82], plaintext_s2[82], plaintext_s1[82], plaintext_s0[82]}), .c ({new_AGEMA_signal_16506, new_AGEMA_signal_16505, new_AGEMA_signal_16504, RoundReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16173, new_AGEMA_signal_16172, new_AGEMA_signal_16171, RoundOutput[83]}), .a ({plaintext_s3[83], plaintext_s2[83], plaintext_s1[83], plaintext_s0[83]}), .c ({new_AGEMA_signal_16908, new_AGEMA_signal_16907, new_AGEMA_signal_16906, RoundReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16176, new_AGEMA_signal_16175, new_AGEMA_signal_16174, RoundOutput[84]}), .a ({plaintext_s3[84], plaintext_s2[84], plaintext_s1[84], plaintext_s0[84]}), .c ({new_AGEMA_signal_16914, new_AGEMA_signal_16913, new_AGEMA_signal_16912, RoundReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15681, new_AGEMA_signal_15680, new_AGEMA_signal_15679, RoundOutput[85]}), .a ({plaintext_s3[85], plaintext_s2[85], plaintext_s1[85], plaintext_s0[85]}), .c ({new_AGEMA_signal_16512, new_AGEMA_signal_16511, new_AGEMA_signal_16510, RoundReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15684, new_AGEMA_signal_15683, new_AGEMA_signal_15682, RoundOutput[86]}), .a ({plaintext_s3[86], plaintext_s2[86], plaintext_s1[86], plaintext_s0[86]}), .c ({new_AGEMA_signal_16518, new_AGEMA_signal_16517, new_AGEMA_signal_16516, RoundReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15687, new_AGEMA_signal_15686, new_AGEMA_signal_15685, RoundOutput[87]}), .a ({plaintext_s3[87], plaintext_s2[87], plaintext_s1[87], plaintext_s0[87]}), .c ({new_AGEMA_signal_16524, new_AGEMA_signal_16523, new_AGEMA_signal_16522, RoundReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15690, new_AGEMA_signal_15689, new_AGEMA_signal_15688, RoundOutput[88]}), .a ({plaintext_s3[88], plaintext_s2[88], plaintext_s1[88], plaintext_s0[88]}), .c ({new_AGEMA_signal_16530, new_AGEMA_signal_16529, new_AGEMA_signal_16528, RoundReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16179, new_AGEMA_signal_16178, new_AGEMA_signal_16177, RoundOutput[89]}), .a ({plaintext_s3[89], plaintext_s2[89], plaintext_s1[89], plaintext_s0[89]}), .c ({new_AGEMA_signal_16920, new_AGEMA_signal_16919, new_AGEMA_signal_16918, RoundReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15696, new_AGEMA_signal_15695, new_AGEMA_signal_15694, RoundOutput[90]}), .a ({plaintext_s3[90], plaintext_s2[90], plaintext_s1[90], plaintext_s0[90]}), .c ({new_AGEMA_signal_16536, new_AGEMA_signal_16535, new_AGEMA_signal_16534, RoundReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16182, new_AGEMA_signal_16181, new_AGEMA_signal_16180, RoundOutput[91]}), .a ({plaintext_s3[91], plaintext_s2[91], plaintext_s1[91], plaintext_s0[91]}), .c ({new_AGEMA_signal_16926, new_AGEMA_signal_16925, new_AGEMA_signal_16924, RoundReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16185, new_AGEMA_signal_16184, new_AGEMA_signal_16183, RoundOutput[92]}), .a ({plaintext_s3[92], plaintext_s2[92], plaintext_s1[92], plaintext_s0[92]}), .c ({new_AGEMA_signal_16932, new_AGEMA_signal_16931, new_AGEMA_signal_16930, RoundReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15699, new_AGEMA_signal_15698, new_AGEMA_signal_15697, RoundOutput[93]}), .a ({plaintext_s3[93], plaintext_s2[93], plaintext_s1[93], plaintext_s0[93]}), .c ({new_AGEMA_signal_16542, new_AGEMA_signal_16541, new_AGEMA_signal_16540, RoundReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15702, new_AGEMA_signal_15701, new_AGEMA_signal_15700, RoundOutput[94]}), .a ({plaintext_s3[94], plaintext_s2[94], plaintext_s1[94], plaintext_s0[94]}), .c ({new_AGEMA_signal_16548, new_AGEMA_signal_16547, new_AGEMA_signal_16546, RoundReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15705, new_AGEMA_signal_15704, new_AGEMA_signal_15703, RoundOutput[95]}), .a ({plaintext_s3[95], plaintext_s2[95], plaintext_s1[95], plaintext_s0[95]}), .c ({new_AGEMA_signal_16554, new_AGEMA_signal_16553, new_AGEMA_signal_16552, RoundReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15708, new_AGEMA_signal_15707, new_AGEMA_signal_15706, RoundOutput[96]}), .a ({plaintext_s3[96], plaintext_s2[96], plaintext_s1[96], plaintext_s0[96]}), .c ({new_AGEMA_signal_16560, new_AGEMA_signal_16559, new_AGEMA_signal_16558, RoundReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16188, new_AGEMA_signal_16187, new_AGEMA_signal_16186, RoundOutput[97]}), .a ({plaintext_s3[97], plaintext_s2[97], plaintext_s1[97], plaintext_s0[97]}), .c ({new_AGEMA_signal_16938, new_AGEMA_signal_16937, new_AGEMA_signal_16936, RoundReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15711, new_AGEMA_signal_15710, new_AGEMA_signal_15709, RoundOutput[98]}), .a ({plaintext_s3[98], plaintext_s2[98], plaintext_s1[98], plaintext_s0[98]}), .c ({new_AGEMA_signal_16566, new_AGEMA_signal_16565, new_AGEMA_signal_16564, RoundReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16191, new_AGEMA_signal_16190, new_AGEMA_signal_16189, RoundOutput[99]}), .a ({plaintext_s3[99], plaintext_s2[99], plaintext_s1[99], plaintext_s0[99]}), .c ({new_AGEMA_signal_16944, new_AGEMA_signal_16943, new_AGEMA_signal_16942, RoundReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16053, new_AGEMA_signal_16052, new_AGEMA_signal_16051, RoundOutput[100]}), .a ({plaintext_s3[100], plaintext_s2[100], plaintext_s1[100], plaintext_s0[100]}), .c ({new_AGEMA_signal_16950, new_AGEMA_signal_16949, new_AGEMA_signal_16948, RoundReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15477, new_AGEMA_signal_15476, new_AGEMA_signal_15475, RoundOutput[101]}), .a ({plaintext_s3[101], plaintext_s2[101], plaintext_s1[101], plaintext_s0[101]}), .c ({new_AGEMA_signal_16572, new_AGEMA_signal_16571, new_AGEMA_signal_16570, RoundReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15480, new_AGEMA_signal_15479, new_AGEMA_signal_15478, RoundOutput[102]}), .a ({plaintext_s3[102], plaintext_s2[102], plaintext_s1[102], plaintext_s0[102]}), .c ({new_AGEMA_signal_16578, new_AGEMA_signal_16577, new_AGEMA_signal_16576, RoundReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15483, new_AGEMA_signal_15482, new_AGEMA_signal_15481, RoundOutput[103]}), .a ({plaintext_s3[103], plaintext_s2[103], plaintext_s1[103], plaintext_s0[103]}), .c ({new_AGEMA_signal_16584, new_AGEMA_signal_16583, new_AGEMA_signal_16582, RoundReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15486, new_AGEMA_signal_15485, new_AGEMA_signal_15484, RoundOutput[104]}), .a ({plaintext_s3[104], plaintext_s2[104], plaintext_s1[104], plaintext_s0[104]}), .c ({new_AGEMA_signal_16590, new_AGEMA_signal_16589, new_AGEMA_signal_16588, RoundReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16056, new_AGEMA_signal_16055, new_AGEMA_signal_16054, RoundOutput[105]}), .a ({plaintext_s3[105], plaintext_s2[105], plaintext_s1[105], plaintext_s0[105]}), .c ({new_AGEMA_signal_16956, new_AGEMA_signal_16955, new_AGEMA_signal_16954, RoundReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15489, new_AGEMA_signal_15488, new_AGEMA_signal_15487, RoundOutput[106]}), .a ({plaintext_s3[106], plaintext_s2[106], plaintext_s1[106], plaintext_s0[106]}), .c ({new_AGEMA_signal_16596, new_AGEMA_signal_16595, new_AGEMA_signal_16594, RoundReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16059, new_AGEMA_signal_16058, new_AGEMA_signal_16057, RoundOutput[107]}), .a ({plaintext_s3[107], plaintext_s2[107], plaintext_s1[107], plaintext_s0[107]}), .c ({new_AGEMA_signal_16962, new_AGEMA_signal_16961, new_AGEMA_signal_16960, RoundReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16062, new_AGEMA_signal_16061, new_AGEMA_signal_16060, RoundOutput[108]}), .a ({plaintext_s3[108], plaintext_s2[108], plaintext_s1[108], plaintext_s0[108]}), .c ({new_AGEMA_signal_16968, new_AGEMA_signal_16967, new_AGEMA_signal_16966, RoundReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15492, new_AGEMA_signal_15491, new_AGEMA_signal_15490, RoundOutput[109]}), .a ({plaintext_s3[109], plaintext_s2[109], plaintext_s1[109], plaintext_s0[109]}), .c ({new_AGEMA_signal_16602, new_AGEMA_signal_16601, new_AGEMA_signal_16600, RoundReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15498, new_AGEMA_signal_15497, new_AGEMA_signal_15496, RoundOutput[110]}), .a ({plaintext_s3[110], plaintext_s2[110], plaintext_s1[110], plaintext_s0[110]}), .c ({new_AGEMA_signal_16608, new_AGEMA_signal_16607, new_AGEMA_signal_16606, RoundReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15501, new_AGEMA_signal_15500, new_AGEMA_signal_15499, RoundOutput[111]}), .a ({plaintext_s3[111], plaintext_s2[111], plaintext_s1[111], plaintext_s0[111]}), .c ({new_AGEMA_signal_16614, new_AGEMA_signal_16613, new_AGEMA_signal_16612, RoundReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15504, new_AGEMA_signal_15503, new_AGEMA_signal_15502, RoundOutput[112]}), .a ({plaintext_s3[112], plaintext_s2[112], plaintext_s1[112], plaintext_s0[112]}), .c ({new_AGEMA_signal_16620, new_AGEMA_signal_16619, new_AGEMA_signal_16618, RoundReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16065, new_AGEMA_signal_16064, new_AGEMA_signal_16063, RoundOutput[113]}), .a ({plaintext_s3[113], plaintext_s2[113], plaintext_s1[113], plaintext_s0[113]}), .c ({new_AGEMA_signal_16974, new_AGEMA_signal_16973, new_AGEMA_signal_16972, RoundReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15507, new_AGEMA_signal_15506, new_AGEMA_signal_15505, RoundOutput[114]}), .a ({plaintext_s3[114], plaintext_s2[114], plaintext_s1[114], plaintext_s0[114]}), .c ({new_AGEMA_signal_16626, new_AGEMA_signal_16625, new_AGEMA_signal_16624, RoundReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16068, new_AGEMA_signal_16067, new_AGEMA_signal_16066, RoundOutput[115]}), .a ({plaintext_s3[115], plaintext_s2[115], plaintext_s1[115], plaintext_s0[115]}), .c ({new_AGEMA_signal_16980, new_AGEMA_signal_16979, new_AGEMA_signal_16978, RoundReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16071, new_AGEMA_signal_16070, new_AGEMA_signal_16069, RoundOutput[116]}), .a ({plaintext_s3[116], plaintext_s2[116], plaintext_s1[116], plaintext_s0[116]}), .c ({new_AGEMA_signal_16986, new_AGEMA_signal_16985, new_AGEMA_signal_16984, RoundReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15510, new_AGEMA_signal_15509, new_AGEMA_signal_15508, RoundOutput[117]}), .a ({plaintext_s3[117], plaintext_s2[117], plaintext_s1[117], plaintext_s0[117]}), .c ({new_AGEMA_signal_16632, new_AGEMA_signal_16631, new_AGEMA_signal_16630, RoundReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15513, new_AGEMA_signal_15512, new_AGEMA_signal_15511, RoundOutput[118]}), .a ({plaintext_s3[118], plaintext_s2[118], plaintext_s1[118], plaintext_s0[118]}), .c ({new_AGEMA_signal_16638, new_AGEMA_signal_16637, new_AGEMA_signal_16636, RoundReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15516, new_AGEMA_signal_15515, new_AGEMA_signal_15514, RoundOutput[119]}), .a ({plaintext_s3[119], plaintext_s2[119], plaintext_s1[119], plaintext_s0[119]}), .c ({new_AGEMA_signal_16644, new_AGEMA_signal_16643, new_AGEMA_signal_16642, RoundReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15519, new_AGEMA_signal_15518, new_AGEMA_signal_15517, RoundOutput[120]}), .a ({plaintext_s3[120], plaintext_s2[120], plaintext_s1[120], plaintext_s0[120]}), .c ({new_AGEMA_signal_16650, new_AGEMA_signal_16649, new_AGEMA_signal_16648, RoundReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16077, new_AGEMA_signal_16076, new_AGEMA_signal_16075, RoundOutput[121]}), .a ({plaintext_s3[121], plaintext_s2[121], plaintext_s1[121], plaintext_s0[121]}), .c ({new_AGEMA_signal_16992, new_AGEMA_signal_16991, new_AGEMA_signal_16990, RoundReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15522, new_AGEMA_signal_15521, new_AGEMA_signal_15520, RoundOutput[122]}), .a ({plaintext_s3[122], plaintext_s2[122], plaintext_s1[122], plaintext_s0[122]}), .c ({new_AGEMA_signal_16656, new_AGEMA_signal_16655, new_AGEMA_signal_16654, RoundReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16080, new_AGEMA_signal_16079, new_AGEMA_signal_16078, RoundOutput[123]}), .a ({plaintext_s3[123], plaintext_s2[123], plaintext_s1[123], plaintext_s0[123]}), .c ({new_AGEMA_signal_16998, new_AGEMA_signal_16997, new_AGEMA_signal_16996, RoundReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16083, new_AGEMA_signal_16082, new_AGEMA_signal_16081, RoundOutput[124]}), .a ({plaintext_s3[124], plaintext_s2[124], plaintext_s1[124], plaintext_s0[124]}), .c ({new_AGEMA_signal_17004, new_AGEMA_signal_17003, new_AGEMA_signal_17002, RoundReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15525, new_AGEMA_signal_15524, new_AGEMA_signal_15523, RoundOutput[125]}), .a ({plaintext_s3[125], plaintext_s2[125], plaintext_s1[125], plaintext_s0[125]}), .c ({new_AGEMA_signal_16662, new_AGEMA_signal_16661, new_AGEMA_signal_16660, RoundReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15528, new_AGEMA_signal_15527, new_AGEMA_signal_15526, RoundOutput[126]}), .a ({plaintext_s3[126], plaintext_s2[126], plaintext_s1[126], plaintext_s0[126]}), .c ({new_AGEMA_signal_16668, new_AGEMA_signal_16667, new_AGEMA_signal_16666, RoundReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15531, new_AGEMA_signal_15530, new_AGEMA_signal_15529, RoundOutput[127]}), .a ({plaintext_s3[127], plaintext_s2[127], plaintext_s1[127], plaintext_s0[127]}), .c ({new_AGEMA_signal_16674, new_AGEMA_signal_16673, new_AGEMA_signal_16672, RoundReg_Inst_ff_SDE_127_next_state}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, new_AGEMA_signal_9874, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_6399, new_AGEMA_signal_6398, new_AGEMA_signal_6397, SubBytesIns_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920]}), .c ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, new_AGEMA_signal_10588, SubBytesIns_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6939, new_AGEMA_signal_6938, new_AGEMA_signal_6937, SubBytesIns_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926]}), .c ({new_AGEMA_signal_9879, new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .b ({ciphertext_s3[0], ciphertext_s2[0], ciphertext_s1[0], ciphertext_s0[0]}), .clk (clk), .r ({Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932]}), .c ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, new_AGEMA_signal_9880, SubBytesIns_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_6411, new_AGEMA_signal_6410, new_AGEMA_signal_6409, SubBytesIns_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938]}), .c ({new_AGEMA_signal_10593, new_AGEMA_signal_10592, new_AGEMA_signal_10591, SubBytesIns_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6402, new_AGEMA_signal_6401, new_AGEMA_signal_6400, SubBytesIns_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944]}), .c ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6948, new_AGEMA_signal_6947, new_AGEMA_signal_6946, SubBytesIns_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950]}), .c ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886, SubBytesIns_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_6408, new_AGEMA_signal_6407, new_AGEMA_signal_6406, SubBytesIns_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956]}), .c ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, new_AGEMA_signal_10594, SubBytesIns_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, new_AGEMA_signal_10585, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_6420, new_AGEMA_signal_6419, new_AGEMA_signal_6418, SubBytesIns_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962]}), .c ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, new_AGEMA_signal_11281, SubBytesIns_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_6942, new_AGEMA_signal_6941, new_AGEMA_signal_6940, SubBytesIns_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968]}), .c ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, new_AGEMA_signal_10597, SubBytesIns_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_9876, new_AGEMA_signal_9875, new_AGEMA_signal_9874, SubBytesIns_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_6405, new_AGEMA_signal_6404, new_AGEMA_signal_6403, SubBytesIns_Inst_Sbox_0_T13}), .clk (clk), .r ({Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974]}), .c ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, new_AGEMA_signal_10600, SubBytesIns_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_9540, new_AGEMA_signal_9539, new_AGEMA_signal_9538, SubBytesIns_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6954, new_AGEMA_signal_6953, new_AGEMA_signal_6952, SubBytesIns_Inst_Sbox_0_T23}), .clk (clk), .r ({Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980]}), .c ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_9537, new_AGEMA_signal_9536, new_AGEMA_signal_9535, SubBytesIns_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_6414, new_AGEMA_signal_6413, new_AGEMA_signal_6412, SubBytesIns_Inst_Sbox_0_T19}), .clk (clk), .r ({Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986]}), .c ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, new_AGEMA_signal_9892, SubBytesIns_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_9873, new_AGEMA_signal_9872, new_AGEMA_signal_9871, SubBytesIns_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5829, new_AGEMA_signal_5828, new_AGEMA_signal_5827, SubBytesIns_Inst_Sbox_0_T3}), .clk (clk), .r ({Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992]}), .c ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, new_AGEMA_signal_10603, SubBytesIns_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_9534, new_AGEMA_signal_9533, new_AGEMA_signal_9532, SubBytesIns_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6417, new_AGEMA_signal_6416, new_AGEMA_signal_6415, SubBytesIns_Inst_Sbox_0_T22}), .clk (clk), .r ({Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998]}), .c ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_9531, new_AGEMA_signal_9530, new_AGEMA_signal_9529, SubBytesIns_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6951, new_AGEMA_signal_6950, new_AGEMA_signal_6949, SubBytesIns_Inst_Sbox_0_T20}), .clk (clk), .r ({Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004]}), .c ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, new_AGEMA_signal_9898, SubBytesIns_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_9870, new_AGEMA_signal_9869, new_AGEMA_signal_9868, SubBytesIns_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5823, new_AGEMA_signal_5822, new_AGEMA_signal_5821, SubBytesIns_Inst_Sbox_0_T1}), .clk (clk), .r ({Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010]}), .c ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_10587, new_AGEMA_signal_10586, new_AGEMA_signal_10585, SubBytesIns_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5832, new_AGEMA_signal_5831, new_AGEMA_signal_5830, SubBytesIns_Inst_Sbox_0_T4}), .clk (clk), .r ({Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016]}), .c ({new_AGEMA_signal_11286, new_AGEMA_signal_11285, new_AGEMA_signal_11284, SubBytesIns_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_9867, new_AGEMA_signal_9866, new_AGEMA_signal_9865, SubBytesIns_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5826, new_AGEMA_signal_5825, new_AGEMA_signal_5824, SubBytesIns_Inst_Sbox_0_T2}), .clk (clk), .r ({Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022]}), .c ({new_AGEMA_signal_10611, new_AGEMA_signal_10610, new_AGEMA_signal_10609, SubBytesIns_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_11286, new_AGEMA_signal_11285, new_AGEMA_signal_11284, SubBytesIns_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, new_AGEMA_signal_10588, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, new_AGEMA_signal_9880, SubBytesIns_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, new_AGEMA_signal_11287, SubBytesIns_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_9879, new_AGEMA_signal_9878, new_AGEMA_signal_9877, SubBytesIns_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, new_AGEMA_signal_10600, SubBytesIns_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, new_AGEMA_signal_11290, SubBytesIns_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_10599, new_AGEMA_signal_10598, new_AGEMA_signal_10597, SubBytesIns_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, new_AGEMA_signal_10603, SubBytesIns_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, new_AGEMA_signal_11293, SubBytesIns_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_10593, new_AGEMA_signal_10592, new_AGEMA_signal_10591, SubBytesIns_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11298, new_AGEMA_signal_11297, new_AGEMA_signal_11296, SubBytesIns_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_11286, new_AGEMA_signal_11285, new_AGEMA_signal_11284, SubBytesIns_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_11298, new_AGEMA_signal_11297, new_AGEMA_signal_11296, SubBytesIns_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_10590, new_AGEMA_signal_10589, new_AGEMA_signal_10588, SubBytesIns_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, new_AGEMA_signal_11290, SubBytesIns_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, new_AGEMA_signal_11875, SubBytesIns_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886, SubBytesIns_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_9897, new_AGEMA_signal_9896, new_AGEMA_signal_9895, SubBytesIns_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, new_AGEMA_signal_10615, SubBytesIns_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, new_AGEMA_signal_10594, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, new_AGEMA_signal_11281, SubBytesIns_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, new_AGEMA_signal_11878, SubBytesIns_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_11283, new_AGEMA_signal_11282, new_AGEMA_signal_11281, SubBytesIns_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, new_AGEMA_signal_11293, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, new_AGEMA_signal_11881, SubBytesIns_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_9900, new_AGEMA_signal_9899, new_AGEMA_signal_9898, SubBytesIns_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, new_AGEMA_signal_11287, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, new_AGEMA_signal_11884, SubBytesIns_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_9882, new_AGEMA_signal_9881, new_AGEMA_signal_9880, SubBytesIns_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_9888, new_AGEMA_signal_9887, new_AGEMA_signal_9886, SubBytesIns_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, new_AGEMA_signal_10618, SubBytesIns_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_9885, new_AGEMA_signal_9884, new_AGEMA_signal_9883, SubBytesIns_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12435, new_AGEMA_signal_12434, new_AGEMA_signal_12433, SubBytesIns_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_10596, new_AGEMA_signal_10595, new_AGEMA_signal_10594, SubBytesIns_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_10608, new_AGEMA_signal_10607, new_AGEMA_signal_10606, SubBytesIns_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, new_AGEMA_signal_11299, SubBytesIns_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_10602, new_AGEMA_signal_10601, new_AGEMA_signal_10600, SubBytesIns_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, new_AGEMA_signal_11302, SubBytesIns_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_9891, new_AGEMA_signal_9890, new_AGEMA_signal_9889, SubBytesIns_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12438, new_AGEMA_signal_12437, new_AGEMA_signal_12436, SubBytesIns_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_9894, new_AGEMA_signal_9893, new_AGEMA_signal_9892, SubBytesIns_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11307, new_AGEMA_signal_11306, new_AGEMA_signal_11305, SubBytesIns_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_10605, new_AGEMA_signal_10604, new_AGEMA_signal_10603, SubBytesIns_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, new_AGEMA_signal_10615, SubBytesIns_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_11310, new_AGEMA_signal_11309, new_AGEMA_signal_11308, SubBytesIns_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_10611, new_AGEMA_signal_10610, new_AGEMA_signal_10609, SubBytesIns_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_11295, new_AGEMA_signal_11294, new_AGEMA_signal_11293, SubBytesIns_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11889, new_AGEMA_signal_11888, new_AGEMA_signal_11887, SubBytesIns_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_11871, new_AGEMA_signal_11870, new_AGEMA_signal_11869, SubBytesIns_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_12441, new_AGEMA_signal_12440, new_AGEMA_signal_12439, SubBytesIns_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_10614, new_AGEMA_signal_10613, new_AGEMA_signal_10612, SubBytesIns_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, new_AGEMA_signal_11875, SubBytesIns_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, new_AGEMA_signal_12442, SubBytesIns_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_11292, new_AGEMA_signal_11291, new_AGEMA_signal_11290, SubBytesIns_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_10620, new_AGEMA_signal_10619, new_AGEMA_signal_10618, SubBytesIns_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, new_AGEMA_signal_11890, SubBytesIns_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_11310, new_AGEMA_signal_11309, new_AGEMA_signal_11308, SubBytesIns_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_11289, new_AGEMA_signal_11288, new_AGEMA_signal_11287, SubBytesIns_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11895, new_AGEMA_signal_11894, new_AGEMA_signal_11893, SubBytesIns_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_11304, new_AGEMA_signal_11303, new_AGEMA_signal_11302, SubBytesIns_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, new_AGEMA_signal_11878, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, new_AGEMA_signal_12445, SubBytesIns_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, new_AGEMA_signal_11881, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12450, new_AGEMA_signal_12449, new_AGEMA_signal_12448, SubBytesIns_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_11877, new_AGEMA_signal_11876, new_AGEMA_signal_11875, SubBytesIns_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_11880, new_AGEMA_signal_11879, new_AGEMA_signal_11878, SubBytesIns_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12453, new_AGEMA_signal_12452, new_AGEMA_signal_12451, SubBytesIns_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_10617, new_AGEMA_signal_10616, new_AGEMA_signal_10615, SubBytesIns_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_11883, new_AGEMA_signal_11882, new_AGEMA_signal_11881, SubBytesIns_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, new_AGEMA_signal_12454, SubBytesIns_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, new_AGEMA_signal_11884, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11301, new_AGEMA_signal_11300, new_AGEMA_signal_11299, SubBytesIns_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_12459, new_AGEMA_signal_12458, new_AGEMA_signal_12457, SubBytesIns_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_11886, new_AGEMA_signal_11885, new_AGEMA_signal_11884, SubBytesIns_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11307, new_AGEMA_signal_11306, new_AGEMA_signal_11305, SubBytesIns_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_12462, new_AGEMA_signal_12461, new_AGEMA_signal_12460, SubBytesIns_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12447, new_AGEMA_signal_12446, new_AGEMA_signal_12445, SubBytesIns_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_12438, new_AGEMA_signal_12437, new_AGEMA_signal_12436, SubBytesIns_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_12453, new_AGEMA_signal_12452, new_AGEMA_signal_12451, SubBytesIns_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_11889, new_AGEMA_signal_11888, new_AGEMA_signal_11887, SubBytesIns_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_12459, new_AGEMA_signal_12458, new_AGEMA_signal_12457, SubBytesIns_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12444, new_AGEMA_signal_12443, new_AGEMA_signal_12442, SubBytesIns_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_12441, new_AGEMA_signal_12440, new_AGEMA_signal_12439, SubBytesIns_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_11892, new_AGEMA_signal_11891, new_AGEMA_signal_11890, SubBytesIns_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_12450, new_AGEMA_signal_12449, new_AGEMA_signal_12448, SubBytesIns_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_12462, new_AGEMA_signal_12461, new_AGEMA_signal_12460, SubBytesIns_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_12435, new_AGEMA_signal_12434, new_AGEMA_signal_12433, SubBytesIns_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_12456, new_AGEMA_signal_12455, new_AGEMA_signal_12454, SubBytesIns_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_11874, new_AGEMA_signal_11873, new_AGEMA_signal_11872, SubBytesIns_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11895, new_AGEMA_signal_11894, new_AGEMA_signal_11893, SubBytesIns_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_6423, new_AGEMA_signal_6422, new_AGEMA_signal_6421, SubBytesIns_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028]}), .c ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, new_AGEMA_signal_10624, SubBytesIns_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6978, new_AGEMA_signal_6977, new_AGEMA_signal_6976, SubBytesIns_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034]}), .c ({new_AGEMA_signal_9915, new_AGEMA_signal_9914, new_AGEMA_signal_9913, SubBytesIns_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .b ({ciphertext_s3[8], ciphertext_s2[8], ciphertext_s1[8], ciphertext_s0[8]}), .clk (clk), .r ({Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040]}), .c ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, new_AGEMA_signal_9916, SubBytesIns_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_6435, new_AGEMA_signal_6434, new_AGEMA_signal_6433, SubBytesIns_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046]}), .c ({new_AGEMA_signal_10629, new_AGEMA_signal_10628, new_AGEMA_signal_10627, SubBytesIns_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6426, new_AGEMA_signal_6425, new_AGEMA_signal_6424, SubBytesIns_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052]}), .c ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6987, new_AGEMA_signal_6986, new_AGEMA_signal_6985, SubBytesIns_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058]}), .c ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922, SubBytesIns_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_6432, new_AGEMA_signal_6431, new_AGEMA_signal_6430, SubBytesIns_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064]}), .c ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, new_AGEMA_signal_10630, SubBytesIns_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, new_AGEMA_signal_10621, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_6444, new_AGEMA_signal_6443, new_AGEMA_signal_6442, SubBytesIns_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070]}), .c ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, new_AGEMA_signal_11311, SubBytesIns_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_6981, new_AGEMA_signal_6980, new_AGEMA_signal_6979, SubBytesIns_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076]}), .c ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, new_AGEMA_signal_10633, SubBytesIns_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_9912, new_AGEMA_signal_9911, new_AGEMA_signal_9910, SubBytesIns_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_6429, new_AGEMA_signal_6428, new_AGEMA_signal_6427, SubBytesIns_Inst_Sbox_1_T13}), .clk (clk), .r ({Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082]}), .c ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, new_AGEMA_signal_10636, SubBytesIns_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_9552, new_AGEMA_signal_9551, new_AGEMA_signal_9550, SubBytesIns_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6993, new_AGEMA_signal_6992, new_AGEMA_signal_6991, SubBytesIns_Inst_Sbox_1_T23}), .clk (clk), .r ({Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088]}), .c ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_9549, new_AGEMA_signal_9548, new_AGEMA_signal_9547, SubBytesIns_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_6438, new_AGEMA_signal_6437, new_AGEMA_signal_6436, SubBytesIns_Inst_Sbox_1_T19}), .clk (clk), .r ({Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094]}), .c ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, new_AGEMA_signal_9928, SubBytesIns_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_9909, new_AGEMA_signal_9908, new_AGEMA_signal_9907, SubBytesIns_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5859, new_AGEMA_signal_5858, new_AGEMA_signal_5857, SubBytesIns_Inst_Sbox_1_T3}), .clk (clk), .r ({Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100]}), .c ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, new_AGEMA_signal_10639, SubBytesIns_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_9546, new_AGEMA_signal_9545, new_AGEMA_signal_9544, SubBytesIns_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6441, new_AGEMA_signal_6440, new_AGEMA_signal_6439, SubBytesIns_Inst_Sbox_1_T22}), .clk (clk), .r ({Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106]}), .c ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_9543, new_AGEMA_signal_9542, new_AGEMA_signal_9541, SubBytesIns_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6990, new_AGEMA_signal_6989, new_AGEMA_signal_6988, SubBytesIns_Inst_Sbox_1_T20}), .clk (clk), .r ({Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112]}), .c ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, new_AGEMA_signal_9934, SubBytesIns_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_9906, new_AGEMA_signal_9905, new_AGEMA_signal_9904, SubBytesIns_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5853, new_AGEMA_signal_5852, new_AGEMA_signal_5851, SubBytesIns_Inst_Sbox_1_T1}), .clk (clk), .r ({Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118]}), .c ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_10623, new_AGEMA_signal_10622, new_AGEMA_signal_10621, SubBytesIns_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5862, new_AGEMA_signal_5861, new_AGEMA_signal_5860, SubBytesIns_Inst_Sbox_1_T4}), .clk (clk), .r ({Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124]}), .c ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, new_AGEMA_signal_11314, SubBytesIns_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_9903, new_AGEMA_signal_9902, new_AGEMA_signal_9901, SubBytesIns_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5856, new_AGEMA_signal_5855, new_AGEMA_signal_5854, SubBytesIns_Inst_Sbox_1_T2}), .clk (clk), .r ({Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130]}), .c ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, new_AGEMA_signal_10645, SubBytesIns_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, new_AGEMA_signal_11314, SubBytesIns_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, new_AGEMA_signal_10624, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, new_AGEMA_signal_9916, SubBytesIns_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, new_AGEMA_signal_11317, SubBytesIns_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_9915, new_AGEMA_signal_9914, new_AGEMA_signal_9913, SubBytesIns_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, new_AGEMA_signal_10636, SubBytesIns_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_11322, new_AGEMA_signal_11321, new_AGEMA_signal_11320, SubBytesIns_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_10635, new_AGEMA_signal_10634, new_AGEMA_signal_10633, SubBytesIns_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, new_AGEMA_signal_10639, SubBytesIns_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, new_AGEMA_signal_11323, SubBytesIns_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_10629, new_AGEMA_signal_10628, new_AGEMA_signal_10627, SubBytesIns_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, new_AGEMA_signal_11326, SubBytesIns_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_11316, new_AGEMA_signal_11315, new_AGEMA_signal_11314, SubBytesIns_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_11328, new_AGEMA_signal_11327, new_AGEMA_signal_11326, SubBytesIns_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_10626, new_AGEMA_signal_10625, new_AGEMA_signal_10624, SubBytesIns_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_11322, new_AGEMA_signal_11321, new_AGEMA_signal_11320, SubBytesIns_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, new_AGEMA_signal_11902, SubBytesIns_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922, SubBytesIns_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_9933, new_AGEMA_signal_9932, new_AGEMA_signal_9931, SubBytesIns_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, new_AGEMA_signal_10651, SubBytesIns_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, new_AGEMA_signal_10630, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, new_AGEMA_signal_11311, SubBytesIns_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, new_AGEMA_signal_11905, SubBytesIns_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_11313, new_AGEMA_signal_11312, new_AGEMA_signal_11311, SubBytesIns_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, new_AGEMA_signal_11323, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, new_AGEMA_signal_11908, SubBytesIns_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_9936, new_AGEMA_signal_9935, new_AGEMA_signal_9934, SubBytesIns_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, new_AGEMA_signal_11317, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, new_AGEMA_signal_11911, SubBytesIns_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_9918, new_AGEMA_signal_9917, new_AGEMA_signal_9916, SubBytesIns_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_9924, new_AGEMA_signal_9923, new_AGEMA_signal_9922, SubBytesIns_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, new_AGEMA_signal_10654, SubBytesIns_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_9921, new_AGEMA_signal_9920, new_AGEMA_signal_9919, SubBytesIns_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, new_AGEMA_signal_12466, SubBytesIns_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_10632, new_AGEMA_signal_10631, new_AGEMA_signal_10630, SubBytesIns_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_10644, new_AGEMA_signal_10643, new_AGEMA_signal_10642, SubBytesIns_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11331, new_AGEMA_signal_11330, new_AGEMA_signal_11329, SubBytesIns_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_10638, new_AGEMA_signal_10637, new_AGEMA_signal_10636, SubBytesIns_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, new_AGEMA_signal_11332, SubBytesIns_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_9927, new_AGEMA_signal_9926, new_AGEMA_signal_9925, SubBytesIns_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12471, new_AGEMA_signal_12470, new_AGEMA_signal_12469, SubBytesIns_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_9930, new_AGEMA_signal_9929, new_AGEMA_signal_9928, SubBytesIns_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11337, new_AGEMA_signal_11336, new_AGEMA_signal_11335, SubBytesIns_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_10641, new_AGEMA_signal_10640, new_AGEMA_signal_10639, SubBytesIns_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, new_AGEMA_signal_10651, SubBytesIns_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, new_AGEMA_signal_11338, SubBytesIns_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_10647, new_AGEMA_signal_10646, new_AGEMA_signal_10645, SubBytesIns_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_11325, new_AGEMA_signal_11324, new_AGEMA_signal_11323, SubBytesIns_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, new_AGEMA_signal_11914, SubBytesIns_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_11898, new_AGEMA_signal_11897, new_AGEMA_signal_11896, SubBytesIns_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_12474, new_AGEMA_signal_12473, new_AGEMA_signal_12472, SubBytesIns_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_10650, new_AGEMA_signal_10649, new_AGEMA_signal_10648, SubBytesIns_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, new_AGEMA_signal_11902, SubBytesIns_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_12477, new_AGEMA_signal_12476, new_AGEMA_signal_12475, SubBytesIns_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_11322, new_AGEMA_signal_11321, new_AGEMA_signal_11320, SubBytesIns_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_10656, new_AGEMA_signal_10655, new_AGEMA_signal_10654, SubBytesIns_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_11919, new_AGEMA_signal_11918, new_AGEMA_signal_11917, SubBytesIns_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_11340, new_AGEMA_signal_11339, new_AGEMA_signal_11338, SubBytesIns_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_11319, new_AGEMA_signal_11318, new_AGEMA_signal_11317, SubBytesIns_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, new_AGEMA_signal_11920, SubBytesIns_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_11334, new_AGEMA_signal_11333, new_AGEMA_signal_11332, SubBytesIns_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, new_AGEMA_signal_11905, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, new_AGEMA_signal_12478, SubBytesIns_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, new_AGEMA_signal_11908, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12483, new_AGEMA_signal_12482, new_AGEMA_signal_12481, SubBytesIns_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_11904, new_AGEMA_signal_11903, new_AGEMA_signal_11902, SubBytesIns_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_11907, new_AGEMA_signal_11906, new_AGEMA_signal_11905, SubBytesIns_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12486, new_AGEMA_signal_12485, new_AGEMA_signal_12484, SubBytesIns_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_10653, new_AGEMA_signal_10652, new_AGEMA_signal_10651, SubBytesIns_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_11910, new_AGEMA_signal_11909, new_AGEMA_signal_11908, SubBytesIns_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12489, new_AGEMA_signal_12488, new_AGEMA_signal_12487, SubBytesIns_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, new_AGEMA_signal_11911, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11331, new_AGEMA_signal_11330, new_AGEMA_signal_11329, SubBytesIns_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, new_AGEMA_signal_12490, SubBytesIns_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_11913, new_AGEMA_signal_11912, new_AGEMA_signal_11911, SubBytesIns_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11337, new_AGEMA_signal_11336, new_AGEMA_signal_11335, SubBytesIns_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_12495, new_AGEMA_signal_12494, new_AGEMA_signal_12493, SubBytesIns_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12480, new_AGEMA_signal_12479, new_AGEMA_signal_12478, SubBytesIns_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_12471, new_AGEMA_signal_12470, new_AGEMA_signal_12469, SubBytesIns_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_12486, new_AGEMA_signal_12485, new_AGEMA_signal_12484, SubBytesIns_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_11916, new_AGEMA_signal_11915, new_AGEMA_signal_11914, SubBytesIns_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_12492, new_AGEMA_signal_12491, new_AGEMA_signal_12490, SubBytesIns_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12477, new_AGEMA_signal_12476, new_AGEMA_signal_12475, SubBytesIns_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_12474, new_AGEMA_signal_12473, new_AGEMA_signal_12472, SubBytesIns_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_11919, new_AGEMA_signal_11918, new_AGEMA_signal_11917, SubBytesIns_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_12483, new_AGEMA_signal_12482, new_AGEMA_signal_12481, SubBytesIns_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_12495, new_AGEMA_signal_12494, new_AGEMA_signal_12493, SubBytesIns_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_12468, new_AGEMA_signal_12467, new_AGEMA_signal_12466, SubBytesIns_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_12489, new_AGEMA_signal_12488, new_AGEMA_signal_12487, SubBytesIns_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_11901, new_AGEMA_signal_11900, new_AGEMA_signal_11899, SubBytesIns_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11922, new_AGEMA_signal_11921, new_AGEMA_signal_11920, SubBytesIns_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_6447, new_AGEMA_signal_6446, new_AGEMA_signal_6445, SubBytesIns_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136]}), .c ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, new_AGEMA_signal_10660, SubBytesIns_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_7017, new_AGEMA_signal_7016, new_AGEMA_signal_7015, SubBytesIns_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142]}), .c ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .b ({ciphertext_s3[16], ciphertext_s2[16], ciphertext_s1[16], ciphertext_s0[16]}), .clk (clk), .r ({Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148]}), .c ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, new_AGEMA_signal_9952, SubBytesIns_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_6459, new_AGEMA_signal_6458, new_AGEMA_signal_6457, SubBytesIns_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154]}), .c ({new_AGEMA_signal_10665, new_AGEMA_signal_10664, new_AGEMA_signal_10663, SubBytesIns_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6450, new_AGEMA_signal_6449, new_AGEMA_signal_6448, SubBytesIns_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160]}), .c ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7026, new_AGEMA_signal_7025, new_AGEMA_signal_7024, SubBytesIns_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166]}), .c ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958, SubBytesIns_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_6456, new_AGEMA_signal_6455, new_AGEMA_signal_6454, SubBytesIns_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172]}), .c ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, new_AGEMA_signal_10666, SubBytesIns_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, new_AGEMA_signal_10657, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_6468, new_AGEMA_signal_6467, new_AGEMA_signal_6466, SubBytesIns_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178]}), .c ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, new_AGEMA_signal_11341, SubBytesIns_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_7020, new_AGEMA_signal_7019, new_AGEMA_signal_7018, SubBytesIns_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184]}), .c ({new_AGEMA_signal_10671, new_AGEMA_signal_10670, new_AGEMA_signal_10669, SubBytesIns_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_9948, new_AGEMA_signal_9947, new_AGEMA_signal_9946, SubBytesIns_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_6453, new_AGEMA_signal_6452, new_AGEMA_signal_6451, SubBytesIns_Inst_Sbox_2_T13}), .clk (clk), .r ({Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190]}), .c ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, new_AGEMA_signal_10672, SubBytesIns_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_9564, new_AGEMA_signal_9563, new_AGEMA_signal_9562, SubBytesIns_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_7032, new_AGEMA_signal_7031, new_AGEMA_signal_7030, SubBytesIns_Inst_Sbox_2_T23}), .clk (clk), .r ({Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196]}), .c ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_9561, new_AGEMA_signal_9560, new_AGEMA_signal_9559, SubBytesIns_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_6462, new_AGEMA_signal_6461, new_AGEMA_signal_6460, SubBytesIns_Inst_Sbox_2_T19}), .clk (clk), .r ({Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202]}), .c ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, new_AGEMA_signal_9964, SubBytesIns_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_9945, new_AGEMA_signal_9944, new_AGEMA_signal_9943, SubBytesIns_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5889, new_AGEMA_signal_5888, new_AGEMA_signal_5887, SubBytesIns_Inst_Sbox_2_T3}), .clk (clk), .r ({Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208]}), .c ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, new_AGEMA_signal_10675, SubBytesIns_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_9558, new_AGEMA_signal_9557, new_AGEMA_signal_9556, SubBytesIns_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6465, new_AGEMA_signal_6464, new_AGEMA_signal_6463, SubBytesIns_Inst_Sbox_2_T22}), .clk (clk), .r ({Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214]}), .c ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_9555, new_AGEMA_signal_9554, new_AGEMA_signal_9553, SubBytesIns_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_7029, new_AGEMA_signal_7028, new_AGEMA_signal_7027, SubBytesIns_Inst_Sbox_2_T20}), .clk (clk), .r ({Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220]}), .c ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, new_AGEMA_signal_9970, SubBytesIns_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_9942, new_AGEMA_signal_9941, new_AGEMA_signal_9940, SubBytesIns_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5883, new_AGEMA_signal_5882, new_AGEMA_signal_5881, SubBytesIns_Inst_Sbox_2_T1}), .clk (clk), .r ({Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226]}), .c ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_10659, new_AGEMA_signal_10658, new_AGEMA_signal_10657, SubBytesIns_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5892, new_AGEMA_signal_5891, new_AGEMA_signal_5890, SubBytesIns_Inst_Sbox_2_T4}), .clk (clk), .r ({Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232]}), .c ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, new_AGEMA_signal_11344, SubBytesIns_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_9939, new_AGEMA_signal_9938, new_AGEMA_signal_9937, SubBytesIns_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5886, new_AGEMA_signal_5885, new_AGEMA_signal_5884, SubBytesIns_Inst_Sbox_2_T2}), .clk (clk), .r ({Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238]}), .c ({new_AGEMA_signal_10683, new_AGEMA_signal_10682, new_AGEMA_signal_10681, SubBytesIns_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, new_AGEMA_signal_11344, SubBytesIns_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, new_AGEMA_signal_10660, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, new_AGEMA_signal_9952, SubBytesIns_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, new_AGEMA_signal_11347, SubBytesIns_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_9951, new_AGEMA_signal_9950, new_AGEMA_signal_9949, SubBytesIns_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, new_AGEMA_signal_10672, SubBytesIns_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, new_AGEMA_signal_11350, SubBytesIns_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_10671, new_AGEMA_signal_10670, new_AGEMA_signal_10669, SubBytesIns_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, new_AGEMA_signal_10675, SubBytesIns_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, new_AGEMA_signal_11353, SubBytesIns_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_10665, new_AGEMA_signal_10664, new_AGEMA_signal_10663, SubBytesIns_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, new_AGEMA_signal_11356, SubBytesIns_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_11346, new_AGEMA_signal_11345, new_AGEMA_signal_11344, SubBytesIns_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_11358, new_AGEMA_signal_11357, new_AGEMA_signal_11356, SubBytesIns_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_10662, new_AGEMA_signal_10661, new_AGEMA_signal_10660, SubBytesIns_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, new_AGEMA_signal_11350, SubBytesIns_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, new_AGEMA_signal_11929, SubBytesIns_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958, SubBytesIns_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_9969, new_AGEMA_signal_9968, new_AGEMA_signal_9967, SubBytesIns_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, new_AGEMA_signal_10687, SubBytesIns_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, new_AGEMA_signal_10666, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, new_AGEMA_signal_11341, SubBytesIns_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, new_AGEMA_signal_11932, SubBytesIns_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_11343, new_AGEMA_signal_11342, new_AGEMA_signal_11341, SubBytesIns_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, new_AGEMA_signal_11353, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, new_AGEMA_signal_11935, SubBytesIns_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_9972, new_AGEMA_signal_9971, new_AGEMA_signal_9970, SubBytesIns_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, new_AGEMA_signal_11347, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, new_AGEMA_signal_11938, SubBytesIns_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_9954, new_AGEMA_signal_9953, new_AGEMA_signal_9952, SubBytesIns_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_9960, new_AGEMA_signal_9959, new_AGEMA_signal_9958, SubBytesIns_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, new_AGEMA_signal_10690, SubBytesIns_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_9957, new_AGEMA_signal_9956, new_AGEMA_signal_9955, SubBytesIns_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12501, new_AGEMA_signal_12500, new_AGEMA_signal_12499, SubBytesIns_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_10668, new_AGEMA_signal_10667, new_AGEMA_signal_10666, SubBytesIns_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_10680, new_AGEMA_signal_10679, new_AGEMA_signal_10678, SubBytesIns_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11361, new_AGEMA_signal_11360, new_AGEMA_signal_11359, SubBytesIns_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_10674, new_AGEMA_signal_10673, new_AGEMA_signal_10672, SubBytesIns_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, new_AGEMA_signal_11362, SubBytesIns_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_9963, new_AGEMA_signal_9962, new_AGEMA_signal_9961, SubBytesIns_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, new_AGEMA_signal_12502, SubBytesIns_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_9966, new_AGEMA_signal_9965, new_AGEMA_signal_9964, SubBytesIns_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11367, new_AGEMA_signal_11366, new_AGEMA_signal_11365, SubBytesIns_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_10677, new_AGEMA_signal_10676, new_AGEMA_signal_10675, SubBytesIns_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, new_AGEMA_signal_10687, SubBytesIns_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, new_AGEMA_signal_11368, SubBytesIns_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_10683, new_AGEMA_signal_10682, new_AGEMA_signal_10681, SubBytesIns_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_11355, new_AGEMA_signal_11354, new_AGEMA_signal_11353, SubBytesIns_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11943, new_AGEMA_signal_11942, new_AGEMA_signal_11941, SubBytesIns_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_11925, new_AGEMA_signal_11924, new_AGEMA_signal_11923, SubBytesIns_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_12507, new_AGEMA_signal_12506, new_AGEMA_signal_12505, SubBytesIns_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_10686, new_AGEMA_signal_10685, new_AGEMA_signal_10684, SubBytesIns_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, new_AGEMA_signal_11929, SubBytesIns_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_12510, new_AGEMA_signal_12509, new_AGEMA_signal_12508, SubBytesIns_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_11352, new_AGEMA_signal_11351, new_AGEMA_signal_11350, SubBytesIns_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_10692, new_AGEMA_signal_10691, new_AGEMA_signal_10690, SubBytesIns_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, new_AGEMA_signal_11944, SubBytesIns_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_11370, new_AGEMA_signal_11369, new_AGEMA_signal_11368, SubBytesIns_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_11349, new_AGEMA_signal_11348, new_AGEMA_signal_11347, SubBytesIns_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11949, new_AGEMA_signal_11948, new_AGEMA_signal_11947, SubBytesIns_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_11364, new_AGEMA_signal_11363, new_AGEMA_signal_11362, SubBytesIns_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, new_AGEMA_signal_11932, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12513, new_AGEMA_signal_12512, new_AGEMA_signal_12511, SubBytesIns_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, new_AGEMA_signal_11935, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, new_AGEMA_signal_12514, SubBytesIns_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_11931, new_AGEMA_signal_11930, new_AGEMA_signal_11929, SubBytesIns_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_11934, new_AGEMA_signal_11933, new_AGEMA_signal_11932, SubBytesIns_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12519, new_AGEMA_signal_12518, new_AGEMA_signal_12517, SubBytesIns_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_10689, new_AGEMA_signal_10688, new_AGEMA_signal_10687, SubBytesIns_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_11937, new_AGEMA_signal_11936, new_AGEMA_signal_11935, SubBytesIns_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12522, new_AGEMA_signal_12521, new_AGEMA_signal_12520, SubBytesIns_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, new_AGEMA_signal_11938, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11361, new_AGEMA_signal_11360, new_AGEMA_signal_11359, SubBytesIns_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_12525, new_AGEMA_signal_12524, new_AGEMA_signal_12523, SubBytesIns_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_11940, new_AGEMA_signal_11939, new_AGEMA_signal_11938, SubBytesIns_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11367, new_AGEMA_signal_11366, new_AGEMA_signal_11365, SubBytesIns_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, new_AGEMA_signal_12526, SubBytesIns_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12513, new_AGEMA_signal_12512, new_AGEMA_signal_12511, SubBytesIns_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_12504, new_AGEMA_signal_12503, new_AGEMA_signal_12502, SubBytesIns_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_12519, new_AGEMA_signal_12518, new_AGEMA_signal_12517, SubBytesIns_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_11943, new_AGEMA_signal_11942, new_AGEMA_signal_11941, SubBytesIns_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_12525, new_AGEMA_signal_12524, new_AGEMA_signal_12523, SubBytesIns_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12510, new_AGEMA_signal_12509, new_AGEMA_signal_12508, SubBytesIns_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_12507, new_AGEMA_signal_12506, new_AGEMA_signal_12505, SubBytesIns_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_11946, new_AGEMA_signal_11945, new_AGEMA_signal_11944, SubBytesIns_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_12516, new_AGEMA_signal_12515, new_AGEMA_signal_12514, SubBytesIns_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_12528, new_AGEMA_signal_12527, new_AGEMA_signal_12526, SubBytesIns_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_12501, new_AGEMA_signal_12500, new_AGEMA_signal_12499, SubBytesIns_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_12522, new_AGEMA_signal_12521, new_AGEMA_signal_12520, SubBytesIns_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_11928, new_AGEMA_signal_11927, new_AGEMA_signal_11926, SubBytesIns_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11949, new_AGEMA_signal_11948, new_AGEMA_signal_11947, SubBytesIns_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_6471, new_AGEMA_signal_6470, new_AGEMA_signal_6469, SubBytesIns_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244]}), .c ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, new_AGEMA_signal_10696, SubBytesIns_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_7056, new_AGEMA_signal_7055, new_AGEMA_signal_7054, SubBytesIns_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250]}), .c ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .b ({ciphertext_s3[24], ciphertext_s2[24], ciphertext_s1[24], ciphertext_s0[24]}), .clk (clk), .r ({Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256]}), .c ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, new_AGEMA_signal_9988, SubBytesIns_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_6483, new_AGEMA_signal_6482, new_AGEMA_signal_6481, SubBytesIns_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262]}), .c ({new_AGEMA_signal_10701, new_AGEMA_signal_10700, new_AGEMA_signal_10699, SubBytesIns_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6474, new_AGEMA_signal_6473, new_AGEMA_signal_6472, SubBytesIns_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268]}), .c ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7065, new_AGEMA_signal_7064, new_AGEMA_signal_7063, SubBytesIns_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274]}), .c ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994, SubBytesIns_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_6480, new_AGEMA_signal_6479, new_AGEMA_signal_6478, SubBytesIns_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280]}), .c ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, new_AGEMA_signal_10702, SubBytesIns_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, new_AGEMA_signal_10693, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_6492, new_AGEMA_signal_6491, new_AGEMA_signal_6490, SubBytesIns_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286]}), .c ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, new_AGEMA_signal_11371, SubBytesIns_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_7059, new_AGEMA_signal_7058, new_AGEMA_signal_7057, SubBytesIns_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292]}), .c ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, new_AGEMA_signal_10705, SubBytesIns_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_9984, new_AGEMA_signal_9983, new_AGEMA_signal_9982, SubBytesIns_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_6477, new_AGEMA_signal_6476, new_AGEMA_signal_6475, SubBytesIns_Inst_Sbox_3_T13}), .clk (clk), .r ({Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298]}), .c ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, new_AGEMA_signal_10708, SubBytesIns_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_9576, new_AGEMA_signal_9575, new_AGEMA_signal_9574, SubBytesIns_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_7071, new_AGEMA_signal_7070, new_AGEMA_signal_7069, SubBytesIns_Inst_Sbox_3_T23}), .clk (clk), .r ({Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304]}), .c ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_9573, new_AGEMA_signal_9572, new_AGEMA_signal_9571, SubBytesIns_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_6486, new_AGEMA_signal_6485, new_AGEMA_signal_6484, SubBytesIns_Inst_Sbox_3_T19}), .clk (clk), .r ({Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310]}), .c ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, new_AGEMA_signal_10000, SubBytesIns_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_9981, new_AGEMA_signal_9980, new_AGEMA_signal_9979, SubBytesIns_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5919, new_AGEMA_signal_5918, new_AGEMA_signal_5917, SubBytesIns_Inst_Sbox_3_T3}), .clk (clk), .r ({Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316]}), .c ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, new_AGEMA_signal_10711, SubBytesIns_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_9570, new_AGEMA_signal_9569, new_AGEMA_signal_9568, SubBytesIns_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6489, new_AGEMA_signal_6488, new_AGEMA_signal_6487, SubBytesIns_Inst_Sbox_3_T22}), .clk (clk), .r ({Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322]}), .c ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_9567, new_AGEMA_signal_9566, new_AGEMA_signal_9565, SubBytesIns_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_7068, new_AGEMA_signal_7067, new_AGEMA_signal_7066, SubBytesIns_Inst_Sbox_3_T20}), .clk (clk), .r ({Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328]}), .c ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006, SubBytesIns_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_9978, new_AGEMA_signal_9977, new_AGEMA_signal_9976, SubBytesIns_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5913, new_AGEMA_signal_5912, new_AGEMA_signal_5911, SubBytesIns_Inst_Sbox_3_T1}), .clk (clk), .r ({Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334]}), .c ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_10695, new_AGEMA_signal_10694, new_AGEMA_signal_10693, SubBytesIns_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5922, new_AGEMA_signal_5921, new_AGEMA_signal_5920, SubBytesIns_Inst_Sbox_3_T4}), .clk (clk), .r ({Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340]}), .c ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, new_AGEMA_signal_11374, SubBytesIns_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_9975, new_AGEMA_signal_9974, new_AGEMA_signal_9973, SubBytesIns_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5916, new_AGEMA_signal_5915, new_AGEMA_signal_5914, SubBytesIns_Inst_Sbox_3_T2}), .clk (clk), .r ({Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346]}), .c ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, new_AGEMA_signal_10717, SubBytesIns_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, new_AGEMA_signal_11374, SubBytesIns_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, new_AGEMA_signal_10696, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, new_AGEMA_signal_9988, SubBytesIns_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, new_AGEMA_signal_11377, SubBytesIns_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_9987, new_AGEMA_signal_9986, new_AGEMA_signal_9985, SubBytesIns_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, new_AGEMA_signal_10708, SubBytesIns_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, new_AGEMA_signal_11380, SubBytesIns_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_10707, new_AGEMA_signal_10706, new_AGEMA_signal_10705, SubBytesIns_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, new_AGEMA_signal_10711, SubBytesIns_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, new_AGEMA_signal_11383, SubBytesIns_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_10701, new_AGEMA_signal_10700, new_AGEMA_signal_10699, SubBytesIns_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, new_AGEMA_signal_11386, SubBytesIns_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_11376, new_AGEMA_signal_11375, new_AGEMA_signal_11374, SubBytesIns_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_11388, new_AGEMA_signal_11387, new_AGEMA_signal_11386, SubBytesIns_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_10698, new_AGEMA_signal_10697, new_AGEMA_signal_10696, SubBytesIns_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, new_AGEMA_signal_11380, SubBytesIns_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, new_AGEMA_signal_11956, SubBytesIns_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994, SubBytesIns_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_10005, new_AGEMA_signal_10004, new_AGEMA_signal_10003, SubBytesIns_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, new_AGEMA_signal_10723, SubBytesIns_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, new_AGEMA_signal_10702, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, new_AGEMA_signal_11371, SubBytesIns_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, new_AGEMA_signal_11959, SubBytesIns_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_11373, new_AGEMA_signal_11372, new_AGEMA_signal_11371, SubBytesIns_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, new_AGEMA_signal_11383, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, new_AGEMA_signal_11962, SubBytesIns_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_10008, new_AGEMA_signal_10007, new_AGEMA_signal_10006, SubBytesIns_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, new_AGEMA_signal_11377, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, new_AGEMA_signal_11965, SubBytesIns_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_9990, new_AGEMA_signal_9989, new_AGEMA_signal_9988, SubBytesIns_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_9996, new_AGEMA_signal_9995, new_AGEMA_signal_9994, SubBytesIns_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, new_AGEMA_signal_10726, SubBytesIns_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_9993, new_AGEMA_signal_9992, new_AGEMA_signal_9991, SubBytesIns_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12534, new_AGEMA_signal_12533, new_AGEMA_signal_12532, SubBytesIns_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_10704, new_AGEMA_signal_10703, new_AGEMA_signal_10702, SubBytesIns_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_10716, new_AGEMA_signal_10715, new_AGEMA_signal_10714, SubBytesIns_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, new_AGEMA_signal_11389, SubBytesIns_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_10710, new_AGEMA_signal_10709, new_AGEMA_signal_10708, SubBytesIns_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, new_AGEMA_signal_11392, SubBytesIns_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_9999, new_AGEMA_signal_9998, new_AGEMA_signal_9997, SubBytesIns_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12537, new_AGEMA_signal_12536, new_AGEMA_signal_12535, SubBytesIns_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_10002, new_AGEMA_signal_10001, new_AGEMA_signal_10000, SubBytesIns_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11397, new_AGEMA_signal_11396, new_AGEMA_signal_11395, SubBytesIns_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_10713, new_AGEMA_signal_10712, new_AGEMA_signal_10711, SubBytesIns_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, new_AGEMA_signal_10723, SubBytesIns_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, new_AGEMA_signal_11398, SubBytesIns_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_10719, new_AGEMA_signal_10718, new_AGEMA_signal_10717, SubBytesIns_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_11385, new_AGEMA_signal_11384, new_AGEMA_signal_11383, SubBytesIns_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, new_AGEMA_signal_11968, SubBytesIns_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_11952, new_AGEMA_signal_11951, new_AGEMA_signal_11950, SubBytesIns_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, new_AGEMA_signal_12538, SubBytesIns_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_10722, new_AGEMA_signal_10721, new_AGEMA_signal_10720, SubBytesIns_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, new_AGEMA_signal_11956, SubBytesIns_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_12543, new_AGEMA_signal_12542, new_AGEMA_signal_12541, SubBytesIns_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_11382, new_AGEMA_signal_11381, new_AGEMA_signal_11380, SubBytesIns_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_10728, new_AGEMA_signal_10727, new_AGEMA_signal_10726, SubBytesIns_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, new_AGEMA_signal_11971, SubBytesIns_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_11400, new_AGEMA_signal_11399, new_AGEMA_signal_11398, SubBytesIns_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_11379, new_AGEMA_signal_11378, new_AGEMA_signal_11377, SubBytesIns_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, new_AGEMA_signal_11974, SubBytesIns_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_11394, new_AGEMA_signal_11393, new_AGEMA_signal_11392, SubBytesIns_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, new_AGEMA_signal_11959, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12546, new_AGEMA_signal_12545, new_AGEMA_signal_12544, SubBytesIns_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, new_AGEMA_signal_11962, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12549, new_AGEMA_signal_12548, new_AGEMA_signal_12547, SubBytesIns_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_11958, new_AGEMA_signal_11957, new_AGEMA_signal_11956, SubBytesIns_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_11961, new_AGEMA_signal_11960, new_AGEMA_signal_11959, SubBytesIns_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, new_AGEMA_signal_12550, SubBytesIns_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_10725, new_AGEMA_signal_10724, new_AGEMA_signal_10723, SubBytesIns_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_11964, new_AGEMA_signal_11963, new_AGEMA_signal_11962, SubBytesIns_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12555, new_AGEMA_signal_12554, new_AGEMA_signal_12553, SubBytesIns_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, new_AGEMA_signal_11965, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11391, new_AGEMA_signal_11390, new_AGEMA_signal_11389, SubBytesIns_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_12558, new_AGEMA_signal_12557, new_AGEMA_signal_12556, SubBytesIns_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_11967, new_AGEMA_signal_11966, new_AGEMA_signal_11965, SubBytesIns_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11397, new_AGEMA_signal_11396, new_AGEMA_signal_11395, SubBytesIns_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_12561, new_AGEMA_signal_12560, new_AGEMA_signal_12559, SubBytesIns_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12546, new_AGEMA_signal_12545, new_AGEMA_signal_12544, SubBytesIns_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_12537, new_AGEMA_signal_12536, new_AGEMA_signal_12535, SubBytesIns_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_12552, new_AGEMA_signal_12551, new_AGEMA_signal_12550, SubBytesIns_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_11970, new_AGEMA_signal_11969, new_AGEMA_signal_11968, SubBytesIns_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_12558, new_AGEMA_signal_12557, new_AGEMA_signal_12556, SubBytesIns_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12543, new_AGEMA_signal_12542, new_AGEMA_signal_12541, SubBytesIns_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_12540, new_AGEMA_signal_12539, new_AGEMA_signal_12538, SubBytesIns_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_11973, new_AGEMA_signal_11972, new_AGEMA_signal_11971, SubBytesIns_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_12549, new_AGEMA_signal_12548, new_AGEMA_signal_12547, SubBytesIns_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_12561, new_AGEMA_signal_12560, new_AGEMA_signal_12559, SubBytesIns_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_12534, new_AGEMA_signal_12533, new_AGEMA_signal_12532, SubBytesIns_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_12555, new_AGEMA_signal_12554, new_AGEMA_signal_12553, SubBytesIns_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_11955, new_AGEMA_signal_11954, new_AGEMA_signal_11953, SubBytesIns_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11976, new_AGEMA_signal_11975, new_AGEMA_signal_11974, SubBytesIns_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M46_U1 ( .a ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_6495, new_AGEMA_signal_6494, new_AGEMA_signal_6493, SubBytesIns_Inst_Sbox_4_T6}), .clk (clk), .r ({Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352]}), .c ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, new_AGEMA_signal_10732, SubBytesIns_Inst_Sbox_4_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M47_U1 ( .a ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_7095, new_AGEMA_signal_7094, new_AGEMA_signal_7093, SubBytesIns_Inst_Sbox_4_T8}), .clk (clk), .r ({Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358]}), .c ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_4_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M48_U1 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .b ({ciphertext_s3[32], ciphertext_s2[32], ciphertext_s1[32], ciphertext_s0[32]}), .clk (clk), .r ({Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364]}), .c ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, new_AGEMA_signal_10024, SubBytesIns_Inst_Sbox_4_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M49_U1 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_6507, new_AGEMA_signal_6506, new_AGEMA_signal_6505, SubBytesIns_Inst_Sbox_4_T16}), .clk (clk), .r ({Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370]}), .c ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, new_AGEMA_signal_10735, SubBytesIns_Inst_Sbox_4_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M50_U1 ( .a ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_6498, new_AGEMA_signal_6497, new_AGEMA_signal_6496, SubBytesIns_Inst_Sbox_4_T9}), .clk (clk), .r ({Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376]}), .c ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_4_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M51_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_7104, new_AGEMA_signal_7103, new_AGEMA_signal_7102, SubBytesIns_Inst_Sbox_4_T17}), .clk (clk), .r ({Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382]}), .c ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030, SubBytesIns_Inst_Sbox_4_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M52_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_6504, new_AGEMA_signal_6503, new_AGEMA_signal_6502, SubBytesIns_Inst_Sbox_4_T15}), .clk (clk), .r ({Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388]}), .c ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, new_AGEMA_signal_10738, SubBytesIns_Inst_Sbox_4_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M53_U1 ( .a ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, new_AGEMA_signal_10729, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_6516, new_AGEMA_signal_6515, new_AGEMA_signal_6514, SubBytesIns_Inst_Sbox_4_T27}), .clk (clk), .r ({Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394]}), .c ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, new_AGEMA_signal_11401, SubBytesIns_Inst_Sbox_4_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M54_U1 ( .a ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_7098, new_AGEMA_signal_7097, new_AGEMA_signal_7096, SubBytesIns_Inst_Sbox_4_T10}), .clk (clk), .r ({Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400]}), .c ({new_AGEMA_signal_10743, new_AGEMA_signal_10742, new_AGEMA_signal_10741, SubBytesIns_Inst_Sbox_4_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M55_U1 ( .a ({new_AGEMA_signal_10020, new_AGEMA_signal_10019, new_AGEMA_signal_10018, SubBytesIns_Inst_Sbox_4_M44}), .b ({new_AGEMA_signal_6501, new_AGEMA_signal_6500, new_AGEMA_signal_6499, SubBytesIns_Inst_Sbox_4_T13}), .clk (clk), .r ({Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406]}), .c ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, new_AGEMA_signal_10744, SubBytesIns_Inst_Sbox_4_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M56_U1 ( .a ({new_AGEMA_signal_9588, new_AGEMA_signal_9587, new_AGEMA_signal_9586, SubBytesIns_Inst_Sbox_4_M40}), .b ({new_AGEMA_signal_7110, new_AGEMA_signal_7109, new_AGEMA_signal_7108, SubBytesIns_Inst_Sbox_4_T23}), .clk (clk), .r ({Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412]}), .c ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_4_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M57_U1 ( .a ({new_AGEMA_signal_9585, new_AGEMA_signal_9584, new_AGEMA_signal_9583, SubBytesIns_Inst_Sbox_4_M39}), .b ({new_AGEMA_signal_6510, new_AGEMA_signal_6509, new_AGEMA_signal_6508, SubBytesIns_Inst_Sbox_4_T19}), .clk (clk), .r ({Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418]}), .c ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, new_AGEMA_signal_10036, SubBytesIns_Inst_Sbox_4_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M58_U1 ( .a ({new_AGEMA_signal_10017, new_AGEMA_signal_10016, new_AGEMA_signal_10015, SubBytesIns_Inst_Sbox_4_M43}), .b ({new_AGEMA_signal_5949, new_AGEMA_signal_5948, new_AGEMA_signal_5947, SubBytesIns_Inst_Sbox_4_T3}), .clk (clk), .r ({Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424]}), .c ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, new_AGEMA_signal_10747, SubBytesIns_Inst_Sbox_4_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M59_U1 ( .a ({new_AGEMA_signal_9582, new_AGEMA_signal_9581, new_AGEMA_signal_9580, SubBytesIns_Inst_Sbox_4_M38}), .b ({new_AGEMA_signal_6513, new_AGEMA_signal_6512, new_AGEMA_signal_6511, SubBytesIns_Inst_Sbox_4_T22}), .clk (clk), .r ({Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430]}), .c ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_4_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M60_U1 ( .a ({new_AGEMA_signal_9579, new_AGEMA_signal_9578, new_AGEMA_signal_9577, SubBytesIns_Inst_Sbox_4_M37}), .b ({new_AGEMA_signal_7107, new_AGEMA_signal_7106, new_AGEMA_signal_7105, SubBytesIns_Inst_Sbox_4_T20}), .clk (clk), .r ({Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436]}), .c ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, new_AGEMA_signal_10042, SubBytesIns_Inst_Sbox_4_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M61_U1 ( .a ({new_AGEMA_signal_10014, new_AGEMA_signal_10013, new_AGEMA_signal_10012, SubBytesIns_Inst_Sbox_4_M42}), .b ({new_AGEMA_signal_5943, new_AGEMA_signal_5942, new_AGEMA_signal_5941, SubBytesIns_Inst_Sbox_4_T1}), .clk (clk), .r ({Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442]}), .c ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M62_U1 ( .a ({new_AGEMA_signal_10731, new_AGEMA_signal_10730, new_AGEMA_signal_10729, SubBytesIns_Inst_Sbox_4_M45}), .b ({new_AGEMA_signal_5952, new_AGEMA_signal_5951, new_AGEMA_signal_5950, SubBytesIns_Inst_Sbox_4_T4}), .clk (clk), .r ({Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448]}), .c ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, new_AGEMA_signal_11404, SubBytesIns_Inst_Sbox_4_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_AND_M63_U1 ( .a ({new_AGEMA_signal_10011, new_AGEMA_signal_10010, new_AGEMA_signal_10009, SubBytesIns_Inst_Sbox_4_M41}), .b ({new_AGEMA_signal_5946, new_AGEMA_signal_5945, new_AGEMA_signal_5944, SubBytesIns_Inst_Sbox_4_T2}), .clk (clk), .r ({Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454]}), .c ({new_AGEMA_signal_10755, new_AGEMA_signal_10754, new_AGEMA_signal_10753, SubBytesIns_Inst_Sbox_4_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L0_U1 ( .a ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}), .b ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, new_AGEMA_signal_11404, SubBytesIns_Inst_Sbox_4_M62}), .c ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L1_U1 ( .a ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_4_M56}), .c ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L2_U1 ( .a ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, new_AGEMA_signal_10732, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, new_AGEMA_signal_10024, SubBytesIns_Inst_Sbox_4_M48}), .c ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, new_AGEMA_signal_11407, SubBytesIns_Inst_Sbox_4_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L3_U1 ( .a ({new_AGEMA_signal_10023, new_AGEMA_signal_10022, new_AGEMA_signal_10021, SubBytesIns_Inst_Sbox_4_M47}), .b ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, new_AGEMA_signal_10744, SubBytesIns_Inst_Sbox_4_M55}), .c ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, new_AGEMA_signal_11410, SubBytesIns_Inst_Sbox_4_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L4_U1 ( .a ({new_AGEMA_signal_10743, new_AGEMA_signal_10742, new_AGEMA_signal_10741, SubBytesIns_Inst_Sbox_4_M54}), .b ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, new_AGEMA_signal_10747, SubBytesIns_Inst_Sbox_4_M58}), .c ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, new_AGEMA_signal_11413, SubBytesIns_Inst_Sbox_4_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L5_U1 ( .a ({new_AGEMA_signal_10737, new_AGEMA_signal_10736, new_AGEMA_signal_10735, SubBytesIns_Inst_Sbox_4_M49}), .b ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, new_AGEMA_signal_11416, SubBytesIns_Inst_Sbox_4_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L6_U1 ( .a ({new_AGEMA_signal_11406, new_AGEMA_signal_11405, new_AGEMA_signal_11404, SubBytesIns_Inst_Sbox_4_M62}), .b ({new_AGEMA_signal_11418, new_AGEMA_signal_11417, new_AGEMA_signal_11416, SubBytesIns_Inst_Sbox_4_L5}), .c ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L7_U1 ( .a ({new_AGEMA_signal_10734, new_AGEMA_signal_10733, new_AGEMA_signal_10732, SubBytesIns_Inst_Sbox_4_M46}), .b ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, new_AGEMA_signal_11410, SubBytesIns_Inst_Sbox_4_L3}), .c ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, new_AGEMA_signal_11983, SubBytesIns_Inst_Sbox_4_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L8_U1 ( .a ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030, SubBytesIns_Inst_Sbox_4_M51}), .b ({new_AGEMA_signal_10041, new_AGEMA_signal_10040, new_AGEMA_signal_10039, SubBytesIns_Inst_Sbox_4_M59}), .c ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, new_AGEMA_signal_10759, SubBytesIns_Inst_Sbox_4_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L9_U1 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, new_AGEMA_signal_10738, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, new_AGEMA_signal_11401, SubBytesIns_Inst_Sbox_4_M53}), .c ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, new_AGEMA_signal_11986, SubBytesIns_Inst_Sbox_4_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L10_U1 ( .a ({new_AGEMA_signal_11403, new_AGEMA_signal_11402, new_AGEMA_signal_11401, SubBytesIns_Inst_Sbox_4_M53}), .b ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, new_AGEMA_signal_11413, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, new_AGEMA_signal_11989, SubBytesIns_Inst_Sbox_4_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L11_U1 ( .a ({new_AGEMA_signal_10044, new_AGEMA_signal_10043, new_AGEMA_signal_10042, SubBytesIns_Inst_Sbox_4_M60}), .b ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, new_AGEMA_signal_11407, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, new_AGEMA_signal_11992, SubBytesIns_Inst_Sbox_4_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L12_U1 ( .a ({new_AGEMA_signal_10026, new_AGEMA_signal_10025, new_AGEMA_signal_10024, SubBytesIns_Inst_Sbox_4_M48}), .b ({new_AGEMA_signal_10032, new_AGEMA_signal_10031, new_AGEMA_signal_10030, SubBytesIns_Inst_Sbox_4_M51}), .c ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, new_AGEMA_signal_10762, SubBytesIns_Inst_Sbox_4_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L13_U1 ( .a ({new_AGEMA_signal_10029, new_AGEMA_signal_10028, new_AGEMA_signal_10027, SubBytesIns_Inst_Sbox_4_M50}), .b ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_12567, new_AGEMA_signal_12566, new_AGEMA_signal_12565, SubBytesIns_Inst_Sbox_4_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L14_U1 ( .a ({new_AGEMA_signal_10740, new_AGEMA_signal_10739, new_AGEMA_signal_10738, SubBytesIns_Inst_Sbox_4_M52}), .b ({new_AGEMA_signal_10752, new_AGEMA_signal_10751, new_AGEMA_signal_10750, SubBytesIns_Inst_Sbox_4_M61}), .c ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, new_AGEMA_signal_11419, SubBytesIns_Inst_Sbox_4_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L15_U1 ( .a ({new_AGEMA_signal_10746, new_AGEMA_signal_10745, new_AGEMA_signal_10744, SubBytesIns_Inst_Sbox_4_M55}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, new_AGEMA_signal_11422, SubBytesIns_Inst_Sbox_4_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L16_U1 ( .a ({new_AGEMA_signal_10035, new_AGEMA_signal_10034, new_AGEMA_signal_10033, SubBytesIns_Inst_Sbox_4_M56}), .b ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}), .c ({new_AGEMA_signal_12570, new_AGEMA_signal_12569, new_AGEMA_signal_12568, SubBytesIns_Inst_Sbox_4_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L17_U1 ( .a ({new_AGEMA_signal_10038, new_AGEMA_signal_10037, new_AGEMA_signal_10036, SubBytesIns_Inst_Sbox_4_M57}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_11427, new_AGEMA_signal_11426, new_AGEMA_signal_11425, SubBytesIns_Inst_Sbox_4_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L18_U1 ( .a ({new_AGEMA_signal_10749, new_AGEMA_signal_10748, new_AGEMA_signal_10747, SubBytesIns_Inst_Sbox_4_M58}), .b ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, new_AGEMA_signal_10759, SubBytesIns_Inst_Sbox_4_L8}), .c ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, new_AGEMA_signal_11428, SubBytesIns_Inst_Sbox_4_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L19_U1 ( .a ({new_AGEMA_signal_10755, new_AGEMA_signal_10754, new_AGEMA_signal_10753, SubBytesIns_Inst_Sbox_4_M63}), .b ({new_AGEMA_signal_11415, new_AGEMA_signal_11414, new_AGEMA_signal_11413, SubBytesIns_Inst_Sbox_4_L4}), .c ({new_AGEMA_signal_11997, new_AGEMA_signal_11996, new_AGEMA_signal_11995, SubBytesIns_Inst_Sbox_4_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L20_U1 ( .a ({new_AGEMA_signal_11979, new_AGEMA_signal_11978, new_AGEMA_signal_11977, SubBytesIns_Inst_Sbox_4_L0}), .b ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .c ({new_AGEMA_signal_12573, new_AGEMA_signal_12572, new_AGEMA_signal_12571, SubBytesIns_Inst_Sbox_4_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L21_U1 ( .a ({new_AGEMA_signal_10758, new_AGEMA_signal_10757, new_AGEMA_signal_10756, SubBytesIns_Inst_Sbox_4_L1}), .b ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, new_AGEMA_signal_11983, SubBytesIns_Inst_Sbox_4_L7}), .c ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, new_AGEMA_signal_12574, SubBytesIns_Inst_Sbox_4_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L22_U1 ( .a ({new_AGEMA_signal_11412, new_AGEMA_signal_11411, new_AGEMA_signal_11410, SubBytesIns_Inst_Sbox_4_L3}), .b ({new_AGEMA_signal_10764, new_AGEMA_signal_10763, new_AGEMA_signal_10762, SubBytesIns_Inst_Sbox_4_L12}), .c ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, new_AGEMA_signal_11998, SubBytesIns_Inst_Sbox_4_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L23_U1 ( .a ({new_AGEMA_signal_11430, new_AGEMA_signal_11429, new_AGEMA_signal_11428, SubBytesIns_Inst_Sbox_4_L18}), .b ({new_AGEMA_signal_11409, new_AGEMA_signal_11408, new_AGEMA_signal_11407, SubBytesIns_Inst_Sbox_4_L2}), .c ({new_AGEMA_signal_12003, new_AGEMA_signal_12002, new_AGEMA_signal_12001, SubBytesIns_Inst_Sbox_4_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L24_U1 ( .a ({new_AGEMA_signal_11424, new_AGEMA_signal_11423, new_AGEMA_signal_11422, SubBytesIns_Inst_Sbox_4_L15}), .b ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, new_AGEMA_signal_11986, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_12579, new_AGEMA_signal_12578, new_AGEMA_signal_12577, SubBytesIns_Inst_Sbox_4_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L25_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, new_AGEMA_signal_11989, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_12582, new_AGEMA_signal_12581, new_AGEMA_signal_12580, SubBytesIns_Inst_Sbox_4_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L26_U1 ( .a ({new_AGEMA_signal_11985, new_AGEMA_signal_11984, new_AGEMA_signal_11983, SubBytesIns_Inst_Sbox_4_L7}), .b ({new_AGEMA_signal_11988, new_AGEMA_signal_11987, new_AGEMA_signal_11986, SubBytesIns_Inst_Sbox_4_L9}), .c ({new_AGEMA_signal_12585, new_AGEMA_signal_12584, new_AGEMA_signal_12583, SubBytesIns_Inst_Sbox_4_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L27_U1 ( .a ({new_AGEMA_signal_10761, new_AGEMA_signal_10760, new_AGEMA_signal_10759, SubBytesIns_Inst_Sbox_4_L8}), .b ({new_AGEMA_signal_11991, new_AGEMA_signal_11990, new_AGEMA_signal_11989, SubBytesIns_Inst_Sbox_4_L10}), .c ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, new_AGEMA_signal_12586, SubBytesIns_Inst_Sbox_4_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L28_U1 ( .a ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, new_AGEMA_signal_11992, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_11421, new_AGEMA_signal_11420, new_AGEMA_signal_11419, SubBytesIns_Inst_Sbox_4_L14}), .c ({new_AGEMA_signal_12591, new_AGEMA_signal_12590, new_AGEMA_signal_12589, SubBytesIns_Inst_Sbox_4_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_L29_U1 ( .a ({new_AGEMA_signal_11994, new_AGEMA_signal_11993, new_AGEMA_signal_11992, SubBytesIns_Inst_Sbox_4_L11}), .b ({new_AGEMA_signal_11427, new_AGEMA_signal_11426, new_AGEMA_signal_11425, SubBytesIns_Inst_Sbox_4_L17}), .c ({new_AGEMA_signal_12594, new_AGEMA_signal_12593, new_AGEMA_signal_12592, SubBytesIns_Inst_Sbox_4_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S0_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_12579, new_AGEMA_signal_12578, new_AGEMA_signal_12577, SubBytesIns_Inst_Sbox_4_L24}), .c ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S1_U1 ( .a ({new_AGEMA_signal_12570, new_AGEMA_signal_12569, new_AGEMA_signal_12568, SubBytesIns_Inst_Sbox_4_L16}), .b ({new_AGEMA_signal_12585, new_AGEMA_signal_12584, new_AGEMA_signal_12583, SubBytesIns_Inst_Sbox_4_L26}), .c ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S2_U1 ( .a ({new_AGEMA_signal_11997, new_AGEMA_signal_11996, new_AGEMA_signal_11995, SubBytesIns_Inst_Sbox_4_L19}), .b ({new_AGEMA_signal_12591, new_AGEMA_signal_12590, new_AGEMA_signal_12589, SubBytesIns_Inst_Sbox_4_L28}), .c ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S3_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_12576, new_AGEMA_signal_12575, new_AGEMA_signal_12574, SubBytesIns_Inst_Sbox_4_L21}), .c ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S4_U1 ( .a ({new_AGEMA_signal_12573, new_AGEMA_signal_12572, new_AGEMA_signal_12571, SubBytesIns_Inst_Sbox_4_L20}), .b ({new_AGEMA_signal_12000, new_AGEMA_signal_11999, new_AGEMA_signal_11998, SubBytesIns_Inst_Sbox_4_L22}), .c ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S5_U1 ( .a ({new_AGEMA_signal_12582, new_AGEMA_signal_12581, new_AGEMA_signal_12580, SubBytesIns_Inst_Sbox_4_L25}), .b ({new_AGEMA_signal_12594, new_AGEMA_signal_12593, new_AGEMA_signal_12592, SubBytesIns_Inst_Sbox_4_L29}), .c ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S6_U1 ( .a ({new_AGEMA_signal_12567, new_AGEMA_signal_12566, new_AGEMA_signal_12565, SubBytesIns_Inst_Sbox_4_L13}), .b ({new_AGEMA_signal_12588, new_AGEMA_signal_12587, new_AGEMA_signal_12586, SubBytesIns_Inst_Sbox_4_L27}), .c ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_4_XOR_S7_U1 ( .a ({new_AGEMA_signal_11982, new_AGEMA_signal_11981, new_AGEMA_signal_11980, SubBytesIns_Inst_Sbox_4_L6}), .b ({new_AGEMA_signal_12003, new_AGEMA_signal_12002, new_AGEMA_signal_12001, SubBytesIns_Inst_Sbox_4_L23}), .c ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M46_U1 ( .a ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_6519, new_AGEMA_signal_6518, new_AGEMA_signal_6517, SubBytesIns_Inst_Sbox_5_T6}), .clk (clk), .r ({Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460]}), .c ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, new_AGEMA_signal_10768, SubBytesIns_Inst_Sbox_5_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M47_U1 ( .a ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_7134, new_AGEMA_signal_7133, new_AGEMA_signal_7132, SubBytesIns_Inst_Sbox_5_T8}), .clk (clk), .r ({Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466]}), .c ({new_AGEMA_signal_10059, new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_5_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M48_U1 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .b ({ciphertext_s3[40], ciphertext_s2[40], ciphertext_s1[40], ciphertext_s0[40]}), .clk (clk), .r ({Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472]}), .c ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, new_AGEMA_signal_10060, SubBytesIns_Inst_Sbox_5_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M49_U1 ( .a ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_6531, new_AGEMA_signal_6530, new_AGEMA_signal_6529, SubBytesIns_Inst_Sbox_5_T16}), .clk (clk), .r ({Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478]}), .c ({new_AGEMA_signal_10773, new_AGEMA_signal_10772, new_AGEMA_signal_10771, SubBytesIns_Inst_Sbox_5_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M50_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_6522, new_AGEMA_signal_6521, new_AGEMA_signal_6520, SubBytesIns_Inst_Sbox_5_T9}), .clk (clk), .r ({Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484]}), .c ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_5_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M51_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_7143, new_AGEMA_signal_7142, new_AGEMA_signal_7141, SubBytesIns_Inst_Sbox_5_T17}), .clk (clk), .r ({Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490]}), .c ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066, SubBytesIns_Inst_Sbox_5_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M52_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_6528, new_AGEMA_signal_6527, new_AGEMA_signal_6526, SubBytesIns_Inst_Sbox_5_T15}), .clk (clk), .r ({Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496]}), .c ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, new_AGEMA_signal_10774, SubBytesIns_Inst_Sbox_5_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M53_U1 ( .a ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, new_AGEMA_signal_10765, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_6540, new_AGEMA_signal_6539, new_AGEMA_signal_6538, SubBytesIns_Inst_Sbox_5_T27}), .clk (clk), .r ({Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502]}), .c ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, new_AGEMA_signal_11431, SubBytesIns_Inst_Sbox_5_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M54_U1 ( .a ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_7137, new_AGEMA_signal_7136, new_AGEMA_signal_7135, SubBytesIns_Inst_Sbox_5_T10}), .clk (clk), .r ({Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508]}), .c ({new_AGEMA_signal_10779, new_AGEMA_signal_10778, new_AGEMA_signal_10777, SubBytesIns_Inst_Sbox_5_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M55_U1 ( .a ({new_AGEMA_signal_10056, new_AGEMA_signal_10055, new_AGEMA_signal_10054, SubBytesIns_Inst_Sbox_5_M44}), .b ({new_AGEMA_signal_6525, new_AGEMA_signal_6524, new_AGEMA_signal_6523, SubBytesIns_Inst_Sbox_5_T13}), .clk (clk), .r ({Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514]}), .c ({new_AGEMA_signal_10782, new_AGEMA_signal_10781, new_AGEMA_signal_10780, SubBytesIns_Inst_Sbox_5_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M56_U1 ( .a ({new_AGEMA_signal_9600, new_AGEMA_signal_9599, new_AGEMA_signal_9598, SubBytesIns_Inst_Sbox_5_M40}), .b ({new_AGEMA_signal_7149, new_AGEMA_signal_7148, new_AGEMA_signal_7147, SubBytesIns_Inst_Sbox_5_T23}), .clk (clk), .r ({Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520]}), .c ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_5_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M57_U1 ( .a ({new_AGEMA_signal_9597, new_AGEMA_signal_9596, new_AGEMA_signal_9595, SubBytesIns_Inst_Sbox_5_M39}), .b ({new_AGEMA_signal_6534, new_AGEMA_signal_6533, new_AGEMA_signal_6532, SubBytesIns_Inst_Sbox_5_T19}), .clk (clk), .r ({Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526]}), .c ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, new_AGEMA_signal_10072, SubBytesIns_Inst_Sbox_5_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M58_U1 ( .a ({new_AGEMA_signal_10053, new_AGEMA_signal_10052, new_AGEMA_signal_10051, SubBytesIns_Inst_Sbox_5_M43}), .b ({new_AGEMA_signal_5979, new_AGEMA_signal_5978, new_AGEMA_signal_5977, SubBytesIns_Inst_Sbox_5_T3}), .clk (clk), .r ({Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532]}), .c ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, new_AGEMA_signal_10783, SubBytesIns_Inst_Sbox_5_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M59_U1 ( .a ({new_AGEMA_signal_9594, new_AGEMA_signal_9593, new_AGEMA_signal_9592, SubBytesIns_Inst_Sbox_5_M38}), .b ({new_AGEMA_signal_6537, new_AGEMA_signal_6536, new_AGEMA_signal_6535, SubBytesIns_Inst_Sbox_5_T22}), .clk (clk), .r ({Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538]}), .c ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_5_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M60_U1 ( .a ({new_AGEMA_signal_9591, new_AGEMA_signal_9590, new_AGEMA_signal_9589, SubBytesIns_Inst_Sbox_5_M37}), .b ({new_AGEMA_signal_7146, new_AGEMA_signal_7145, new_AGEMA_signal_7144, SubBytesIns_Inst_Sbox_5_T20}), .clk (clk), .r ({Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544]}), .c ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, new_AGEMA_signal_10078, SubBytesIns_Inst_Sbox_5_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M61_U1 ( .a ({new_AGEMA_signal_10050, new_AGEMA_signal_10049, new_AGEMA_signal_10048, SubBytesIns_Inst_Sbox_5_M42}), .b ({new_AGEMA_signal_5973, new_AGEMA_signal_5972, new_AGEMA_signal_5971, SubBytesIns_Inst_Sbox_5_T1}), .clk (clk), .r ({Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550]}), .c ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M62_U1 ( .a ({new_AGEMA_signal_10767, new_AGEMA_signal_10766, new_AGEMA_signal_10765, SubBytesIns_Inst_Sbox_5_M45}), .b ({new_AGEMA_signal_5982, new_AGEMA_signal_5981, new_AGEMA_signal_5980, SubBytesIns_Inst_Sbox_5_T4}), .clk (clk), .r ({Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556]}), .c ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, new_AGEMA_signal_11434, SubBytesIns_Inst_Sbox_5_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_AND_M63_U1 ( .a ({new_AGEMA_signal_10047, new_AGEMA_signal_10046, new_AGEMA_signal_10045, SubBytesIns_Inst_Sbox_5_M41}), .b ({new_AGEMA_signal_5976, new_AGEMA_signal_5975, new_AGEMA_signal_5974, SubBytesIns_Inst_Sbox_5_T2}), .clk (clk), .r ({Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562]}), .c ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, new_AGEMA_signal_10789, SubBytesIns_Inst_Sbox_5_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L0_U1 ( .a ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}), .b ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, new_AGEMA_signal_11434, SubBytesIns_Inst_Sbox_5_M62}), .c ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L1_U1 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_5_M56}), .c ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L2_U1 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, new_AGEMA_signal_10768, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, new_AGEMA_signal_10060, SubBytesIns_Inst_Sbox_5_M48}), .c ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, new_AGEMA_signal_11437, SubBytesIns_Inst_Sbox_5_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L3_U1 ( .a ({new_AGEMA_signal_10059, new_AGEMA_signal_10058, new_AGEMA_signal_10057, SubBytesIns_Inst_Sbox_5_M47}), .b ({new_AGEMA_signal_10782, new_AGEMA_signal_10781, new_AGEMA_signal_10780, SubBytesIns_Inst_Sbox_5_M55}), .c ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, new_AGEMA_signal_11440, SubBytesIns_Inst_Sbox_5_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L4_U1 ( .a ({new_AGEMA_signal_10779, new_AGEMA_signal_10778, new_AGEMA_signal_10777, SubBytesIns_Inst_Sbox_5_M54}), .b ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, new_AGEMA_signal_10783, SubBytesIns_Inst_Sbox_5_M58}), .c ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, new_AGEMA_signal_11443, SubBytesIns_Inst_Sbox_5_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L5_U1 ( .a ({new_AGEMA_signal_10773, new_AGEMA_signal_10772, new_AGEMA_signal_10771, SubBytesIns_Inst_Sbox_5_M49}), .b ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, new_AGEMA_signal_11446, SubBytesIns_Inst_Sbox_5_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L6_U1 ( .a ({new_AGEMA_signal_11436, new_AGEMA_signal_11435, new_AGEMA_signal_11434, SubBytesIns_Inst_Sbox_5_M62}), .b ({new_AGEMA_signal_11448, new_AGEMA_signal_11447, new_AGEMA_signal_11446, SubBytesIns_Inst_Sbox_5_L5}), .c ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L7_U1 ( .a ({new_AGEMA_signal_10770, new_AGEMA_signal_10769, new_AGEMA_signal_10768, SubBytesIns_Inst_Sbox_5_M46}), .b ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, new_AGEMA_signal_11440, SubBytesIns_Inst_Sbox_5_L3}), .c ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, new_AGEMA_signal_12010, SubBytesIns_Inst_Sbox_5_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L8_U1 ( .a ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066, SubBytesIns_Inst_Sbox_5_M51}), .b ({new_AGEMA_signal_10077, new_AGEMA_signal_10076, new_AGEMA_signal_10075, SubBytesIns_Inst_Sbox_5_M59}), .c ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, new_AGEMA_signal_10795, SubBytesIns_Inst_Sbox_5_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L9_U1 ( .a ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, new_AGEMA_signal_10774, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, new_AGEMA_signal_11431, SubBytesIns_Inst_Sbox_5_M53}), .c ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, new_AGEMA_signal_12013, SubBytesIns_Inst_Sbox_5_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L10_U1 ( .a ({new_AGEMA_signal_11433, new_AGEMA_signal_11432, new_AGEMA_signal_11431, SubBytesIns_Inst_Sbox_5_M53}), .b ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, new_AGEMA_signal_11443, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, new_AGEMA_signal_12016, SubBytesIns_Inst_Sbox_5_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L11_U1 ( .a ({new_AGEMA_signal_10080, new_AGEMA_signal_10079, new_AGEMA_signal_10078, SubBytesIns_Inst_Sbox_5_M60}), .b ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, new_AGEMA_signal_11437, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, new_AGEMA_signal_12019, SubBytesIns_Inst_Sbox_5_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L12_U1 ( .a ({new_AGEMA_signal_10062, new_AGEMA_signal_10061, new_AGEMA_signal_10060, SubBytesIns_Inst_Sbox_5_M48}), .b ({new_AGEMA_signal_10068, new_AGEMA_signal_10067, new_AGEMA_signal_10066, SubBytesIns_Inst_Sbox_5_M51}), .c ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, new_AGEMA_signal_10798, SubBytesIns_Inst_Sbox_5_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L13_U1 ( .a ({new_AGEMA_signal_10065, new_AGEMA_signal_10064, new_AGEMA_signal_10063, SubBytesIns_Inst_Sbox_5_M50}), .b ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, new_AGEMA_signal_12598, SubBytesIns_Inst_Sbox_5_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L14_U1 ( .a ({new_AGEMA_signal_10776, new_AGEMA_signal_10775, new_AGEMA_signal_10774, SubBytesIns_Inst_Sbox_5_M52}), .b ({new_AGEMA_signal_10788, new_AGEMA_signal_10787, new_AGEMA_signal_10786, SubBytesIns_Inst_Sbox_5_M61}), .c ({new_AGEMA_signal_11451, new_AGEMA_signal_11450, new_AGEMA_signal_11449, SubBytesIns_Inst_Sbox_5_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L15_U1 ( .a ({new_AGEMA_signal_10782, new_AGEMA_signal_10781, new_AGEMA_signal_10780, SubBytesIns_Inst_Sbox_5_M55}), .b ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, new_AGEMA_signal_11452, SubBytesIns_Inst_Sbox_5_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L16_U1 ( .a ({new_AGEMA_signal_10071, new_AGEMA_signal_10070, new_AGEMA_signal_10069, SubBytesIns_Inst_Sbox_5_M56}), .b ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}), .c ({new_AGEMA_signal_12603, new_AGEMA_signal_12602, new_AGEMA_signal_12601, SubBytesIns_Inst_Sbox_5_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L17_U1 ( .a ({new_AGEMA_signal_10074, new_AGEMA_signal_10073, new_AGEMA_signal_10072, SubBytesIns_Inst_Sbox_5_M57}), .b ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_11457, new_AGEMA_signal_11456, new_AGEMA_signal_11455, SubBytesIns_Inst_Sbox_5_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L18_U1 ( .a ({new_AGEMA_signal_10785, new_AGEMA_signal_10784, new_AGEMA_signal_10783, SubBytesIns_Inst_Sbox_5_M58}), .b ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, new_AGEMA_signal_10795, SubBytesIns_Inst_Sbox_5_L8}), .c ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, new_AGEMA_signal_11458, SubBytesIns_Inst_Sbox_5_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L19_U1 ( .a ({new_AGEMA_signal_10791, new_AGEMA_signal_10790, new_AGEMA_signal_10789, SubBytesIns_Inst_Sbox_5_M63}), .b ({new_AGEMA_signal_11445, new_AGEMA_signal_11444, new_AGEMA_signal_11443, SubBytesIns_Inst_Sbox_5_L4}), .c ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, new_AGEMA_signal_12022, SubBytesIns_Inst_Sbox_5_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L20_U1 ( .a ({new_AGEMA_signal_12006, new_AGEMA_signal_12005, new_AGEMA_signal_12004, SubBytesIns_Inst_Sbox_5_L0}), .b ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .c ({new_AGEMA_signal_12606, new_AGEMA_signal_12605, new_AGEMA_signal_12604, SubBytesIns_Inst_Sbox_5_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L21_U1 ( .a ({new_AGEMA_signal_10794, new_AGEMA_signal_10793, new_AGEMA_signal_10792, SubBytesIns_Inst_Sbox_5_L1}), .b ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, new_AGEMA_signal_12010, SubBytesIns_Inst_Sbox_5_L7}), .c ({new_AGEMA_signal_12609, new_AGEMA_signal_12608, new_AGEMA_signal_12607, SubBytesIns_Inst_Sbox_5_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L22_U1 ( .a ({new_AGEMA_signal_11442, new_AGEMA_signal_11441, new_AGEMA_signal_11440, SubBytesIns_Inst_Sbox_5_L3}), .b ({new_AGEMA_signal_10800, new_AGEMA_signal_10799, new_AGEMA_signal_10798, SubBytesIns_Inst_Sbox_5_L12}), .c ({new_AGEMA_signal_12027, new_AGEMA_signal_12026, new_AGEMA_signal_12025, SubBytesIns_Inst_Sbox_5_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L23_U1 ( .a ({new_AGEMA_signal_11460, new_AGEMA_signal_11459, new_AGEMA_signal_11458, SubBytesIns_Inst_Sbox_5_L18}), .b ({new_AGEMA_signal_11439, new_AGEMA_signal_11438, new_AGEMA_signal_11437, SubBytesIns_Inst_Sbox_5_L2}), .c ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, new_AGEMA_signal_12028, SubBytesIns_Inst_Sbox_5_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L24_U1 ( .a ({new_AGEMA_signal_11454, new_AGEMA_signal_11453, new_AGEMA_signal_11452, SubBytesIns_Inst_Sbox_5_L15}), .b ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, new_AGEMA_signal_12013, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, new_AGEMA_signal_12610, SubBytesIns_Inst_Sbox_5_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L25_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, new_AGEMA_signal_12016, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_12615, new_AGEMA_signal_12614, new_AGEMA_signal_12613, SubBytesIns_Inst_Sbox_5_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L26_U1 ( .a ({new_AGEMA_signal_12012, new_AGEMA_signal_12011, new_AGEMA_signal_12010, SubBytesIns_Inst_Sbox_5_L7}), .b ({new_AGEMA_signal_12015, new_AGEMA_signal_12014, new_AGEMA_signal_12013, SubBytesIns_Inst_Sbox_5_L9}), .c ({new_AGEMA_signal_12618, new_AGEMA_signal_12617, new_AGEMA_signal_12616, SubBytesIns_Inst_Sbox_5_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L27_U1 ( .a ({new_AGEMA_signal_10797, new_AGEMA_signal_10796, new_AGEMA_signal_10795, SubBytesIns_Inst_Sbox_5_L8}), .b ({new_AGEMA_signal_12018, new_AGEMA_signal_12017, new_AGEMA_signal_12016, SubBytesIns_Inst_Sbox_5_L10}), .c ({new_AGEMA_signal_12621, new_AGEMA_signal_12620, new_AGEMA_signal_12619, SubBytesIns_Inst_Sbox_5_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L28_U1 ( .a ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, new_AGEMA_signal_12019, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_11451, new_AGEMA_signal_11450, new_AGEMA_signal_11449, SubBytesIns_Inst_Sbox_5_L14}), .c ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, new_AGEMA_signal_12622, SubBytesIns_Inst_Sbox_5_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_L29_U1 ( .a ({new_AGEMA_signal_12021, new_AGEMA_signal_12020, new_AGEMA_signal_12019, SubBytesIns_Inst_Sbox_5_L11}), .b ({new_AGEMA_signal_11457, new_AGEMA_signal_11456, new_AGEMA_signal_11455, SubBytesIns_Inst_Sbox_5_L17}), .c ({new_AGEMA_signal_12627, new_AGEMA_signal_12626, new_AGEMA_signal_12625, SubBytesIns_Inst_Sbox_5_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S0_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12612, new_AGEMA_signal_12611, new_AGEMA_signal_12610, SubBytesIns_Inst_Sbox_5_L24}), .c ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S1_U1 ( .a ({new_AGEMA_signal_12603, new_AGEMA_signal_12602, new_AGEMA_signal_12601, SubBytesIns_Inst_Sbox_5_L16}), .b ({new_AGEMA_signal_12618, new_AGEMA_signal_12617, new_AGEMA_signal_12616, SubBytesIns_Inst_Sbox_5_L26}), .c ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S2_U1 ( .a ({new_AGEMA_signal_12024, new_AGEMA_signal_12023, new_AGEMA_signal_12022, SubBytesIns_Inst_Sbox_5_L19}), .b ({new_AGEMA_signal_12624, new_AGEMA_signal_12623, new_AGEMA_signal_12622, SubBytesIns_Inst_Sbox_5_L28}), .c ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S3_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12609, new_AGEMA_signal_12608, new_AGEMA_signal_12607, SubBytesIns_Inst_Sbox_5_L21}), .c ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S4_U1 ( .a ({new_AGEMA_signal_12606, new_AGEMA_signal_12605, new_AGEMA_signal_12604, SubBytesIns_Inst_Sbox_5_L20}), .b ({new_AGEMA_signal_12027, new_AGEMA_signal_12026, new_AGEMA_signal_12025, SubBytesIns_Inst_Sbox_5_L22}), .c ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S5_U1 ( .a ({new_AGEMA_signal_12615, new_AGEMA_signal_12614, new_AGEMA_signal_12613, SubBytesIns_Inst_Sbox_5_L25}), .b ({new_AGEMA_signal_12627, new_AGEMA_signal_12626, new_AGEMA_signal_12625, SubBytesIns_Inst_Sbox_5_L29}), .c ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S6_U1 ( .a ({new_AGEMA_signal_12600, new_AGEMA_signal_12599, new_AGEMA_signal_12598, SubBytesIns_Inst_Sbox_5_L13}), .b ({new_AGEMA_signal_12621, new_AGEMA_signal_12620, new_AGEMA_signal_12619, SubBytesIns_Inst_Sbox_5_L27}), .c ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_5_XOR_S7_U1 ( .a ({new_AGEMA_signal_12009, new_AGEMA_signal_12008, new_AGEMA_signal_12007, SubBytesIns_Inst_Sbox_5_L6}), .b ({new_AGEMA_signal_12030, new_AGEMA_signal_12029, new_AGEMA_signal_12028, SubBytesIns_Inst_Sbox_5_L23}), .c ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M46_U1 ( .a ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, new_AGEMA_signal_10090, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_6543, new_AGEMA_signal_6542, new_AGEMA_signal_6541, SubBytesIns_Inst_Sbox_6_T6}), .clk (clk), .r ({Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568]}), .c ({new_AGEMA_signal_10806, new_AGEMA_signal_10805, new_AGEMA_signal_10804, SubBytesIns_Inst_Sbox_6_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M47_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_7173, new_AGEMA_signal_7172, new_AGEMA_signal_7171, SubBytesIns_Inst_Sbox_6_T8}), .clk (clk), .r ({Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574]}), .c ({new_AGEMA_signal_10095, new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_6_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M48_U1 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .b ({ciphertext_s3[48], ciphertext_s2[48], ciphertext_s1[48], ciphertext_s0[48]}), .clk (clk), .r ({Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580]}), .c ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, new_AGEMA_signal_10096, SubBytesIns_Inst_Sbox_6_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M49_U1 ( .a ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_6555, new_AGEMA_signal_6554, new_AGEMA_signal_6553, SubBytesIns_Inst_Sbox_6_T16}), .clk (clk), .r ({Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586]}), .c ({new_AGEMA_signal_10809, new_AGEMA_signal_10808, new_AGEMA_signal_10807, SubBytesIns_Inst_Sbox_6_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M50_U1 ( .a ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_6546, new_AGEMA_signal_6545, new_AGEMA_signal_6544, SubBytesIns_Inst_Sbox_6_T9}), .clk (clk), .r ({Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592]}), .c ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_6_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M51_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_7182, new_AGEMA_signal_7181, new_AGEMA_signal_7180, SubBytesIns_Inst_Sbox_6_T17}), .clk (clk), .r ({Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598]}), .c ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, new_AGEMA_signal_10102, SubBytesIns_Inst_Sbox_6_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M52_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_6552, new_AGEMA_signal_6551, new_AGEMA_signal_6550, SubBytesIns_Inst_Sbox_6_T15}), .clk (clk), .r ({Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604]}), .c ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, new_AGEMA_signal_10810, SubBytesIns_Inst_Sbox_6_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M53_U1 ( .a ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, new_AGEMA_signal_10801, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_6564, new_AGEMA_signal_6563, new_AGEMA_signal_6562, SubBytesIns_Inst_Sbox_6_T27}), .clk (clk), .r ({Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610]}), .c ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, new_AGEMA_signal_11461, SubBytesIns_Inst_Sbox_6_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M54_U1 ( .a ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_7176, new_AGEMA_signal_7175, new_AGEMA_signal_7174, SubBytesIns_Inst_Sbox_6_T10}), .clk (clk), .r ({Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616]}), .c ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, new_AGEMA_signal_10813, SubBytesIns_Inst_Sbox_6_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M55_U1 ( .a ({new_AGEMA_signal_10092, new_AGEMA_signal_10091, new_AGEMA_signal_10090, SubBytesIns_Inst_Sbox_6_M44}), .b ({new_AGEMA_signal_6549, new_AGEMA_signal_6548, new_AGEMA_signal_6547, SubBytesIns_Inst_Sbox_6_T13}), .clk (clk), .r ({Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622]}), .c ({new_AGEMA_signal_10818, new_AGEMA_signal_10817, new_AGEMA_signal_10816, SubBytesIns_Inst_Sbox_6_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M56_U1 ( .a ({new_AGEMA_signal_9612, new_AGEMA_signal_9611, new_AGEMA_signal_9610, SubBytesIns_Inst_Sbox_6_M40}), .b ({new_AGEMA_signal_7188, new_AGEMA_signal_7187, new_AGEMA_signal_7186, SubBytesIns_Inst_Sbox_6_T23}), .clk (clk), .r ({Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628]}), .c ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_6_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M57_U1 ( .a ({new_AGEMA_signal_9609, new_AGEMA_signal_9608, new_AGEMA_signal_9607, SubBytesIns_Inst_Sbox_6_M39}), .b ({new_AGEMA_signal_6558, new_AGEMA_signal_6557, new_AGEMA_signal_6556, SubBytesIns_Inst_Sbox_6_T19}), .clk (clk), .r ({Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634]}), .c ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, new_AGEMA_signal_10108, SubBytesIns_Inst_Sbox_6_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M58_U1 ( .a ({new_AGEMA_signal_10089, new_AGEMA_signal_10088, new_AGEMA_signal_10087, SubBytesIns_Inst_Sbox_6_M43}), .b ({new_AGEMA_signal_6009, new_AGEMA_signal_6008, new_AGEMA_signal_6007, SubBytesIns_Inst_Sbox_6_T3}), .clk (clk), .r ({Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640]}), .c ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, new_AGEMA_signal_10819, SubBytesIns_Inst_Sbox_6_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M59_U1 ( .a ({new_AGEMA_signal_9606, new_AGEMA_signal_9605, new_AGEMA_signal_9604, SubBytesIns_Inst_Sbox_6_M38}), .b ({new_AGEMA_signal_6561, new_AGEMA_signal_6560, new_AGEMA_signal_6559, SubBytesIns_Inst_Sbox_6_T22}), .clk (clk), .r ({Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646]}), .c ({new_AGEMA_signal_10113, new_AGEMA_signal_10112, new_AGEMA_signal_10111, SubBytesIns_Inst_Sbox_6_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M60_U1 ( .a ({new_AGEMA_signal_9603, new_AGEMA_signal_9602, new_AGEMA_signal_9601, SubBytesIns_Inst_Sbox_6_M37}), .b ({new_AGEMA_signal_7185, new_AGEMA_signal_7184, new_AGEMA_signal_7183, SubBytesIns_Inst_Sbox_6_T20}), .clk (clk), .r ({Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652]}), .c ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, new_AGEMA_signal_10114, SubBytesIns_Inst_Sbox_6_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M61_U1 ( .a ({new_AGEMA_signal_10086, new_AGEMA_signal_10085, new_AGEMA_signal_10084, SubBytesIns_Inst_Sbox_6_M42}), .b ({new_AGEMA_signal_6003, new_AGEMA_signal_6002, new_AGEMA_signal_6001, SubBytesIns_Inst_Sbox_6_T1}), .clk (clk), .r ({Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658]}), .c ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M62_U1 ( .a ({new_AGEMA_signal_10803, new_AGEMA_signal_10802, new_AGEMA_signal_10801, SubBytesIns_Inst_Sbox_6_M45}), .b ({new_AGEMA_signal_6012, new_AGEMA_signal_6011, new_AGEMA_signal_6010, SubBytesIns_Inst_Sbox_6_T4}), .clk (clk), .r ({Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664]}), .c ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, new_AGEMA_signal_11464, SubBytesIns_Inst_Sbox_6_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_AND_M63_U1 ( .a ({new_AGEMA_signal_10083, new_AGEMA_signal_10082, new_AGEMA_signal_10081, SubBytesIns_Inst_Sbox_6_M41}), .b ({new_AGEMA_signal_6006, new_AGEMA_signal_6005, new_AGEMA_signal_6004, SubBytesIns_Inst_Sbox_6_T2}), .clk (clk), .r ({Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670]}), .c ({new_AGEMA_signal_10827, new_AGEMA_signal_10826, new_AGEMA_signal_10825, SubBytesIns_Inst_Sbox_6_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L0_U1 ( .a ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}), .b ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, new_AGEMA_signal_11464, SubBytesIns_Inst_Sbox_6_M62}), .c ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L1_U1 ( .a ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_6_M56}), .c ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L2_U1 ( .a ({new_AGEMA_signal_10806, new_AGEMA_signal_10805, new_AGEMA_signal_10804, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, new_AGEMA_signal_10096, SubBytesIns_Inst_Sbox_6_M48}), .c ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, new_AGEMA_signal_11467, SubBytesIns_Inst_Sbox_6_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L3_U1 ( .a ({new_AGEMA_signal_10095, new_AGEMA_signal_10094, new_AGEMA_signal_10093, SubBytesIns_Inst_Sbox_6_M47}), .b ({new_AGEMA_signal_10818, new_AGEMA_signal_10817, new_AGEMA_signal_10816, SubBytesIns_Inst_Sbox_6_M55}), .c ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, new_AGEMA_signal_11470, SubBytesIns_Inst_Sbox_6_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L4_U1 ( .a ({new_AGEMA_signal_10815, new_AGEMA_signal_10814, new_AGEMA_signal_10813, SubBytesIns_Inst_Sbox_6_M54}), .b ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, new_AGEMA_signal_10819, SubBytesIns_Inst_Sbox_6_M58}), .c ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, new_AGEMA_signal_11473, SubBytesIns_Inst_Sbox_6_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L5_U1 ( .a ({new_AGEMA_signal_10809, new_AGEMA_signal_10808, new_AGEMA_signal_10807, SubBytesIns_Inst_Sbox_6_M49}), .b ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, new_AGEMA_signal_11476, SubBytesIns_Inst_Sbox_6_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L6_U1 ( .a ({new_AGEMA_signal_11466, new_AGEMA_signal_11465, new_AGEMA_signal_11464, SubBytesIns_Inst_Sbox_6_M62}), .b ({new_AGEMA_signal_11478, new_AGEMA_signal_11477, new_AGEMA_signal_11476, SubBytesIns_Inst_Sbox_6_L5}), .c ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L7_U1 ( .a ({new_AGEMA_signal_10806, new_AGEMA_signal_10805, new_AGEMA_signal_10804, SubBytesIns_Inst_Sbox_6_M46}), .b ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, new_AGEMA_signal_11470, SubBytesIns_Inst_Sbox_6_L3}), .c ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, new_AGEMA_signal_12037, SubBytesIns_Inst_Sbox_6_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L8_U1 ( .a ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, new_AGEMA_signal_10102, SubBytesIns_Inst_Sbox_6_M51}), .b ({new_AGEMA_signal_10113, new_AGEMA_signal_10112, new_AGEMA_signal_10111, SubBytesIns_Inst_Sbox_6_M59}), .c ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, new_AGEMA_signal_10831, SubBytesIns_Inst_Sbox_6_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L9_U1 ( .a ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, new_AGEMA_signal_10810, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, new_AGEMA_signal_11461, SubBytesIns_Inst_Sbox_6_M53}), .c ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, new_AGEMA_signal_12040, SubBytesIns_Inst_Sbox_6_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L10_U1 ( .a ({new_AGEMA_signal_11463, new_AGEMA_signal_11462, new_AGEMA_signal_11461, SubBytesIns_Inst_Sbox_6_M53}), .b ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, new_AGEMA_signal_11473, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, new_AGEMA_signal_12043, SubBytesIns_Inst_Sbox_6_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L11_U1 ( .a ({new_AGEMA_signal_10116, new_AGEMA_signal_10115, new_AGEMA_signal_10114, SubBytesIns_Inst_Sbox_6_M60}), .b ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, new_AGEMA_signal_11467, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, new_AGEMA_signal_12046, SubBytesIns_Inst_Sbox_6_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L12_U1 ( .a ({new_AGEMA_signal_10098, new_AGEMA_signal_10097, new_AGEMA_signal_10096, SubBytesIns_Inst_Sbox_6_M48}), .b ({new_AGEMA_signal_10104, new_AGEMA_signal_10103, new_AGEMA_signal_10102, SubBytesIns_Inst_Sbox_6_M51}), .c ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, new_AGEMA_signal_10834, SubBytesIns_Inst_Sbox_6_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L13_U1 ( .a ({new_AGEMA_signal_10101, new_AGEMA_signal_10100, new_AGEMA_signal_10099, SubBytesIns_Inst_Sbox_6_M50}), .b ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_12633, new_AGEMA_signal_12632, new_AGEMA_signal_12631, SubBytesIns_Inst_Sbox_6_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L14_U1 ( .a ({new_AGEMA_signal_10812, new_AGEMA_signal_10811, new_AGEMA_signal_10810, SubBytesIns_Inst_Sbox_6_M52}), .b ({new_AGEMA_signal_10824, new_AGEMA_signal_10823, new_AGEMA_signal_10822, SubBytesIns_Inst_Sbox_6_M61}), .c ({new_AGEMA_signal_11481, new_AGEMA_signal_11480, new_AGEMA_signal_11479, SubBytesIns_Inst_Sbox_6_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L15_U1 ( .a ({new_AGEMA_signal_10818, new_AGEMA_signal_10817, new_AGEMA_signal_10816, SubBytesIns_Inst_Sbox_6_M55}), .b ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, new_AGEMA_signal_11482, SubBytesIns_Inst_Sbox_6_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L16_U1 ( .a ({new_AGEMA_signal_10107, new_AGEMA_signal_10106, new_AGEMA_signal_10105, SubBytesIns_Inst_Sbox_6_M56}), .b ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}), .c ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, new_AGEMA_signal_12634, SubBytesIns_Inst_Sbox_6_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L17_U1 ( .a ({new_AGEMA_signal_10110, new_AGEMA_signal_10109, new_AGEMA_signal_10108, SubBytesIns_Inst_Sbox_6_M57}), .b ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_11487, new_AGEMA_signal_11486, new_AGEMA_signal_11485, SubBytesIns_Inst_Sbox_6_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L18_U1 ( .a ({new_AGEMA_signal_10821, new_AGEMA_signal_10820, new_AGEMA_signal_10819, SubBytesIns_Inst_Sbox_6_M58}), .b ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, new_AGEMA_signal_10831, SubBytesIns_Inst_Sbox_6_L8}), .c ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, new_AGEMA_signal_11488, SubBytesIns_Inst_Sbox_6_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L19_U1 ( .a ({new_AGEMA_signal_10827, new_AGEMA_signal_10826, new_AGEMA_signal_10825, SubBytesIns_Inst_Sbox_6_M63}), .b ({new_AGEMA_signal_11475, new_AGEMA_signal_11474, new_AGEMA_signal_11473, SubBytesIns_Inst_Sbox_6_L4}), .c ({new_AGEMA_signal_12051, new_AGEMA_signal_12050, new_AGEMA_signal_12049, SubBytesIns_Inst_Sbox_6_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L20_U1 ( .a ({new_AGEMA_signal_12033, new_AGEMA_signal_12032, new_AGEMA_signal_12031, SubBytesIns_Inst_Sbox_6_L0}), .b ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .c ({new_AGEMA_signal_12639, new_AGEMA_signal_12638, new_AGEMA_signal_12637, SubBytesIns_Inst_Sbox_6_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L21_U1 ( .a ({new_AGEMA_signal_10830, new_AGEMA_signal_10829, new_AGEMA_signal_10828, SubBytesIns_Inst_Sbox_6_L1}), .b ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, new_AGEMA_signal_12037, SubBytesIns_Inst_Sbox_6_L7}), .c ({new_AGEMA_signal_12642, new_AGEMA_signal_12641, new_AGEMA_signal_12640, SubBytesIns_Inst_Sbox_6_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L22_U1 ( .a ({new_AGEMA_signal_11472, new_AGEMA_signal_11471, new_AGEMA_signal_11470, SubBytesIns_Inst_Sbox_6_L3}), .b ({new_AGEMA_signal_10836, new_AGEMA_signal_10835, new_AGEMA_signal_10834, SubBytesIns_Inst_Sbox_6_L12}), .c ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, new_AGEMA_signal_12052, SubBytesIns_Inst_Sbox_6_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L23_U1 ( .a ({new_AGEMA_signal_11490, new_AGEMA_signal_11489, new_AGEMA_signal_11488, SubBytesIns_Inst_Sbox_6_L18}), .b ({new_AGEMA_signal_11469, new_AGEMA_signal_11468, new_AGEMA_signal_11467, SubBytesIns_Inst_Sbox_6_L2}), .c ({new_AGEMA_signal_12057, new_AGEMA_signal_12056, new_AGEMA_signal_12055, SubBytesIns_Inst_Sbox_6_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L24_U1 ( .a ({new_AGEMA_signal_11484, new_AGEMA_signal_11483, new_AGEMA_signal_11482, SubBytesIns_Inst_Sbox_6_L15}), .b ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, new_AGEMA_signal_12040, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_12645, new_AGEMA_signal_12644, new_AGEMA_signal_12643, SubBytesIns_Inst_Sbox_6_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L25_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, new_AGEMA_signal_12043, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, new_AGEMA_signal_12646, SubBytesIns_Inst_Sbox_6_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L26_U1 ( .a ({new_AGEMA_signal_12039, new_AGEMA_signal_12038, new_AGEMA_signal_12037, SubBytesIns_Inst_Sbox_6_L7}), .b ({new_AGEMA_signal_12042, new_AGEMA_signal_12041, new_AGEMA_signal_12040, SubBytesIns_Inst_Sbox_6_L9}), .c ({new_AGEMA_signal_12651, new_AGEMA_signal_12650, new_AGEMA_signal_12649, SubBytesIns_Inst_Sbox_6_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L27_U1 ( .a ({new_AGEMA_signal_10833, new_AGEMA_signal_10832, new_AGEMA_signal_10831, SubBytesIns_Inst_Sbox_6_L8}), .b ({new_AGEMA_signal_12045, new_AGEMA_signal_12044, new_AGEMA_signal_12043, SubBytesIns_Inst_Sbox_6_L10}), .c ({new_AGEMA_signal_12654, new_AGEMA_signal_12653, new_AGEMA_signal_12652, SubBytesIns_Inst_Sbox_6_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L28_U1 ( .a ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, new_AGEMA_signal_12046, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_11481, new_AGEMA_signal_11480, new_AGEMA_signal_11479, SubBytesIns_Inst_Sbox_6_L14}), .c ({new_AGEMA_signal_12657, new_AGEMA_signal_12656, new_AGEMA_signal_12655, SubBytesIns_Inst_Sbox_6_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_L29_U1 ( .a ({new_AGEMA_signal_12048, new_AGEMA_signal_12047, new_AGEMA_signal_12046, SubBytesIns_Inst_Sbox_6_L11}), .b ({new_AGEMA_signal_11487, new_AGEMA_signal_11486, new_AGEMA_signal_11485, SubBytesIns_Inst_Sbox_6_L17}), .c ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, new_AGEMA_signal_12658, SubBytesIns_Inst_Sbox_6_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S0_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12645, new_AGEMA_signal_12644, new_AGEMA_signal_12643, SubBytesIns_Inst_Sbox_6_L24}), .c ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S1_U1 ( .a ({new_AGEMA_signal_12636, new_AGEMA_signal_12635, new_AGEMA_signal_12634, SubBytesIns_Inst_Sbox_6_L16}), .b ({new_AGEMA_signal_12651, new_AGEMA_signal_12650, new_AGEMA_signal_12649, SubBytesIns_Inst_Sbox_6_L26}), .c ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S2_U1 ( .a ({new_AGEMA_signal_12051, new_AGEMA_signal_12050, new_AGEMA_signal_12049, SubBytesIns_Inst_Sbox_6_L19}), .b ({new_AGEMA_signal_12657, new_AGEMA_signal_12656, new_AGEMA_signal_12655, SubBytesIns_Inst_Sbox_6_L28}), .c ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S3_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12642, new_AGEMA_signal_12641, new_AGEMA_signal_12640, SubBytesIns_Inst_Sbox_6_L21}), .c ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S4_U1 ( .a ({new_AGEMA_signal_12639, new_AGEMA_signal_12638, new_AGEMA_signal_12637, SubBytesIns_Inst_Sbox_6_L20}), .b ({new_AGEMA_signal_12054, new_AGEMA_signal_12053, new_AGEMA_signal_12052, SubBytesIns_Inst_Sbox_6_L22}), .c ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S5_U1 ( .a ({new_AGEMA_signal_12648, new_AGEMA_signal_12647, new_AGEMA_signal_12646, SubBytesIns_Inst_Sbox_6_L25}), .b ({new_AGEMA_signal_12660, new_AGEMA_signal_12659, new_AGEMA_signal_12658, SubBytesIns_Inst_Sbox_6_L29}), .c ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S6_U1 ( .a ({new_AGEMA_signal_12633, new_AGEMA_signal_12632, new_AGEMA_signal_12631, SubBytesIns_Inst_Sbox_6_L13}), .b ({new_AGEMA_signal_12654, new_AGEMA_signal_12653, new_AGEMA_signal_12652, SubBytesIns_Inst_Sbox_6_L27}), .c ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_6_XOR_S7_U1 ( .a ({new_AGEMA_signal_12036, new_AGEMA_signal_12035, new_AGEMA_signal_12034, SubBytesIns_Inst_Sbox_6_L6}), .b ({new_AGEMA_signal_12057, new_AGEMA_signal_12056, new_AGEMA_signal_12055, SubBytesIns_Inst_Sbox_6_L23}), .c ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M46_U1 ( .a ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, new_AGEMA_signal_10126, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_6567, new_AGEMA_signal_6566, new_AGEMA_signal_6565, SubBytesIns_Inst_Sbox_7_T6}), .clk (clk), .r ({Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676]}), .c ({new_AGEMA_signal_10842, new_AGEMA_signal_10841, new_AGEMA_signal_10840, SubBytesIns_Inst_Sbox_7_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M47_U1 ( .a ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_7212, new_AGEMA_signal_7211, new_AGEMA_signal_7210, SubBytesIns_Inst_Sbox_7_T8}), .clk (clk), .r ({Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682]}), .c ({new_AGEMA_signal_10131, new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_7_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M48_U1 ( .a ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .b ({ciphertext_s3[56], ciphertext_s2[56], ciphertext_s1[56], ciphertext_s0[56]}), .clk (clk), .r ({Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688]}), .c ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, new_AGEMA_signal_10132, SubBytesIns_Inst_Sbox_7_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M49_U1 ( .a ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_6579, new_AGEMA_signal_6578, new_AGEMA_signal_6577, SubBytesIns_Inst_Sbox_7_T16}), .clk (clk), .r ({Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694]}), .c ({new_AGEMA_signal_10845, new_AGEMA_signal_10844, new_AGEMA_signal_10843, SubBytesIns_Inst_Sbox_7_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M50_U1 ( .a ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_6570, new_AGEMA_signal_6569, new_AGEMA_signal_6568, SubBytesIns_Inst_Sbox_7_T9}), .clk (clk), .r ({Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700]}), .c ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_7_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M51_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_7221, new_AGEMA_signal_7220, new_AGEMA_signal_7219, SubBytesIns_Inst_Sbox_7_T17}), .clk (clk), .r ({Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706]}), .c ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, new_AGEMA_signal_10138, SubBytesIns_Inst_Sbox_7_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M52_U1 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_6576, new_AGEMA_signal_6575, new_AGEMA_signal_6574, SubBytesIns_Inst_Sbox_7_T15}), .clk (clk), .r ({Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712]}), .c ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, new_AGEMA_signal_10846, SubBytesIns_Inst_Sbox_7_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M53_U1 ( .a ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, new_AGEMA_signal_10837, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_6588, new_AGEMA_signal_6587, new_AGEMA_signal_6586, SubBytesIns_Inst_Sbox_7_T27}), .clk (clk), .r ({Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718]}), .c ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, new_AGEMA_signal_11491, SubBytesIns_Inst_Sbox_7_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M54_U1 ( .a ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_7215, new_AGEMA_signal_7214, new_AGEMA_signal_7213, SubBytesIns_Inst_Sbox_7_T10}), .clk (clk), .r ({Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724]}), .c ({new_AGEMA_signal_10851, new_AGEMA_signal_10850, new_AGEMA_signal_10849, SubBytesIns_Inst_Sbox_7_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M55_U1 ( .a ({new_AGEMA_signal_10128, new_AGEMA_signal_10127, new_AGEMA_signal_10126, SubBytesIns_Inst_Sbox_7_M44}), .b ({new_AGEMA_signal_6573, new_AGEMA_signal_6572, new_AGEMA_signal_6571, SubBytesIns_Inst_Sbox_7_T13}), .clk (clk), .r ({Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730]}), .c ({new_AGEMA_signal_10854, new_AGEMA_signal_10853, new_AGEMA_signal_10852, SubBytesIns_Inst_Sbox_7_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M56_U1 ( .a ({new_AGEMA_signal_9624, new_AGEMA_signal_9623, new_AGEMA_signal_9622, SubBytesIns_Inst_Sbox_7_M40}), .b ({new_AGEMA_signal_7227, new_AGEMA_signal_7226, new_AGEMA_signal_7225, SubBytesIns_Inst_Sbox_7_T23}), .clk (clk), .r ({Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736]}), .c ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_7_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M57_U1 ( .a ({new_AGEMA_signal_9621, new_AGEMA_signal_9620, new_AGEMA_signal_9619, SubBytesIns_Inst_Sbox_7_M39}), .b ({new_AGEMA_signal_6582, new_AGEMA_signal_6581, new_AGEMA_signal_6580, SubBytesIns_Inst_Sbox_7_T19}), .clk (clk), .r ({Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742]}), .c ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, new_AGEMA_signal_10144, SubBytesIns_Inst_Sbox_7_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M58_U1 ( .a ({new_AGEMA_signal_10125, new_AGEMA_signal_10124, new_AGEMA_signal_10123, SubBytesIns_Inst_Sbox_7_M43}), .b ({new_AGEMA_signal_6039, new_AGEMA_signal_6038, new_AGEMA_signal_6037, SubBytesIns_Inst_Sbox_7_T3}), .clk (clk), .r ({Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748]}), .c ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, new_AGEMA_signal_10855, SubBytesIns_Inst_Sbox_7_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M59_U1 ( .a ({new_AGEMA_signal_9618, new_AGEMA_signal_9617, new_AGEMA_signal_9616, SubBytesIns_Inst_Sbox_7_M38}), .b ({new_AGEMA_signal_6585, new_AGEMA_signal_6584, new_AGEMA_signal_6583, SubBytesIns_Inst_Sbox_7_T22}), .clk (clk), .r ({Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754]}), .c ({new_AGEMA_signal_10149, new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_7_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M60_U1 ( .a ({new_AGEMA_signal_9615, new_AGEMA_signal_9614, new_AGEMA_signal_9613, SubBytesIns_Inst_Sbox_7_M37}), .b ({new_AGEMA_signal_7224, new_AGEMA_signal_7223, new_AGEMA_signal_7222, SubBytesIns_Inst_Sbox_7_T20}), .clk (clk), .r ({Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760]}), .c ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, new_AGEMA_signal_10150, SubBytesIns_Inst_Sbox_7_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M61_U1 ( .a ({new_AGEMA_signal_10122, new_AGEMA_signal_10121, new_AGEMA_signal_10120, SubBytesIns_Inst_Sbox_7_M42}), .b ({new_AGEMA_signal_6033, new_AGEMA_signal_6032, new_AGEMA_signal_6031, SubBytesIns_Inst_Sbox_7_T1}), .clk (clk), .r ({Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766]}), .c ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M62_U1 ( .a ({new_AGEMA_signal_10839, new_AGEMA_signal_10838, new_AGEMA_signal_10837, SubBytesIns_Inst_Sbox_7_M45}), .b ({new_AGEMA_signal_6042, new_AGEMA_signal_6041, new_AGEMA_signal_6040, SubBytesIns_Inst_Sbox_7_T4}), .clk (clk), .r ({Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772]}), .c ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, new_AGEMA_signal_11494, SubBytesIns_Inst_Sbox_7_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_AND_M63_U1 ( .a ({new_AGEMA_signal_10119, new_AGEMA_signal_10118, new_AGEMA_signal_10117, SubBytesIns_Inst_Sbox_7_M41}), .b ({new_AGEMA_signal_6036, new_AGEMA_signal_6035, new_AGEMA_signal_6034, SubBytesIns_Inst_Sbox_7_T2}), .clk (clk), .r ({Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778]}), .c ({new_AGEMA_signal_10863, new_AGEMA_signal_10862, new_AGEMA_signal_10861, SubBytesIns_Inst_Sbox_7_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L0_U1 ( .a ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}), .b ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, new_AGEMA_signal_11494, SubBytesIns_Inst_Sbox_7_M62}), .c ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L1_U1 ( .a ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_7_M56}), .c ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L2_U1 ( .a ({new_AGEMA_signal_10842, new_AGEMA_signal_10841, new_AGEMA_signal_10840, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, new_AGEMA_signal_10132, SubBytesIns_Inst_Sbox_7_M48}), .c ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, new_AGEMA_signal_11497, SubBytesIns_Inst_Sbox_7_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L3_U1 ( .a ({new_AGEMA_signal_10131, new_AGEMA_signal_10130, new_AGEMA_signal_10129, SubBytesIns_Inst_Sbox_7_M47}), .b ({new_AGEMA_signal_10854, new_AGEMA_signal_10853, new_AGEMA_signal_10852, SubBytesIns_Inst_Sbox_7_M55}), .c ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, new_AGEMA_signal_11500, SubBytesIns_Inst_Sbox_7_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L4_U1 ( .a ({new_AGEMA_signal_10851, new_AGEMA_signal_10850, new_AGEMA_signal_10849, SubBytesIns_Inst_Sbox_7_M54}), .b ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, new_AGEMA_signal_10855, SubBytesIns_Inst_Sbox_7_M58}), .c ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, new_AGEMA_signal_11503, SubBytesIns_Inst_Sbox_7_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L5_U1 ( .a ({new_AGEMA_signal_10845, new_AGEMA_signal_10844, new_AGEMA_signal_10843, SubBytesIns_Inst_Sbox_7_M49}), .b ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, new_AGEMA_signal_11506, SubBytesIns_Inst_Sbox_7_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L6_U1 ( .a ({new_AGEMA_signal_11496, new_AGEMA_signal_11495, new_AGEMA_signal_11494, SubBytesIns_Inst_Sbox_7_M62}), .b ({new_AGEMA_signal_11508, new_AGEMA_signal_11507, new_AGEMA_signal_11506, SubBytesIns_Inst_Sbox_7_L5}), .c ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L7_U1 ( .a ({new_AGEMA_signal_10842, new_AGEMA_signal_10841, new_AGEMA_signal_10840, SubBytesIns_Inst_Sbox_7_M46}), .b ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, new_AGEMA_signal_11500, SubBytesIns_Inst_Sbox_7_L3}), .c ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, new_AGEMA_signal_12064, SubBytesIns_Inst_Sbox_7_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L8_U1 ( .a ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, new_AGEMA_signal_10138, SubBytesIns_Inst_Sbox_7_M51}), .b ({new_AGEMA_signal_10149, new_AGEMA_signal_10148, new_AGEMA_signal_10147, SubBytesIns_Inst_Sbox_7_M59}), .c ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, new_AGEMA_signal_10867, SubBytesIns_Inst_Sbox_7_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L9_U1 ( .a ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, new_AGEMA_signal_10846, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, new_AGEMA_signal_11491, SubBytesIns_Inst_Sbox_7_M53}), .c ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, new_AGEMA_signal_12067, SubBytesIns_Inst_Sbox_7_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L10_U1 ( .a ({new_AGEMA_signal_11493, new_AGEMA_signal_11492, new_AGEMA_signal_11491, SubBytesIns_Inst_Sbox_7_M53}), .b ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, new_AGEMA_signal_11503, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, new_AGEMA_signal_12070, SubBytesIns_Inst_Sbox_7_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L11_U1 ( .a ({new_AGEMA_signal_10152, new_AGEMA_signal_10151, new_AGEMA_signal_10150, SubBytesIns_Inst_Sbox_7_M60}), .b ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, new_AGEMA_signal_11497, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, new_AGEMA_signal_12073, SubBytesIns_Inst_Sbox_7_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L12_U1 ( .a ({new_AGEMA_signal_10134, new_AGEMA_signal_10133, new_AGEMA_signal_10132, SubBytesIns_Inst_Sbox_7_M48}), .b ({new_AGEMA_signal_10140, new_AGEMA_signal_10139, new_AGEMA_signal_10138, SubBytesIns_Inst_Sbox_7_M51}), .c ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, new_AGEMA_signal_10870, SubBytesIns_Inst_Sbox_7_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L13_U1 ( .a ({new_AGEMA_signal_10137, new_AGEMA_signal_10136, new_AGEMA_signal_10135, SubBytesIns_Inst_Sbox_7_M50}), .b ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_12666, new_AGEMA_signal_12665, new_AGEMA_signal_12664, SubBytesIns_Inst_Sbox_7_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L14_U1 ( .a ({new_AGEMA_signal_10848, new_AGEMA_signal_10847, new_AGEMA_signal_10846, SubBytesIns_Inst_Sbox_7_M52}), .b ({new_AGEMA_signal_10860, new_AGEMA_signal_10859, new_AGEMA_signal_10858, SubBytesIns_Inst_Sbox_7_M61}), .c ({new_AGEMA_signal_11511, new_AGEMA_signal_11510, new_AGEMA_signal_11509, SubBytesIns_Inst_Sbox_7_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L15_U1 ( .a ({new_AGEMA_signal_10854, new_AGEMA_signal_10853, new_AGEMA_signal_10852, SubBytesIns_Inst_Sbox_7_M55}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, new_AGEMA_signal_11512, SubBytesIns_Inst_Sbox_7_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L16_U1 ( .a ({new_AGEMA_signal_10143, new_AGEMA_signal_10142, new_AGEMA_signal_10141, SubBytesIns_Inst_Sbox_7_M56}), .b ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}), .c ({new_AGEMA_signal_12669, new_AGEMA_signal_12668, new_AGEMA_signal_12667, SubBytesIns_Inst_Sbox_7_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L17_U1 ( .a ({new_AGEMA_signal_10146, new_AGEMA_signal_10145, new_AGEMA_signal_10144, SubBytesIns_Inst_Sbox_7_M57}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, new_AGEMA_signal_11515, SubBytesIns_Inst_Sbox_7_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L18_U1 ( .a ({new_AGEMA_signal_10857, new_AGEMA_signal_10856, new_AGEMA_signal_10855, SubBytesIns_Inst_Sbox_7_M58}), .b ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, new_AGEMA_signal_10867, SubBytesIns_Inst_Sbox_7_L8}), .c ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, new_AGEMA_signal_11518, SubBytesIns_Inst_Sbox_7_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L19_U1 ( .a ({new_AGEMA_signal_10863, new_AGEMA_signal_10862, new_AGEMA_signal_10861, SubBytesIns_Inst_Sbox_7_M63}), .b ({new_AGEMA_signal_11505, new_AGEMA_signal_11504, new_AGEMA_signal_11503, SubBytesIns_Inst_Sbox_7_L4}), .c ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, new_AGEMA_signal_12076, SubBytesIns_Inst_Sbox_7_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L20_U1 ( .a ({new_AGEMA_signal_12060, new_AGEMA_signal_12059, new_AGEMA_signal_12058, SubBytesIns_Inst_Sbox_7_L0}), .b ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .c ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, new_AGEMA_signal_12670, SubBytesIns_Inst_Sbox_7_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L21_U1 ( .a ({new_AGEMA_signal_10866, new_AGEMA_signal_10865, new_AGEMA_signal_10864, SubBytesIns_Inst_Sbox_7_L1}), .b ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, new_AGEMA_signal_12064, SubBytesIns_Inst_Sbox_7_L7}), .c ({new_AGEMA_signal_12675, new_AGEMA_signal_12674, new_AGEMA_signal_12673, SubBytesIns_Inst_Sbox_7_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L22_U1 ( .a ({new_AGEMA_signal_11502, new_AGEMA_signal_11501, new_AGEMA_signal_11500, SubBytesIns_Inst_Sbox_7_L3}), .b ({new_AGEMA_signal_10872, new_AGEMA_signal_10871, new_AGEMA_signal_10870, SubBytesIns_Inst_Sbox_7_L12}), .c ({new_AGEMA_signal_12081, new_AGEMA_signal_12080, new_AGEMA_signal_12079, SubBytesIns_Inst_Sbox_7_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L23_U1 ( .a ({new_AGEMA_signal_11520, new_AGEMA_signal_11519, new_AGEMA_signal_11518, SubBytesIns_Inst_Sbox_7_L18}), .b ({new_AGEMA_signal_11499, new_AGEMA_signal_11498, new_AGEMA_signal_11497, SubBytesIns_Inst_Sbox_7_L2}), .c ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, new_AGEMA_signal_12082, SubBytesIns_Inst_Sbox_7_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L24_U1 ( .a ({new_AGEMA_signal_11514, new_AGEMA_signal_11513, new_AGEMA_signal_11512, SubBytesIns_Inst_Sbox_7_L15}), .b ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, new_AGEMA_signal_12067, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_12678, new_AGEMA_signal_12677, new_AGEMA_signal_12676, SubBytesIns_Inst_Sbox_7_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L25_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, new_AGEMA_signal_12070, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, new_AGEMA_signal_12679, SubBytesIns_Inst_Sbox_7_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L26_U1 ( .a ({new_AGEMA_signal_12066, new_AGEMA_signal_12065, new_AGEMA_signal_12064, SubBytesIns_Inst_Sbox_7_L7}), .b ({new_AGEMA_signal_12069, new_AGEMA_signal_12068, new_AGEMA_signal_12067, SubBytesIns_Inst_Sbox_7_L9}), .c ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, new_AGEMA_signal_12682, SubBytesIns_Inst_Sbox_7_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L27_U1 ( .a ({new_AGEMA_signal_10869, new_AGEMA_signal_10868, new_AGEMA_signal_10867, SubBytesIns_Inst_Sbox_7_L8}), .b ({new_AGEMA_signal_12072, new_AGEMA_signal_12071, new_AGEMA_signal_12070, SubBytesIns_Inst_Sbox_7_L10}), .c ({new_AGEMA_signal_12687, new_AGEMA_signal_12686, new_AGEMA_signal_12685, SubBytesIns_Inst_Sbox_7_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L28_U1 ( .a ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, new_AGEMA_signal_12073, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_11511, new_AGEMA_signal_11510, new_AGEMA_signal_11509, SubBytesIns_Inst_Sbox_7_L14}), .c ({new_AGEMA_signal_12690, new_AGEMA_signal_12689, new_AGEMA_signal_12688, SubBytesIns_Inst_Sbox_7_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_L29_U1 ( .a ({new_AGEMA_signal_12075, new_AGEMA_signal_12074, new_AGEMA_signal_12073, SubBytesIns_Inst_Sbox_7_L11}), .b ({new_AGEMA_signal_11517, new_AGEMA_signal_11516, new_AGEMA_signal_11515, SubBytesIns_Inst_Sbox_7_L17}), .c ({new_AGEMA_signal_12693, new_AGEMA_signal_12692, new_AGEMA_signal_12691, SubBytesIns_Inst_Sbox_7_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S0_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12678, new_AGEMA_signal_12677, new_AGEMA_signal_12676, SubBytesIns_Inst_Sbox_7_L24}), .c ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S1_U1 ( .a ({new_AGEMA_signal_12669, new_AGEMA_signal_12668, new_AGEMA_signal_12667, SubBytesIns_Inst_Sbox_7_L16}), .b ({new_AGEMA_signal_12684, new_AGEMA_signal_12683, new_AGEMA_signal_12682, SubBytesIns_Inst_Sbox_7_L26}), .c ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S2_U1 ( .a ({new_AGEMA_signal_12078, new_AGEMA_signal_12077, new_AGEMA_signal_12076, SubBytesIns_Inst_Sbox_7_L19}), .b ({new_AGEMA_signal_12690, new_AGEMA_signal_12689, new_AGEMA_signal_12688, SubBytesIns_Inst_Sbox_7_L28}), .c ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S3_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12675, new_AGEMA_signal_12674, new_AGEMA_signal_12673, SubBytesIns_Inst_Sbox_7_L21}), .c ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S4_U1 ( .a ({new_AGEMA_signal_12672, new_AGEMA_signal_12671, new_AGEMA_signal_12670, SubBytesIns_Inst_Sbox_7_L20}), .b ({new_AGEMA_signal_12081, new_AGEMA_signal_12080, new_AGEMA_signal_12079, SubBytesIns_Inst_Sbox_7_L22}), .c ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S5_U1 ( .a ({new_AGEMA_signal_12681, new_AGEMA_signal_12680, new_AGEMA_signal_12679, SubBytesIns_Inst_Sbox_7_L25}), .b ({new_AGEMA_signal_12693, new_AGEMA_signal_12692, new_AGEMA_signal_12691, SubBytesIns_Inst_Sbox_7_L29}), .c ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S6_U1 ( .a ({new_AGEMA_signal_12666, new_AGEMA_signal_12665, new_AGEMA_signal_12664, SubBytesIns_Inst_Sbox_7_L13}), .b ({new_AGEMA_signal_12687, new_AGEMA_signal_12686, new_AGEMA_signal_12685, SubBytesIns_Inst_Sbox_7_L27}), .c ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_7_XOR_S7_U1 ( .a ({new_AGEMA_signal_12063, new_AGEMA_signal_12062, new_AGEMA_signal_12061, SubBytesIns_Inst_Sbox_7_L6}), .b ({new_AGEMA_signal_12084, new_AGEMA_signal_12083, new_AGEMA_signal_12082, SubBytesIns_Inst_Sbox_7_L23}), .c ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M46_U1 ( .a ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, new_AGEMA_signal_10162, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_6591, new_AGEMA_signal_6590, new_AGEMA_signal_6589, SubBytesIns_Inst_Sbox_8_T6}), .clk (clk), .r ({Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784]}), .c ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, new_AGEMA_signal_10876, SubBytesIns_Inst_Sbox_8_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M47_U1 ( .a ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_7251, new_AGEMA_signal_7250, new_AGEMA_signal_7249, SubBytesIns_Inst_Sbox_8_T8}), .clk (clk), .r ({Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790]}), .c ({new_AGEMA_signal_10167, new_AGEMA_signal_10166, new_AGEMA_signal_10165, SubBytesIns_Inst_Sbox_8_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M48_U1 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .b ({ciphertext_s3[64], ciphertext_s2[64], ciphertext_s1[64], ciphertext_s0[64]}), .clk (clk), .r ({Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796]}), .c ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, new_AGEMA_signal_10168, SubBytesIns_Inst_Sbox_8_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M49_U1 ( .a ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, new_AGEMA_signal_10159, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_6603, new_AGEMA_signal_6602, new_AGEMA_signal_6601, SubBytesIns_Inst_Sbox_8_T16}), .clk (clk), .r ({Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802]}), .c ({new_AGEMA_signal_10881, new_AGEMA_signal_10880, new_AGEMA_signal_10879, SubBytesIns_Inst_Sbox_8_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M50_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_6594, new_AGEMA_signal_6593, new_AGEMA_signal_6592, SubBytesIns_Inst_Sbox_8_T9}), .clk (clk), .r ({Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808]}), .c ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, new_AGEMA_signal_10171, SubBytesIns_Inst_Sbox_8_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M51_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_7260, new_AGEMA_signal_7259, new_AGEMA_signal_7258, SubBytesIns_Inst_Sbox_8_T17}), .clk (clk), .r ({Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814]}), .c ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, new_AGEMA_signal_10174, SubBytesIns_Inst_Sbox_8_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M52_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_6600, new_AGEMA_signal_6599, new_AGEMA_signal_6598, SubBytesIns_Inst_Sbox_8_T15}), .clk (clk), .r ({Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820]}), .c ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, new_AGEMA_signal_10882, SubBytesIns_Inst_Sbox_8_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M53_U1 ( .a ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, new_AGEMA_signal_10873, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_6612, new_AGEMA_signal_6611, new_AGEMA_signal_6610, SubBytesIns_Inst_Sbox_8_T27}), .clk (clk), .r ({Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826]}), .c ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, new_AGEMA_signal_11521, SubBytesIns_Inst_Sbox_8_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M54_U1 ( .a ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_7254, new_AGEMA_signal_7253, new_AGEMA_signal_7252, SubBytesIns_Inst_Sbox_8_T10}), .clk (clk), .r ({Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832]}), .c ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, new_AGEMA_signal_10885, SubBytesIns_Inst_Sbox_8_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M55_U1 ( .a ({new_AGEMA_signal_10164, new_AGEMA_signal_10163, new_AGEMA_signal_10162, SubBytesIns_Inst_Sbox_8_M44}), .b ({new_AGEMA_signal_6597, new_AGEMA_signal_6596, new_AGEMA_signal_6595, SubBytesIns_Inst_Sbox_8_T13}), .clk (clk), .r ({Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838]}), .c ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, new_AGEMA_signal_10888, SubBytesIns_Inst_Sbox_8_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M56_U1 ( .a ({new_AGEMA_signal_9636, new_AGEMA_signal_9635, new_AGEMA_signal_9634, SubBytesIns_Inst_Sbox_8_M40}), .b ({new_AGEMA_signal_7266, new_AGEMA_signal_7265, new_AGEMA_signal_7264, SubBytesIns_Inst_Sbox_8_T23}), .clk (clk), .r ({Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844]}), .c ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, new_AGEMA_signal_10177, SubBytesIns_Inst_Sbox_8_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M57_U1 ( .a ({new_AGEMA_signal_9633, new_AGEMA_signal_9632, new_AGEMA_signal_9631, SubBytesIns_Inst_Sbox_8_M39}), .b ({new_AGEMA_signal_6606, new_AGEMA_signal_6605, new_AGEMA_signal_6604, SubBytesIns_Inst_Sbox_8_T19}), .clk (clk), .r ({Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850]}), .c ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, new_AGEMA_signal_10180, SubBytesIns_Inst_Sbox_8_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M58_U1 ( .a ({new_AGEMA_signal_10161, new_AGEMA_signal_10160, new_AGEMA_signal_10159, SubBytesIns_Inst_Sbox_8_M43}), .b ({new_AGEMA_signal_6069, new_AGEMA_signal_6068, new_AGEMA_signal_6067, SubBytesIns_Inst_Sbox_8_T3}), .clk (clk), .r ({Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856]}), .c ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, new_AGEMA_signal_10891, SubBytesIns_Inst_Sbox_8_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M59_U1 ( .a ({new_AGEMA_signal_9630, new_AGEMA_signal_9629, new_AGEMA_signal_9628, SubBytesIns_Inst_Sbox_8_M38}), .b ({new_AGEMA_signal_6609, new_AGEMA_signal_6608, new_AGEMA_signal_6607, SubBytesIns_Inst_Sbox_8_T22}), .clk (clk), .r ({Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862]}), .c ({new_AGEMA_signal_10185, new_AGEMA_signal_10184, new_AGEMA_signal_10183, SubBytesIns_Inst_Sbox_8_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M60_U1 ( .a ({new_AGEMA_signal_9627, new_AGEMA_signal_9626, new_AGEMA_signal_9625, SubBytesIns_Inst_Sbox_8_M37}), .b ({new_AGEMA_signal_7263, new_AGEMA_signal_7262, new_AGEMA_signal_7261, SubBytesIns_Inst_Sbox_8_T20}), .clk (clk), .r ({Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868]}), .c ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, new_AGEMA_signal_10186, SubBytesIns_Inst_Sbox_8_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M61_U1 ( .a ({new_AGEMA_signal_10158, new_AGEMA_signal_10157, new_AGEMA_signal_10156, SubBytesIns_Inst_Sbox_8_M42}), .b ({new_AGEMA_signal_6063, new_AGEMA_signal_6062, new_AGEMA_signal_6061, SubBytesIns_Inst_Sbox_8_T1}), .clk (clk), .r ({Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874]}), .c ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M62_U1 ( .a ({new_AGEMA_signal_10875, new_AGEMA_signal_10874, new_AGEMA_signal_10873, SubBytesIns_Inst_Sbox_8_M45}), .b ({new_AGEMA_signal_6072, new_AGEMA_signal_6071, new_AGEMA_signal_6070, SubBytesIns_Inst_Sbox_8_T4}), .clk (clk), .r ({Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880]}), .c ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, new_AGEMA_signal_11524, SubBytesIns_Inst_Sbox_8_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_AND_M63_U1 ( .a ({new_AGEMA_signal_10155, new_AGEMA_signal_10154, new_AGEMA_signal_10153, SubBytesIns_Inst_Sbox_8_M41}), .b ({new_AGEMA_signal_6066, new_AGEMA_signal_6065, new_AGEMA_signal_6064, SubBytesIns_Inst_Sbox_8_T2}), .clk (clk), .r ({Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886]}), .c ({new_AGEMA_signal_10899, new_AGEMA_signal_10898, new_AGEMA_signal_10897, SubBytesIns_Inst_Sbox_8_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L0_U1 ( .a ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}), .b ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, new_AGEMA_signal_11524, SubBytesIns_Inst_Sbox_8_M62}), .c ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L1_U1 ( .a ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, new_AGEMA_signal_10171, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, new_AGEMA_signal_10177, SubBytesIns_Inst_Sbox_8_M56}), .c ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L2_U1 ( .a ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, new_AGEMA_signal_10876, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, new_AGEMA_signal_10168, SubBytesIns_Inst_Sbox_8_M48}), .c ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, new_AGEMA_signal_11527, SubBytesIns_Inst_Sbox_8_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L3_U1 ( .a ({new_AGEMA_signal_10167, new_AGEMA_signal_10166, new_AGEMA_signal_10165, SubBytesIns_Inst_Sbox_8_M47}), .b ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, new_AGEMA_signal_10888, SubBytesIns_Inst_Sbox_8_M55}), .c ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, new_AGEMA_signal_11530, SubBytesIns_Inst_Sbox_8_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L4_U1 ( .a ({new_AGEMA_signal_10887, new_AGEMA_signal_10886, new_AGEMA_signal_10885, SubBytesIns_Inst_Sbox_8_M54}), .b ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, new_AGEMA_signal_10891, SubBytesIns_Inst_Sbox_8_M58}), .c ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, new_AGEMA_signal_11533, SubBytesIns_Inst_Sbox_8_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L5_U1 ( .a ({new_AGEMA_signal_10881, new_AGEMA_signal_10880, new_AGEMA_signal_10879, SubBytesIns_Inst_Sbox_8_M49}), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, new_AGEMA_signal_11536, SubBytesIns_Inst_Sbox_8_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L6_U1 ( .a ({new_AGEMA_signal_11526, new_AGEMA_signal_11525, new_AGEMA_signal_11524, SubBytesIns_Inst_Sbox_8_M62}), .b ({new_AGEMA_signal_11538, new_AGEMA_signal_11537, new_AGEMA_signal_11536, SubBytesIns_Inst_Sbox_8_L5}), .c ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L7_U1 ( .a ({new_AGEMA_signal_10878, new_AGEMA_signal_10877, new_AGEMA_signal_10876, SubBytesIns_Inst_Sbox_8_M46}), .b ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, new_AGEMA_signal_11530, SubBytesIns_Inst_Sbox_8_L3}), .c ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, new_AGEMA_signal_12091, SubBytesIns_Inst_Sbox_8_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L8_U1 ( .a ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, new_AGEMA_signal_10174, SubBytesIns_Inst_Sbox_8_M51}), .b ({new_AGEMA_signal_10185, new_AGEMA_signal_10184, new_AGEMA_signal_10183, SubBytesIns_Inst_Sbox_8_M59}), .c ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, new_AGEMA_signal_10903, SubBytesIns_Inst_Sbox_8_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L9_U1 ( .a ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, new_AGEMA_signal_10882, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, new_AGEMA_signal_11521, SubBytesIns_Inst_Sbox_8_M53}), .c ({new_AGEMA_signal_12096, new_AGEMA_signal_12095, new_AGEMA_signal_12094, SubBytesIns_Inst_Sbox_8_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L10_U1 ( .a ({new_AGEMA_signal_11523, new_AGEMA_signal_11522, new_AGEMA_signal_11521, SubBytesIns_Inst_Sbox_8_M53}), .b ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, new_AGEMA_signal_11533, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, new_AGEMA_signal_12097, SubBytesIns_Inst_Sbox_8_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L11_U1 ( .a ({new_AGEMA_signal_10188, new_AGEMA_signal_10187, new_AGEMA_signal_10186, SubBytesIns_Inst_Sbox_8_M60}), .b ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, new_AGEMA_signal_11527, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, new_AGEMA_signal_12100, SubBytesIns_Inst_Sbox_8_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L12_U1 ( .a ({new_AGEMA_signal_10170, new_AGEMA_signal_10169, new_AGEMA_signal_10168, SubBytesIns_Inst_Sbox_8_M48}), .b ({new_AGEMA_signal_10176, new_AGEMA_signal_10175, new_AGEMA_signal_10174, SubBytesIns_Inst_Sbox_8_M51}), .c ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, new_AGEMA_signal_10906, SubBytesIns_Inst_Sbox_8_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L13_U1 ( .a ({new_AGEMA_signal_10173, new_AGEMA_signal_10172, new_AGEMA_signal_10171, SubBytesIns_Inst_Sbox_8_M50}), .b ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_12699, new_AGEMA_signal_12698, new_AGEMA_signal_12697, SubBytesIns_Inst_Sbox_8_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L14_U1 ( .a ({new_AGEMA_signal_10884, new_AGEMA_signal_10883, new_AGEMA_signal_10882, SubBytesIns_Inst_Sbox_8_M52}), .b ({new_AGEMA_signal_10896, new_AGEMA_signal_10895, new_AGEMA_signal_10894, SubBytesIns_Inst_Sbox_8_M61}), .c ({new_AGEMA_signal_11541, new_AGEMA_signal_11540, new_AGEMA_signal_11539, SubBytesIns_Inst_Sbox_8_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L15_U1 ( .a ({new_AGEMA_signal_10890, new_AGEMA_signal_10889, new_AGEMA_signal_10888, SubBytesIns_Inst_Sbox_8_M55}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, new_AGEMA_signal_11542, SubBytesIns_Inst_Sbox_8_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L16_U1 ( .a ({new_AGEMA_signal_10179, new_AGEMA_signal_10178, new_AGEMA_signal_10177, SubBytesIns_Inst_Sbox_8_M56}), .b ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}), .c ({new_AGEMA_signal_12702, new_AGEMA_signal_12701, new_AGEMA_signal_12700, SubBytesIns_Inst_Sbox_8_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L17_U1 ( .a ({new_AGEMA_signal_10182, new_AGEMA_signal_10181, new_AGEMA_signal_10180, SubBytesIns_Inst_Sbox_8_M57}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_11547, new_AGEMA_signal_11546, new_AGEMA_signal_11545, SubBytesIns_Inst_Sbox_8_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L18_U1 ( .a ({new_AGEMA_signal_10893, new_AGEMA_signal_10892, new_AGEMA_signal_10891, SubBytesIns_Inst_Sbox_8_M58}), .b ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, new_AGEMA_signal_10903, SubBytesIns_Inst_Sbox_8_L8}), .c ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, new_AGEMA_signal_11548, SubBytesIns_Inst_Sbox_8_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L19_U1 ( .a ({new_AGEMA_signal_10899, new_AGEMA_signal_10898, new_AGEMA_signal_10897, SubBytesIns_Inst_Sbox_8_M63}), .b ({new_AGEMA_signal_11535, new_AGEMA_signal_11534, new_AGEMA_signal_11533, SubBytesIns_Inst_Sbox_8_L4}), .c ({new_AGEMA_signal_12105, new_AGEMA_signal_12104, new_AGEMA_signal_12103, SubBytesIns_Inst_Sbox_8_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L20_U1 ( .a ({new_AGEMA_signal_12087, new_AGEMA_signal_12086, new_AGEMA_signal_12085, SubBytesIns_Inst_Sbox_8_L0}), .b ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .c ({new_AGEMA_signal_12705, new_AGEMA_signal_12704, new_AGEMA_signal_12703, SubBytesIns_Inst_Sbox_8_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L21_U1 ( .a ({new_AGEMA_signal_10902, new_AGEMA_signal_10901, new_AGEMA_signal_10900, SubBytesIns_Inst_Sbox_8_L1}), .b ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, new_AGEMA_signal_12091, SubBytesIns_Inst_Sbox_8_L7}), .c ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, new_AGEMA_signal_12706, SubBytesIns_Inst_Sbox_8_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L22_U1 ( .a ({new_AGEMA_signal_11532, new_AGEMA_signal_11531, new_AGEMA_signal_11530, SubBytesIns_Inst_Sbox_8_L3}), .b ({new_AGEMA_signal_10908, new_AGEMA_signal_10907, new_AGEMA_signal_10906, SubBytesIns_Inst_Sbox_8_L12}), .c ({new_AGEMA_signal_12108, new_AGEMA_signal_12107, new_AGEMA_signal_12106, SubBytesIns_Inst_Sbox_8_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L23_U1 ( .a ({new_AGEMA_signal_11550, new_AGEMA_signal_11549, new_AGEMA_signal_11548, SubBytesIns_Inst_Sbox_8_L18}), .b ({new_AGEMA_signal_11529, new_AGEMA_signal_11528, new_AGEMA_signal_11527, SubBytesIns_Inst_Sbox_8_L2}), .c ({new_AGEMA_signal_12111, new_AGEMA_signal_12110, new_AGEMA_signal_12109, SubBytesIns_Inst_Sbox_8_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L24_U1 ( .a ({new_AGEMA_signal_11544, new_AGEMA_signal_11543, new_AGEMA_signal_11542, SubBytesIns_Inst_Sbox_8_L15}), .b ({new_AGEMA_signal_12096, new_AGEMA_signal_12095, new_AGEMA_signal_12094, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, new_AGEMA_signal_12709, SubBytesIns_Inst_Sbox_8_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L25_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, new_AGEMA_signal_12097, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_12714, new_AGEMA_signal_12713, new_AGEMA_signal_12712, SubBytesIns_Inst_Sbox_8_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L26_U1 ( .a ({new_AGEMA_signal_12093, new_AGEMA_signal_12092, new_AGEMA_signal_12091, SubBytesIns_Inst_Sbox_8_L7}), .b ({new_AGEMA_signal_12096, new_AGEMA_signal_12095, new_AGEMA_signal_12094, SubBytesIns_Inst_Sbox_8_L9}), .c ({new_AGEMA_signal_12717, new_AGEMA_signal_12716, new_AGEMA_signal_12715, SubBytesIns_Inst_Sbox_8_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L27_U1 ( .a ({new_AGEMA_signal_10905, new_AGEMA_signal_10904, new_AGEMA_signal_10903, SubBytesIns_Inst_Sbox_8_L8}), .b ({new_AGEMA_signal_12099, new_AGEMA_signal_12098, new_AGEMA_signal_12097, SubBytesIns_Inst_Sbox_8_L10}), .c ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, new_AGEMA_signal_12718, SubBytesIns_Inst_Sbox_8_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L28_U1 ( .a ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, new_AGEMA_signal_12100, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_11541, new_AGEMA_signal_11540, new_AGEMA_signal_11539, SubBytesIns_Inst_Sbox_8_L14}), .c ({new_AGEMA_signal_12723, new_AGEMA_signal_12722, new_AGEMA_signal_12721, SubBytesIns_Inst_Sbox_8_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_L29_U1 ( .a ({new_AGEMA_signal_12102, new_AGEMA_signal_12101, new_AGEMA_signal_12100, SubBytesIns_Inst_Sbox_8_L11}), .b ({new_AGEMA_signal_11547, new_AGEMA_signal_11546, new_AGEMA_signal_11545, SubBytesIns_Inst_Sbox_8_L17}), .c ({new_AGEMA_signal_12726, new_AGEMA_signal_12725, new_AGEMA_signal_12724, SubBytesIns_Inst_Sbox_8_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S0_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12711, new_AGEMA_signal_12710, new_AGEMA_signal_12709, SubBytesIns_Inst_Sbox_8_L24}), .c ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S1_U1 ( .a ({new_AGEMA_signal_12702, new_AGEMA_signal_12701, new_AGEMA_signal_12700, SubBytesIns_Inst_Sbox_8_L16}), .b ({new_AGEMA_signal_12717, new_AGEMA_signal_12716, new_AGEMA_signal_12715, SubBytesIns_Inst_Sbox_8_L26}), .c ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S2_U1 ( .a ({new_AGEMA_signal_12105, new_AGEMA_signal_12104, new_AGEMA_signal_12103, SubBytesIns_Inst_Sbox_8_L19}), .b ({new_AGEMA_signal_12723, new_AGEMA_signal_12722, new_AGEMA_signal_12721, SubBytesIns_Inst_Sbox_8_L28}), .c ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S3_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12708, new_AGEMA_signal_12707, new_AGEMA_signal_12706, SubBytesIns_Inst_Sbox_8_L21}), .c ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S4_U1 ( .a ({new_AGEMA_signal_12705, new_AGEMA_signal_12704, new_AGEMA_signal_12703, SubBytesIns_Inst_Sbox_8_L20}), .b ({new_AGEMA_signal_12108, new_AGEMA_signal_12107, new_AGEMA_signal_12106, SubBytesIns_Inst_Sbox_8_L22}), .c ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S5_U1 ( .a ({new_AGEMA_signal_12714, new_AGEMA_signal_12713, new_AGEMA_signal_12712, SubBytesIns_Inst_Sbox_8_L25}), .b ({new_AGEMA_signal_12726, new_AGEMA_signal_12725, new_AGEMA_signal_12724, SubBytesIns_Inst_Sbox_8_L29}), .c ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S6_U1 ( .a ({new_AGEMA_signal_12699, new_AGEMA_signal_12698, new_AGEMA_signal_12697, SubBytesIns_Inst_Sbox_8_L13}), .b ({new_AGEMA_signal_12720, new_AGEMA_signal_12719, new_AGEMA_signal_12718, SubBytesIns_Inst_Sbox_8_L27}), .c ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_8_XOR_S7_U1 ( .a ({new_AGEMA_signal_12090, new_AGEMA_signal_12089, new_AGEMA_signal_12088, SubBytesIns_Inst_Sbox_8_L6}), .b ({new_AGEMA_signal_12111, new_AGEMA_signal_12110, new_AGEMA_signal_12109, SubBytesIns_Inst_Sbox_8_L23}), .c ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M46_U1 ( .a ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, new_AGEMA_signal_10198, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_6615, new_AGEMA_signal_6614, new_AGEMA_signal_6613, SubBytesIns_Inst_Sbox_9_T6}), .clk (clk), .r ({Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892]}), .c ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, new_AGEMA_signal_10912, SubBytesIns_Inst_Sbox_9_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M47_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_7290, new_AGEMA_signal_7289, new_AGEMA_signal_7288, SubBytesIns_Inst_Sbox_9_T8}), .clk (clk), .r ({Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898]}), .c ({new_AGEMA_signal_10203, new_AGEMA_signal_10202, new_AGEMA_signal_10201, SubBytesIns_Inst_Sbox_9_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M48_U1 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .b ({ciphertext_s3[72], ciphertext_s2[72], ciphertext_s1[72], ciphertext_s0[72]}), .clk (clk), .r ({Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904]}), .c ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, new_AGEMA_signal_10204, SubBytesIns_Inst_Sbox_9_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M49_U1 ( .a ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, new_AGEMA_signal_10195, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_6627, new_AGEMA_signal_6626, new_AGEMA_signal_6625, SubBytesIns_Inst_Sbox_9_T16}), .clk (clk), .r ({Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910]}), .c ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, new_AGEMA_signal_10915, SubBytesIns_Inst_Sbox_9_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M50_U1 ( .a ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_6618, new_AGEMA_signal_6617, new_AGEMA_signal_6616, SubBytesIns_Inst_Sbox_9_T9}), .clk (clk), .r ({Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916]}), .c ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, new_AGEMA_signal_10207, SubBytesIns_Inst_Sbox_9_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M51_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_7299, new_AGEMA_signal_7298, new_AGEMA_signal_7297, SubBytesIns_Inst_Sbox_9_T17}), .clk (clk), .r ({Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922]}), .c ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, new_AGEMA_signal_10210, SubBytesIns_Inst_Sbox_9_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M52_U1 ( .a ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_6624, new_AGEMA_signal_6623, new_AGEMA_signal_6622, SubBytesIns_Inst_Sbox_9_T15}), .clk (clk), .r ({Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928]}), .c ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, new_AGEMA_signal_10918, SubBytesIns_Inst_Sbox_9_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M53_U1 ( .a ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, new_AGEMA_signal_10909, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_6636, new_AGEMA_signal_6635, new_AGEMA_signal_6634, SubBytesIns_Inst_Sbox_9_T27}), .clk (clk), .r ({Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934]}), .c ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, new_AGEMA_signal_11551, SubBytesIns_Inst_Sbox_9_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M54_U1 ( .a ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_7293, new_AGEMA_signal_7292, new_AGEMA_signal_7291, SubBytesIns_Inst_Sbox_9_T10}), .clk (clk), .r ({Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940]}), .c ({new_AGEMA_signal_10923, new_AGEMA_signal_10922, new_AGEMA_signal_10921, SubBytesIns_Inst_Sbox_9_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M55_U1 ( .a ({new_AGEMA_signal_10200, new_AGEMA_signal_10199, new_AGEMA_signal_10198, SubBytesIns_Inst_Sbox_9_M44}), .b ({new_AGEMA_signal_6621, new_AGEMA_signal_6620, new_AGEMA_signal_6619, SubBytesIns_Inst_Sbox_9_T13}), .clk (clk), .r ({Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946]}), .c ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, new_AGEMA_signal_10924, SubBytesIns_Inst_Sbox_9_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M56_U1 ( .a ({new_AGEMA_signal_9648, new_AGEMA_signal_9647, new_AGEMA_signal_9646, SubBytesIns_Inst_Sbox_9_M40}), .b ({new_AGEMA_signal_7305, new_AGEMA_signal_7304, new_AGEMA_signal_7303, SubBytesIns_Inst_Sbox_9_T23}), .clk (clk), .r ({Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952]}), .c ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, new_AGEMA_signal_10213, SubBytesIns_Inst_Sbox_9_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M57_U1 ( .a ({new_AGEMA_signal_9645, new_AGEMA_signal_9644, new_AGEMA_signal_9643, SubBytesIns_Inst_Sbox_9_M39}), .b ({new_AGEMA_signal_6630, new_AGEMA_signal_6629, new_AGEMA_signal_6628, SubBytesIns_Inst_Sbox_9_T19}), .clk (clk), .r ({Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958]}), .c ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, new_AGEMA_signal_10216, SubBytesIns_Inst_Sbox_9_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M58_U1 ( .a ({new_AGEMA_signal_10197, new_AGEMA_signal_10196, new_AGEMA_signal_10195, SubBytesIns_Inst_Sbox_9_M43}), .b ({new_AGEMA_signal_6099, new_AGEMA_signal_6098, new_AGEMA_signal_6097, SubBytesIns_Inst_Sbox_9_T3}), .clk (clk), .r ({Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964]}), .c ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, new_AGEMA_signal_10927, SubBytesIns_Inst_Sbox_9_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M59_U1 ( .a ({new_AGEMA_signal_9642, new_AGEMA_signal_9641, new_AGEMA_signal_9640, SubBytesIns_Inst_Sbox_9_M38}), .b ({new_AGEMA_signal_6633, new_AGEMA_signal_6632, new_AGEMA_signal_6631, SubBytesIns_Inst_Sbox_9_T22}), .clk (clk), .r ({Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970]}), .c ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, new_AGEMA_signal_10219, SubBytesIns_Inst_Sbox_9_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M60_U1 ( .a ({new_AGEMA_signal_9639, new_AGEMA_signal_9638, new_AGEMA_signal_9637, SubBytesIns_Inst_Sbox_9_M37}), .b ({new_AGEMA_signal_7302, new_AGEMA_signal_7301, new_AGEMA_signal_7300, SubBytesIns_Inst_Sbox_9_T20}), .clk (clk), .r ({Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976]}), .c ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, new_AGEMA_signal_10222, SubBytesIns_Inst_Sbox_9_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M61_U1 ( .a ({new_AGEMA_signal_10194, new_AGEMA_signal_10193, new_AGEMA_signal_10192, SubBytesIns_Inst_Sbox_9_M42}), .b ({new_AGEMA_signal_6093, new_AGEMA_signal_6092, new_AGEMA_signal_6091, SubBytesIns_Inst_Sbox_9_T1}), .clk (clk), .r ({Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982]}), .c ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M62_U1 ( .a ({new_AGEMA_signal_10911, new_AGEMA_signal_10910, new_AGEMA_signal_10909, SubBytesIns_Inst_Sbox_9_M45}), .b ({new_AGEMA_signal_6102, new_AGEMA_signal_6101, new_AGEMA_signal_6100, SubBytesIns_Inst_Sbox_9_T4}), .clk (clk), .r ({Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988]}), .c ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, new_AGEMA_signal_11554, SubBytesIns_Inst_Sbox_9_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_AND_M63_U1 ( .a ({new_AGEMA_signal_10191, new_AGEMA_signal_10190, new_AGEMA_signal_10189, SubBytesIns_Inst_Sbox_9_M41}), .b ({new_AGEMA_signal_6096, new_AGEMA_signal_6095, new_AGEMA_signal_6094, SubBytesIns_Inst_Sbox_9_T2}), .clk (clk), .r ({Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994]}), .c ({new_AGEMA_signal_10935, new_AGEMA_signal_10934, new_AGEMA_signal_10933, SubBytesIns_Inst_Sbox_9_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L0_U1 ( .a ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}), .b ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, new_AGEMA_signal_11554, SubBytesIns_Inst_Sbox_9_M62}), .c ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L1_U1 ( .a ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, new_AGEMA_signal_10207, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, new_AGEMA_signal_10213, SubBytesIns_Inst_Sbox_9_M56}), .c ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L2_U1 ( .a ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, new_AGEMA_signal_10912, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, new_AGEMA_signal_10204, SubBytesIns_Inst_Sbox_9_M48}), .c ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, new_AGEMA_signal_11557, SubBytesIns_Inst_Sbox_9_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L3_U1 ( .a ({new_AGEMA_signal_10203, new_AGEMA_signal_10202, new_AGEMA_signal_10201, SubBytesIns_Inst_Sbox_9_M47}), .b ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, new_AGEMA_signal_10924, SubBytesIns_Inst_Sbox_9_M55}), .c ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, new_AGEMA_signal_11560, SubBytesIns_Inst_Sbox_9_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L4_U1 ( .a ({new_AGEMA_signal_10923, new_AGEMA_signal_10922, new_AGEMA_signal_10921, SubBytesIns_Inst_Sbox_9_M54}), .b ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, new_AGEMA_signal_10927, SubBytesIns_Inst_Sbox_9_M58}), .c ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, new_AGEMA_signal_11563, SubBytesIns_Inst_Sbox_9_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L5_U1 ( .a ({new_AGEMA_signal_10917, new_AGEMA_signal_10916, new_AGEMA_signal_10915, SubBytesIns_Inst_Sbox_9_M49}), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, new_AGEMA_signal_11566, SubBytesIns_Inst_Sbox_9_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L6_U1 ( .a ({new_AGEMA_signal_11556, new_AGEMA_signal_11555, new_AGEMA_signal_11554, SubBytesIns_Inst_Sbox_9_M62}), .b ({new_AGEMA_signal_11568, new_AGEMA_signal_11567, new_AGEMA_signal_11566, SubBytesIns_Inst_Sbox_9_L5}), .c ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L7_U1 ( .a ({new_AGEMA_signal_10914, new_AGEMA_signal_10913, new_AGEMA_signal_10912, SubBytesIns_Inst_Sbox_9_M46}), .b ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, new_AGEMA_signal_11560, SubBytesIns_Inst_Sbox_9_L3}), .c ({new_AGEMA_signal_12120, new_AGEMA_signal_12119, new_AGEMA_signal_12118, SubBytesIns_Inst_Sbox_9_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L8_U1 ( .a ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, new_AGEMA_signal_10210, SubBytesIns_Inst_Sbox_9_M51}), .b ({new_AGEMA_signal_10221, new_AGEMA_signal_10220, new_AGEMA_signal_10219, SubBytesIns_Inst_Sbox_9_M59}), .c ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, new_AGEMA_signal_10939, SubBytesIns_Inst_Sbox_9_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L9_U1 ( .a ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, new_AGEMA_signal_10918, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, new_AGEMA_signal_11551, SubBytesIns_Inst_Sbox_9_M53}), .c ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, new_AGEMA_signal_12121, SubBytesIns_Inst_Sbox_9_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L10_U1 ( .a ({new_AGEMA_signal_11553, new_AGEMA_signal_11552, new_AGEMA_signal_11551, SubBytesIns_Inst_Sbox_9_M53}), .b ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, new_AGEMA_signal_11563, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, new_AGEMA_signal_12124, SubBytesIns_Inst_Sbox_9_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L11_U1 ( .a ({new_AGEMA_signal_10224, new_AGEMA_signal_10223, new_AGEMA_signal_10222, SubBytesIns_Inst_Sbox_9_M60}), .b ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, new_AGEMA_signal_11557, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, new_AGEMA_signal_12127, SubBytesIns_Inst_Sbox_9_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L12_U1 ( .a ({new_AGEMA_signal_10206, new_AGEMA_signal_10205, new_AGEMA_signal_10204, SubBytesIns_Inst_Sbox_9_M48}), .b ({new_AGEMA_signal_10212, new_AGEMA_signal_10211, new_AGEMA_signal_10210, SubBytesIns_Inst_Sbox_9_M51}), .c ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, new_AGEMA_signal_10942, SubBytesIns_Inst_Sbox_9_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L13_U1 ( .a ({new_AGEMA_signal_10209, new_AGEMA_signal_10208, new_AGEMA_signal_10207, SubBytesIns_Inst_Sbox_9_M50}), .b ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, new_AGEMA_signal_12730, SubBytesIns_Inst_Sbox_9_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L14_U1 ( .a ({new_AGEMA_signal_10920, new_AGEMA_signal_10919, new_AGEMA_signal_10918, SubBytesIns_Inst_Sbox_9_M52}), .b ({new_AGEMA_signal_10932, new_AGEMA_signal_10931, new_AGEMA_signal_10930, SubBytesIns_Inst_Sbox_9_M61}), .c ({new_AGEMA_signal_11571, new_AGEMA_signal_11570, new_AGEMA_signal_11569, SubBytesIns_Inst_Sbox_9_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L15_U1 ( .a ({new_AGEMA_signal_10926, new_AGEMA_signal_10925, new_AGEMA_signal_10924, SubBytesIns_Inst_Sbox_9_M55}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, new_AGEMA_signal_11572, SubBytesIns_Inst_Sbox_9_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L16_U1 ( .a ({new_AGEMA_signal_10215, new_AGEMA_signal_10214, new_AGEMA_signal_10213, SubBytesIns_Inst_Sbox_9_M56}), .b ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}), .c ({new_AGEMA_signal_12735, new_AGEMA_signal_12734, new_AGEMA_signal_12733, SubBytesIns_Inst_Sbox_9_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L17_U1 ( .a ({new_AGEMA_signal_10218, new_AGEMA_signal_10217, new_AGEMA_signal_10216, SubBytesIns_Inst_Sbox_9_M57}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_11577, new_AGEMA_signal_11576, new_AGEMA_signal_11575, SubBytesIns_Inst_Sbox_9_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L18_U1 ( .a ({new_AGEMA_signal_10929, new_AGEMA_signal_10928, new_AGEMA_signal_10927, SubBytesIns_Inst_Sbox_9_M58}), .b ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, new_AGEMA_signal_10939, SubBytesIns_Inst_Sbox_9_L8}), .c ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, new_AGEMA_signal_11578, SubBytesIns_Inst_Sbox_9_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L19_U1 ( .a ({new_AGEMA_signal_10935, new_AGEMA_signal_10934, new_AGEMA_signal_10933, SubBytesIns_Inst_Sbox_9_M63}), .b ({new_AGEMA_signal_11565, new_AGEMA_signal_11564, new_AGEMA_signal_11563, SubBytesIns_Inst_Sbox_9_L4}), .c ({new_AGEMA_signal_12132, new_AGEMA_signal_12131, new_AGEMA_signal_12130, SubBytesIns_Inst_Sbox_9_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L20_U1 ( .a ({new_AGEMA_signal_12114, new_AGEMA_signal_12113, new_AGEMA_signal_12112, SubBytesIns_Inst_Sbox_9_L0}), .b ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .c ({new_AGEMA_signal_12738, new_AGEMA_signal_12737, new_AGEMA_signal_12736, SubBytesIns_Inst_Sbox_9_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L21_U1 ( .a ({new_AGEMA_signal_10938, new_AGEMA_signal_10937, new_AGEMA_signal_10936, SubBytesIns_Inst_Sbox_9_L1}), .b ({new_AGEMA_signal_12120, new_AGEMA_signal_12119, new_AGEMA_signal_12118, SubBytesIns_Inst_Sbox_9_L7}), .c ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, new_AGEMA_signal_12739, SubBytesIns_Inst_Sbox_9_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L22_U1 ( .a ({new_AGEMA_signal_11562, new_AGEMA_signal_11561, new_AGEMA_signal_11560, SubBytesIns_Inst_Sbox_9_L3}), .b ({new_AGEMA_signal_10944, new_AGEMA_signal_10943, new_AGEMA_signal_10942, SubBytesIns_Inst_Sbox_9_L12}), .c ({new_AGEMA_signal_12135, new_AGEMA_signal_12134, new_AGEMA_signal_12133, SubBytesIns_Inst_Sbox_9_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L23_U1 ( .a ({new_AGEMA_signal_11580, new_AGEMA_signal_11579, new_AGEMA_signal_11578, SubBytesIns_Inst_Sbox_9_L18}), .b ({new_AGEMA_signal_11559, new_AGEMA_signal_11558, new_AGEMA_signal_11557, SubBytesIns_Inst_Sbox_9_L2}), .c ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, new_AGEMA_signal_12136, SubBytesIns_Inst_Sbox_9_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L24_U1 ( .a ({new_AGEMA_signal_11574, new_AGEMA_signal_11573, new_AGEMA_signal_11572, SubBytesIns_Inst_Sbox_9_L15}), .b ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, new_AGEMA_signal_12121, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, new_AGEMA_signal_12742, SubBytesIns_Inst_Sbox_9_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L25_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, new_AGEMA_signal_12124, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_12747, new_AGEMA_signal_12746, new_AGEMA_signal_12745, SubBytesIns_Inst_Sbox_9_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L26_U1 ( .a ({new_AGEMA_signal_12120, new_AGEMA_signal_12119, new_AGEMA_signal_12118, SubBytesIns_Inst_Sbox_9_L7}), .b ({new_AGEMA_signal_12123, new_AGEMA_signal_12122, new_AGEMA_signal_12121, SubBytesIns_Inst_Sbox_9_L9}), .c ({new_AGEMA_signal_12750, new_AGEMA_signal_12749, new_AGEMA_signal_12748, SubBytesIns_Inst_Sbox_9_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L27_U1 ( .a ({new_AGEMA_signal_10941, new_AGEMA_signal_10940, new_AGEMA_signal_10939, SubBytesIns_Inst_Sbox_9_L8}), .b ({new_AGEMA_signal_12126, new_AGEMA_signal_12125, new_AGEMA_signal_12124, SubBytesIns_Inst_Sbox_9_L10}), .c ({new_AGEMA_signal_12753, new_AGEMA_signal_12752, new_AGEMA_signal_12751, SubBytesIns_Inst_Sbox_9_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L28_U1 ( .a ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, new_AGEMA_signal_12127, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_11571, new_AGEMA_signal_11570, new_AGEMA_signal_11569, SubBytesIns_Inst_Sbox_9_L14}), .c ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, new_AGEMA_signal_12754, SubBytesIns_Inst_Sbox_9_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_L29_U1 ( .a ({new_AGEMA_signal_12129, new_AGEMA_signal_12128, new_AGEMA_signal_12127, SubBytesIns_Inst_Sbox_9_L11}), .b ({new_AGEMA_signal_11577, new_AGEMA_signal_11576, new_AGEMA_signal_11575, SubBytesIns_Inst_Sbox_9_L17}), .c ({new_AGEMA_signal_12759, new_AGEMA_signal_12758, new_AGEMA_signal_12757, SubBytesIns_Inst_Sbox_9_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S0_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12744, new_AGEMA_signal_12743, new_AGEMA_signal_12742, SubBytesIns_Inst_Sbox_9_L24}), .c ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S1_U1 ( .a ({new_AGEMA_signal_12735, new_AGEMA_signal_12734, new_AGEMA_signal_12733, SubBytesIns_Inst_Sbox_9_L16}), .b ({new_AGEMA_signal_12750, new_AGEMA_signal_12749, new_AGEMA_signal_12748, SubBytesIns_Inst_Sbox_9_L26}), .c ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S2_U1 ( .a ({new_AGEMA_signal_12132, new_AGEMA_signal_12131, new_AGEMA_signal_12130, SubBytesIns_Inst_Sbox_9_L19}), .b ({new_AGEMA_signal_12756, new_AGEMA_signal_12755, new_AGEMA_signal_12754, SubBytesIns_Inst_Sbox_9_L28}), .c ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S3_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12741, new_AGEMA_signal_12740, new_AGEMA_signal_12739, SubBytesIns_Inst_Sbox_9_L21}), .c ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S4_U1 ( .a ({new_AGEMA_signal_12738, new_AGEMA_signal_12737, new_AGEMA_signal_12736, SubBytesIns_Inst_Sbox_9_L20}), .b ({new_AGEMA_signal_12135, new_AGEMA_signal_12134, new_AGEMA_signal_12133, SubBytesIns_Inst_Sbox_9_L22}), .c ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S5_U1 ( .a ({new_AGEMA_signal_12747, new_AGEMA_signal_12746, new_AGEMA_signal_12745, SubBytesIns_Inst_Sbox_9_L25}), .b ({new_AGEMA_signal_12759, new_AGEMA_signal_12758, new_AGEMA_signal_12757, SubBytesIns_Inst_Sbox_9_L29}), .c ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S6_U1 ( .a ({new_AGEMA_signal_12732, new_AGEMA_signal_12731, new_AGEMA_signal_12730, SubBytesIns_Inst_Sbox_9_L13}), .b ({new_AGEMA_signal_12753, new_AGEMA_signal_12752, new_AGEMA_signal_12751, SubBytesIns_Inst_Sbox_9_L27}), .c ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_9_XOR_S7_U1 ( .a ({new_AGEMA_signal_12117, new_AGEMA_signal_12116, new_AGEMA_signal_12115, SubBytesIns_Inst_Sbox_9_L6}), .b ({new_AGEMA_signal_12138, new_AGEMA_signal_12137, new_AGEMA_signal_12136, SubBytesIns_Inst_Sbox_9_L23}), .c ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M46_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, new_AGEMA_signal_10234, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_6639, new_AGEMA_signal_6638, new_AGEMA_signal_6637, SubBytesIns_Inst_Sbox_10_T6}), .clk (clk), .r ({Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000]}), .c ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, new_AGEMA_signal_10948, SubBytesIns_Inst_Sbox_10_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M47_U1 ( .a ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_7329, new_AGEMA_signal_7328, new_AGEMA_signal_7327, SubBytesIns_Inst_Sbox_10_T8}), .clk (clk), .r ({Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006]}), .c ({new_AGEMA_signal_10239, new_AGEMA_signal_10238, new_AGEMA_signal_10237, SubBytesIns_Inst_Sbox_10_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M48_U1 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .b ({ciphertext_s3[80], ciphertext_s2[80], ciphertext_s1[80], ciphertext_s0[80]}), .clk (clk), .r ({Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012]}), .c ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, new_AGEMA_signal_10240, SubBytesIns_Inst_Sbox_10_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M49_U1 ( .a ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, new_AGEMA_signal_10231, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_6651, new_AGEMA_signal_6650, new_AGEMA_signal_6649, SubBytesIns_Inst_Sbox_10_T16}), .clk (clk), .r ({Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018]}), .c ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, new_AGEMA_signal_10951, SubBytesIns_Inst_Sbox_10_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M50_U1 ( .a ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_6642, new_AGEMA_signal_6641, new_AGEMA_signal_6640, SubBytesIns_Inst_Sbox_10_T9}), .clk (clk), .r ({Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024]}), .c ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, new_AGEMA_signal_10243, SubBytesIns_Inst_Sbox_10_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M51_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_7338, new_AGEMA_signal_7337, new_AGEMA_signal_7336, SubBytesIns_Inst_Sbox_10_T17}), .clk (clk), .r ({Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030]}), .c ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, new_AGEMA_signal_10246, SubBytesIns_Inst_Sbox_10_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M52_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_6648, new_AGEMA_signal_6647, new_AGEMA_signal_6646, SubBytesIns_Inst_Sbox_10_T15}), .clk (clk), .r ({Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036]}), .c ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, new_AGEMA_signal_10954, SubBytesIns_Inst_Sbox_10_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M53_U1 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, new_AGEMA_signal_10945, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_6660, new_AGEMA_signal_6659, new_AGEMA_signal_6658, SubBytesIns_Inst_Sbox_10_T27}), .clk (clk), .r ({Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042]}), .c ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, new_AGEMA_signal_11581, SubBytesIns_Inst_Sbox_10_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M54_U1 ( .a ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_7332, new_AGEMA_signal_7331, new_AGEMA_signal_7330, SubBytesIns_Inst_Sbox_10_T10}), .clk (clk), .r ({Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048]}), .c ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, new_AGEMA_signal_10957, SubBytesIns_Inst_Sbox_10_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M55_U1 ( .a ({new_AGEMA_signal_10236, new_AGEMA_signal_10235, new_AGEMA_signal_10234, SubBytesIns_Inst_Sbox_10_M44}), .b ({new_AGEMA_signal_6645, new_AGEMA_signal_6644, new_AGEMA_signal_6643, SubBytesIns_Inst_Sbox_10_T13}), .clk (clk), .r ({Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054]}), .c ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, new_AGEMA_signal_10960, SubBytesIns_Inst_Sbox_10_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M56_U1 ( .a ({new_AGEMA_signal_9660, new_AGEMA_signal_9659, new_AGEMA_signal_9658, SubBytesIns_Inst_Sbox_10_M40}), .b ({new_AGEMA_signal_7344, new_AGEMA_signal_7343, new_AGEMA_signal_7342, SubBytesIns_Inst_Sbox_10_T23}), .clk (clk), .r ({Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060]}), .c ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, new_AGEMA_signal_10249, SubBytesIns_Inst_Sbox_10_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M57_U1 ( .a ({new_AGEMA_signal_9657, new_AGEMA_signal_9656, new_AGEMA_signal_9655, SubBytesIns_Inst_Sbox_10_M39}), .b ({new_AGEMA_signal_6654, new_AGEMA_signal_6653, new_AGEMA_signal_6652, SubBytesIns_Inst_Sbox_10_T19}), .clk (clk), .r ({Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066]}), .c ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, new_AGEMA_signal_10252, SubBytesIns_Inst_Sbox_10_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M58_U1 ( .a ({new_AGEMA_signal_10233, new_AGEMA_signal_10232, new_AGEMA_signal_10231, SubBytesIns_Inst_Sbox_10_M43}), .b ({new_AGEMA_signal_6129, new_AGEMA_signal_6128, new_AGEMA_signal_6127, SubBytesIns_Inst_Sbox_10_T3}), .clk (clk), .r ({Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072]}), .c ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, new_AGEMA_signal_10963, SubBytesIns_Inst_Sbox_10_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M59_U1 ( .a ({new_AGEMA_signal_9654, new_AGEMA_signal_9653, new_AGEMA_signal_9652, SubBytesIns_Inst_Sbox_10_M38}), .b ({new_AGEMA_signal_6657, new_AGEMA_signal_6656, new_AGEMA_signal_6655, SubBytesIns_Inst_Sbox_10_T22}), .clk (clk), .r ({Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078]}), .c ({new_AGEMA_signal_10257, new_AGEMA_signal_10256, new_AGEMA_signal_10255, SubBytesIns_Inst_Sbox_10_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M60_U1 ( .a ({new_AGEMA_signal_9651, new_AGEMA_signal_9650, new_AGEMA_signal_9649, SubBytesIns_Inst_Sbox_10_M37}), .b ({new_AGEMA_signal_7341, new_AGEMA_signal_7340, new_AGEMA_signal_7339, SubBytesIns_Inst_Sbox_10_T20}), .clk (clk), .r ({Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084]}), .c ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, new_AGEMA_signal_10258, SubBytesIns_Inst_Sbox_10_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M61_U1 ( .a ({new_AGEMA_signal_10230, new_AGEMA_signal_10229, new_AGEMA_signal_10228, SubBytesIns_Inst_Sbox_10_M42}), .b ({new_AGEMA_signal_6123, new_AGEMA_signal_6122, new_AGEMA_signal_6121, SubBytesIns_Inst_Sbox_10_T1}), .clk (clk), .r ({Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090]}), .c ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M62_U1 ( .a ({new_AGEMA_signal_10947, new_AGEMA_signal_10946, new_AGEMA_signal_10945, SubBytesIns_Inst_Sbox_10_M45}), .b ({new_AGEMA_signal_6132, new_AGEMA_signal_6131, new_AGEMA_signal_6130, SubBytesIns_Inst_Sbox_10_T4}), .clk (clk), .r ({Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096]}), .c ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, new_AGEMA_signal_11584, SubBytesIns_Inst_Sbox_10_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_AND_M63_U1 ( .a ({new_AGEMA_signal_10227, new_AGEMA_signal_10226, new_AGEMA_signal_10225, SubBytesIns_Inst_Sbox_10_M41}), .b ({new_AGEMA_signal_6126, new_AGEMA_signal_6125, new_AGEMA_signal_6124, SubBytesIns_Inst_Sbox_10_T2}), .clk (clk), .r ({Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102]}), .c ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, new_AGEMA_signal_10969, SubBytesIns_Inst_Sbox_10_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L0_U1 ( .a ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}), .b ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, new_AGEMA_signal_11584, SubBytesIns_Inst_Sbox_10_M62}), .c ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L1_U1 ( .a ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, new_AGEMA_signal_10243, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, new_AGEMA_signal_10249, SubBytesIns_Inst_Sbox_10_M56}), .c ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L2_U1 ( .a ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, new_AGEMA_signal_10948, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, new_AGEMA_signal_10240, SubBytesIns_Inst_Sbox_10_M48}), .c ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, new_AGEMA_signal_11587, SubBytesIns_Inst_Sbox_10_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L3_U1 ( .a ({new_AGEMA_signal_10239, new_AGEMA_signal_10238, new_AGEMA_signal_10237, SubBytesIns_Inst_Sbox_10_M47}), .b ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, new_AGEMA_signal_10960, SubBytesIns_Inst_Sbox_10_M55}), .c ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, new_AGEMA_signal_11590, SubBytesIns_Inst_Sbox_10_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L4_U1 ( .a ({new_AGEMA_signal_10959, new_AGEMA_signal_10958, new_AGEMA_signal_10957, SubBytesIns_Inst_Sbox_10_M54}), .b ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, new_AGEMA_signal_10963, SubBytesIns_Inst_Sbox_10_M58}), .c ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, new_AGEMA_signal_11593, SubBytesIns_Inst_Sbox_10_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L5_U1 ( .a ({new_AGEMA_signal_10953, new_AGEMA_signal_10952, new_AGEMA_signal_10951, SubBytesIns_Inst_Sbox_10_M49}), .b ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, new_AGEMA_signal_11596, SubBytesIns_Inst_Sbox_10_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L6_U1 ( .a ({new_AGEMA_signal_11586, new_AGEMA_signal_11585, new_AGEMA_signal_11584, SubBytesIns_Inst_Sbox_10_M62}), .b ({new_AGEMA_signal_11598, new_AGEMA_signal_11597, new_AGEMA_signal_11596, SubBytesIns_Inst_Sbox_10_L5}), .c ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L7_U1 ( .a ({new_AGEMA_signal_10950, new_AGEMA_signal_10949, new_AGEMA_signal_10948, SubBytesIns_Inst_Sbox_10_M46}), .b ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, new_AGEMA_signal_11590, SubBytesIns_Inst_Sbox_10_L3}), .c ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, new_AGEMA_signal_12145, SubBytesIns_Inst_Sbox_10_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L8_U1 ( .a ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, new_AGEMA_signal_10246, SubBytesIns_Inst_Sbox_10_M51}), .b ({new_AGEMA_signal_10257, new_AGEMA_signal_10256, new_AGEMA_signal_10255, SubBytesIns_Inst_Sbox_10_M59}), .c ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, new_AGEMA_signal_10975, SubBytesIns_Inst_Sbox_10_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L9_U1 ( .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, new_AGEMA_signal_10954, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, new_AGEMA_signal_11581, SubBytesIns_Inst_Sbox_10_M53}), .c ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, new_AGEMA_signal_12148, SubBytesIns_Inst_Sbox_10_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L10_U1 ( .a ({new_AGEMA_signal_11583, new_AGEMA_signal_11582, new_AGEMA_signal_11581, SubBytesIns_Inst_Sbox_10_M53}), .b ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, new_AGEMA_signal_11593, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, new_AGEMA_signal_12151, SubBytesIns_Inst_Sbox_10_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L11_U1 ( .a ({new_AGEMA_signal_10260, new_AGEMA_signal_10259, new_AGEMA_signal_10258, SubBytesIns_Inst_Sbox_10_M60}), .b ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, new_AGEMA_signal_11587, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_12156, new_AGEMA_signal_12155, new_AGEMA_signal_12154, SubBytesIns_Inst_Sbox_10_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L12_U1 ( .a ({new_AGEMA_signal_10242, new_AGEMA_signal_10241, new_AGEMA_signal_10240, SubBytesIns_Inst_Sbox_10_M48}), .b ({new_AGEMA_signal_10248, new_AGEMA_signal_10247, new_AGEMA_signal_10246, SubBytesIns_Inst_Sbox_10_M51}), .c ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, new_AGEMA_signal_10978, SubBytesIns_Inst_Sbox_10_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L13_U1 ( .a ({new_AGEMA_signal_10245, new_AGEMA_signal_10244, new_AGEMA_signal_10243, SubBytesIns_Inst_Sbox_10_M50}), .b ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_12765, new_AGEMA_signal_12764, new_AGEMA_signal_12763, SubBytesIns_Inst_Sbox_10_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L14_U1 ( .a ({new_AGEMA_signal_10956, new_AGEMA_signal_10955, new_AGEMA_signal_10954, SubBytesIns_Inst_Sbox_10_M52}), .b ({new_AGEMA_signal_10968, new_AGEMA_signal_10967, new_AGEMA_signal_10966, SubBytesIns_Inst_Sbox_10_M61}), .c ({new_AGEMA_signal_11601, new_AGEMA_signal_11600, new_AGEMA_signal_11599, SubBytesIns_Inst_Sbox_10_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L15_U1 ( .a ({new_AGEMA_signal_10962, new_AGEMA_signal_10961, new_AGEMA_signal_10960, SubBytesIns_Inst_Sbox_10_M55}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, new_AGEMA_signal_11602, SubBytesIns_Inst_Sbox_10_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L16_U1 ( .a ({new_AGEMA_signal_10251, new_AGEMA_signal_10250, new_AGEMA_signal_10249, SubBytesIns_Inst_Sbox_10_M56}), .b ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}), .c ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, new_AGEMA_signal_12766, SubBytesIns_Inst_Sbox_10_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L17_U1 ( .a ({new_AGEMA_signal_10254, new_AGEMA_signal_10253, new_AGEMA_signal_10252, SubBytesIns_Inst_Sbox_10_M57}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_11607, new_AGEMA_signal_11606, new_AGEMA_signal_11605, SubBytesIns_Inst_Sbox_10_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L18_U1 ( .a ({new_AGEMA_signal_10965, new_AGEMA_signal_10964, new_AGEMA_signal_10963, SubBytesIns_Inst_Sbox_10_M58}), .b ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, new_AGEMA_signal_10975, SubBytesIns_Inst_Sbox_10_L8}), .c ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, new_AGEMA_signal_11608, SubBytesIns_Inst_Sbox_10_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L19_U1 ( .a ({new_AGEMA_signal_10971, new_AGEMA_signal_10970, new_AGEMA_signal_10969, SubBytesIns_Inst_Sbox_10_M63}), .b ({new_AGEMA_signal_11595, new_AGEMA_signal_11594, new_AGEMA_signal_11593, SubBytesIns_Inst_Sbox_10_L4}), .c ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, new_AGEMA_signal_12157, SubBytesIns_Inst_Sbox_10_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L20_U1 ( .a ({new_AGEMA_signal_12141, new_AGEMA_signal_12140, new_AGEMA_signal_12139, SubBytesIns_Inst_Sbox_10_L0}), .b ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .c ({new_AGEMA_signal_12771, new_AGEMA_signal_12770, new_AGEMA_signal_12769, SubBytesIns_Inst_Sbox_10_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L21_U1 ( .a ({new_AGEMA_signal_10974, new_AGEMA_signal_10973, new_AGEMA_signal_10972, SubBytesIns_Inst_Sbox_10_L1}), .b ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, new_AGEMA_signal_12145, SubBytesIns_Inst_Sbox_10_L7}), .c ({new_AGEMA_signal_12774, new_AGEMA_signal_12773, new_AGEMA_signal_12772, SubBytesIns_Inst_Sbox_10_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L22_U1 ( .a ({new_AGEMA_signal_11592, new_AGEMA_signal_11591, new_AGEMA_signal_11590, SubBytesIns_Inst_Sbox_10_L3}), .b ({new_AGEMA_signal_10980, new_AGEMA_signal_10979, new_AGEMA_signal_10978, SubBytesIns_Inst_Sbox_10_L12}), .c ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, new_AGEMA_signal_12160, SubBytesIns_Inst_Sbox_10_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L23_U1 ( .a ({new_AGEMA_signal_11610, new_AGEMA_signal_11609, new_AGEMA_signal_11608, SubBytesIns_Inst_Sbox_10_L18}), .b ({new_AGEMA_signal_11589, new_AGEMA_signal_11588, new_AGEMA_signal_11587, SubBytesIns_Inst_Sbox_10_L2}), .c ({new_AGEMA_signal_12165, new_AGEMA_signal_12164, new_AGEMA_signal_12163, SubBytesIns_Inst_Sbox_10_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L24_U1 ( .a ({new_AGEMA_signal_11604, new_AGEMA_signal_11603, new_AGEMA_signal_11602, SubBytesIns_Inst_Sbox_10_L15}), .b ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, new_AGEMA_signal_12148, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_12777, new_AGEMA_signal_12776, new_AGEMA_signal_12775, SubBytesIns_Inst_Sbox_10_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L25_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, new_AGEMA_signal_12151, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, new_AGEMA_signal_12778, SubBytesIns_Inst_Sbox_10_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L26_U1 ( .a ({new_AGEMA_signal_12147, new_AGEMA_signal_12146, new_AGEMA_signal_12145, SubBytesIns_Inst_Sbox_10_L7}), .b ({new_AGEMA_signal_12150, new_AGEMA_signal_12149, new_AGEMA_signal_12148, SubBytesIns_Inst_Sbox_10_L9}), .c ({new_AGEMA_signal_12783, new_AGEMA_signal_12782, new_AGEMA_signal_12781, SubBytesIns_Inst_Sbox_10_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L27_U1 ( .a ({new_AGEMA_signal_10977, new_AGEMA_signal_10976, new_AGEMA_signal_10975, SubBytesIns_Inst_Sbox_10_L8}), .b ({new_AGEMA_signal_12153, new_AGEMA_signal_12152, new_AGEMA_signal_12151, SubBytesIns_Inst_Sbox_10_L10}), .c ({new_AGEMA_signal_12786, new_AGEMA_signal_12785, new_AGEMA_signal_12784, SubBytesIns_Inst_Sbox_10_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L28_U1 ( .a ({new_AGEMA_signal_12156, new_AGEMA_signal_12155, new_AGEMA_signal_12154, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_11601, new_AGEMA_signal_11600, new_AGEMA_signal_11599, SubBytesIns_Inst_Sbox_10_L14}), .c ({new_AGEMA_signal_12789, new_AGEMA_signal_12788, new_AGEMA_signal_12787, SubBytesIns_Inst_Sbox_10_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_L29_U1 ( .a ({new_AGEMA_signal_12156, new_AGEMA_signal_12155, new_AGEMA_signal_12154, SubBytesIns_Inst_Sbox_10_L11}), .b ({new_AGEMA_signal_11607, new_AGEMA_signal_11606, new_AGEMA_signal_11605, SubBytesIns_Inst_Sbox_10_L17}), .c ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, new_AGEMA_signal_12790, SubBytesIns_Inst_Sbox_10_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S0_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12777, new_AGEMA_signal_12776, new_AGEMA_signal_12775, SubBytesIns_Inst_Sbox_10_L24}), .c ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S1_U1 ( .a ({new_AGEMA_signal_12768, new_AGEMA_signal_12767, new_AGEMA_signal_12766, SubBytesIns_Inst_Sbox_10_L16}), .b ({new_AGEMA_signal_12783, new_AGEMA_signal_12782, new_AGEMA_signal_12781, SubBytesIns_Inst_Sbox_10_L26}), .c ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S2_U1 ( .a ({new_AGEMA_signal_12159, new_AGEMA_signal_12158, new_AGEMA_signal_12157, SubBytesIns_Inst_Sbox_10_L19}), .b ({new_AGEMA_signal_12789, new_AGEMA_signal_12788, new_AGEMA_signal_12787, SubBytesIns_Inst_Sbox_10_L28}), .c ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S3_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12774, new_AGEMA_signal_12773, new_AGEMA_signal_12772, SubBytesIns_Inst_Sbox_10_L21}), .c ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S4_U1 ( .a ({new_AGEMA_signal_12771, new_AGEMA_signal_12770, new_AGEMA_signal_12769, SubBytesIns_Inst_Sbox_10_L20}), .b ({new_AGEMA_signal_12162, new_AGEMA_signal_12161, new_AGEMA_signal_12160, SubBytesIns_Inst_Sbox_10_L22}), .c ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S5_U1 ( .a ({new_AGEMA_signal_12780, new_AGEMA_signal_12779, new_AGEMA_signal_12778, SubBytesIns_Inst_Sbox_10_L25}), .b ({new_AGEMA_signal_12792, new_AGEMA_signal_12791, new_AGEMA_signal_12790, SubBytesIns_Inst_Sbox_10_L29}), .c ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S6_U1 ( .a ({new_AGEMA_signal_12765, new_AGEMA_signal_12764, new_AGEMA_signal_12763, SubBytesIns_Inst_Sbox_10_L13}), .b ({new_AGEMA_signal_12786, new_AGEMA_signal_12785, new_AGEMA_signal_12784, SubBytesIns_Inst_Sbox_10_L27}), .c ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_10_XOR_S7_U1 ( .a ({new_AGEMA_signal_12144, new_AGEMA_signal_12143, new_AGEMA_signal_12142, SubBytesIns_Inst_Sbox_10_L6}), .b ({new_AGEMA_signal_12165, new_AGEMA_signal_12164, new_AGEMA_signal_12163, SubBytesIns_Inst_Sbox_10_L23}), .c ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M46_U1 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, new_AGEMA_signal_10270, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_6663, new_AGEMA_signal_6662, new_AGEMA_signal_6661, SubBytesIns_Inst_Sbox_11_T6}), .clk (clk), .r ({Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108]}), .c ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, new_AGEMA_signal_10984, SubBytesIns_Inst_Sbox_11_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M47_U1 ( .a ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_7368, new_AGEMA_signal_7367, new_AGEMA_signal_7366, SubBytesIns_Inst_Sbox_11_T8}), .clk (clk), .r ({Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114]}), .c ({new_AGEMA_signal_10275, new_AGEMA_signal_10274, new_AGEMA_signal_10273, SubBytesIns_Inst_Sbox_11_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M48_U1 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .b ({ciphertext_s3[88], ciphertext_s2[88], ciphertext_s1[88], ciphertext_s0[88]}), .clk (clk), .r ({Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120]}), .c ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, new_AGEMA_signal_10276, SubBytesIns_Inst_Sbox_11_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M49_U1 ( .a ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, new_AGEMA_signal_10267, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_6675, new_AGEMA_signal_6674, new_AGEMA_signal_6673, SubBytesIns_Inst_Sbox_11_T16}), .clk (clk), .r ({Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126]}), .c ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, new_AGEMA_signal_10987, SubBytesIns_Inst_Sbox_11_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M50_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_6666, new_AGEMA_signal_6665, new_AGEMA_signal_6664, SubBytesIns_Inst_Sbox_11_T9}), .clk (clk), .r ({Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132]}), .c ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, new_AGEMA_signal_10279, SubBytesIns_Inst_Sbox_11_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M51_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_7377, new_AGEMA_signal_7376, new_AGEMA_signal_7375, SubBytesIns_Inst_Sbox_11_T17}), .clk (clk), .r ({Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138]}), .c ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, new_AGEMA_signal_10282, SubBytesIns_Inst_Sbox_11_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M52_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_6672, new_AGEMA_signal_6671, new_AGEMA_signal_6670, SubBytesIns_Inst_Sbox_11_T15}), .clk (clk), .r ({Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144]}), .c ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, new_AGEMA_signal_10990, SubBytesIns_Inst_Sbox_11_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M53_U1 ( .a ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, new_AGEMA_signal_10981, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_6684, new_AGEMA_signal_6683, new_AGEMA_signal_6682, SubBytesIns_Inst_Sbox_11_T27}), .clk (clk), .r ({Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150]}), .c ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, new_AGEMA_signal_11611, SubBytesIns_Inst_Sbox_11_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M54_U1 ( .a ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_7371, new_AGEMA_signal_7370, new_AGEMA_signal_7369, SubBytesIns_Inst_Sbox_11_T10}), .clk (clk), .r ({Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156]}), .c ({new_AGEMA_signal_10995, new_AGEMA_signal_10994, new_AGEMA_signal_10993, SubBytesIns_Inst_Sbox_11_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M55_U1 ( .a ({new_AGEMA_signal_10272, new_AGEMA_signal_10271, new_AGEMA_signal_10270, SubBytesIns_Inst_Sbox_11_M44}), .b ({new_AGEMA_signal_6669, new_AGEMA_signal_6668, new_AGEMA_signal_6667, SubBytesIns_Inst_Sbox_11_T13}), .clk (clk), .r ({Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162]}), .c ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, new_AGEMA_signal_10996, SubBytesIns_Inst_Sbox_11_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M56_U1 ( .a ({new_AGEMA_signal_9672, new_AGEMA_signal_9671, new_AGEMA_signal_9670, SubBytesIns_Inst_Sbox_11_M40}), .b ({new_AGEMA_signal_7383, new_AGEMA_signal_7382, new_AGEMA_signal_7381, SubBytesIns_Inst_Sbox_11_T23}), .clk (clk), .r ({Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168]}), .c ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, new_AGEMA_signal_10285, SubBytesIns_Inst_Sbox_11_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M57_U1 ( .a ({new_AGEMA_signal_9669, new_AGEMA_signal_9668, new_AGEMA_signal_9667, SubBytesIns_Inst_Sbox_11_M39}), .b ({new_AGEMA_signal_6678, new_AGEMA_signal_6677, new_AGEMA_signal_6676, SubBytesIns_Inst_Sbox_11_T19}), .clk (clk), .r ({Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174]}), .c ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, new_AGEMA_signal_10288, SubBytesIns_Inst_Sbox_11_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M58_U1 ( .a ({new_AGEMA_signal_10269, new_AGEMA_signal_10268, new_AGEMA_signal_10267, SubBytesIns_Inst_Sbox_11_M43}), .b ({new_AGEMA_signal_6159, new_AGEMA_signal_6158, new_AGEMA_signal_6157, SubBytesIns_Inst_Sbox_11_T3}), .clk (clk), .r ({Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180]}), .c ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, new_AGEMA_signal_10999, SubBytesIns_Inst_Sbox_11_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M59_U1 ( .a ({new_AGEMA_signal_9666, new_AGEMA_signal_9665, new_AGEMA_signal_9664, SubBytesIns_Inst_Sbox_11_M38}), .b ({new_AGEMA_signal_6681, new_AGEMA_signal_6680, new_AGEMA_signal_6679, SubBytesIns_Inst_Sbox_11_T22}), .clk (clk), .r ({Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186]}), .c ({new_AGEMA_signal_10293, new_AGEMA_signal_10292, new_AGEMA_signal_10291, SubBytesIns_Inst_Sbox_11_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M60_U1 ( .a ({new_AGEMA_signal_9663, new_AGEMA_signal_9662, new_AGEMA_signal_9661, SubBytesIns_Inst_Sbox_11_M37}), .b ({new_AGEMA_signal_7380, new_AGEMA_signal_7379, new_AGEMA_signal_7378, SubBytesIns_Inst_Sbox_11_T20}), .clk (clk), .r ({Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192]}), .c ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, new_AGEMA_signal_10294, SubBytesIns_Inst_Sbox_11_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M61_U1 ( .a ({new_AGEMA_signal_10266, new_AGEMA_signal_10265, new_AGEMA_signal_10264, SubBytesIns_Inst_Sbox_11_M42}), .b ({new_AGEMA_signal_6153, new_AGEMA_signal_6152, new_AGEMA_signal_6151, SubBytesIns_Inst_Sbox_11_T1}), .clk (clk), .r ({Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198]}), .c ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M62_U1 ( .a ({new_AGEMA_signal_10983, new_AGEMA_signal_10982, new_AGEMA_signal_10981, SubBytesIns_Inst_Sbox_11_M45}), .b ({new_AGEMA_signal_6162, new_AGEMA_signal_6161, new_AGEMA_signal_6160, SubBytesIns_Inst_Sbox_11_T4}), .clk (clk), .r ({Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204]}), .c ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, new_AGEMA_signal_11614, SubBytesIns_Inst_Sbox_11_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_AND_M63_U1 ( .a ({new_AGEMA_signal_10263, new_AGEMA_signal_10262, new_AGEMA_signal_10261, SubBytesIns_Inst_Sbox_11_M41}), .b ({new_AGEMA_signal_6156, new_AGEMA_signal_6155, new_AGEMA_signal_6154, SubBytesIns_Inst_Sbox_11_T2}), .clk (clk), .r ({Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210]}), .c ({new_AGEMA_signal_11007, new_AGEMA_signal_11006, new_AGEMA_signal_11005, SubBytesIns_Inst_Sbox_11_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L0_U1 ( .a ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}), .b ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, new_AGEMA_signal_11614, SubBytesIns_Inst_Sbox_11_M62}), .c ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L1_U1 ( .a ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, new_AGEMA_signal_10279, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, new_AGEMA_signal_10285, SubBytesIns_Inst_Sbox_11_M56}), .c ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L2_U1 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, new_AGEMA_signal_10984, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, new_AGEMA_signal_10276, SubBytesIns_Inst_Sbox_11_M48}), .c ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, new_AGEMA_signal_11617, SubBytesIns_Inst_Sbox_11_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L3_U1 ( .a ({new_AGEMA_signal_10275, new_AGEMA_signal_10274, new_AGEMA_signal_10273, SubBytesIns_Inst_Sbox_11_M47}), .b ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, new_AGEMA_signal_10996, SubBytesIns_Inst_Sbox_11_M55}), .c ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, new_AGEMA_signal_11620, SubBytesIns_Inst_Sbox_11_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L4_U1 ( .a ({new_AGEMA_signal_10995, new_AGEMA_signal_10994, new_AGEMA_signal_10993, SubBytesIns_Inst_Sbox_11_M54}), .b ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, new_AGEMA_signal_10999, SubBytesIns_Inst_Sbox_11_M58}), .c ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, new_AGEMA_signal_11623, SubBytesIns_Inst_Sbox_11_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L5_U1 ( .a ({new_AGEMA_signal_10989, new_AGEMA_signal_10988, new_AGEMA_signal_10987, SubBytesIns_Inst_Sbox_11_M49}), .b ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, new_AGEMA_signal_11626, SubBytesIns_Inst_Sbox_11_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L6_U1 ( .a ({new_AGEMA_signal_11616, new_AGEMA_signal_11615, new_AGEMA_signal_11614, SubBytesIns_Inst_Sbox_11_M62}), .b ({new_AGEMA_signal_11628, new_AGEMA_signal_11627, new_AGEMA_signal_11626, SubBytesIns_Inst_Sbox_11_L5}), .c ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L7_U1 ( .a ({new_AGEMA_signal_10986, new_AGEMA_signal_10985, new_AGEMA_signal_10984, SubBytesIns_Inst_Sbox_11_M46}), .b ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, new_AGEMA_signal_11620, SubBytesIns_Inst_Sbox_11_L3}), .c ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, new_AGEMA_signal_12172, SubBytesIns_Inst_Sbox_11_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L8_U1 ( .a ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, new_AGEMA_signal_10282, SubBytesIns_Inst_Sbox_11_M51}), .b ({new_AGEMA_signal_10293, new_AGEMA_signal_10292, new_AGEMA_signal_10291, SubBytesIns_Inst_Sbox_11_M59}), .c ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, new_AGEMA_signal_11011, SubBytesIns_Inst_Sbox_11_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L9_U1 ( .a ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, new_AGEMA_signal_10990, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, new_AGEMA_signal_11611, SubBytesIns_Inst_Sbox_11_M53}), .c ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, new_AGEMA_signal_12175, SubBytesIns_Inst_Sbox_11_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L10_U1 ( .a ({new_AGEMA_signal_11613, new_AGEMA_signal_11612, new_AGEMA_signal_11611, SubBytesIns_Inst_Sbox_11_M53}), .b ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, new_AGEMA_signal_11623, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_12180, new_AGEMA_signal_12179, new_AGEMA_signal_12178, SubBytesIns_Inst_Sbox_11_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L11_U1 ( .a ({new_AGEMA_signal_10296, new_AGEMA_signal_10295, new_AGEMA_signal_10294, SubBytesIns_Inst_Sbox_11_M60}), .b ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, new_AGEMA_signal_11617, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, new_AGEMA_signal_12181, SubBytesIns_Inst_Sbox_11_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L12_U1 ( .a ({new_AGEMA_signal_10278, new_AGEMA_signal_10277, new_AGEMA_signal_10276, SubBytesIns_Inst_Sbox_11_M48}), .b ({new_AGEMA_signal_10284, new_AGEMA_signal_10283, new_AGEMA_signal_10282, SubBytesIns_Inst_Sbox_11_M51}), .c ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, new_AGEMA_signal_11014, SubBytesIns_Inst_Sbox_11_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L13_U1 ( .a ({new_AGEMA_signal_10281, new_AGEMA_signal_10280, new_AGEMA_signal_10279, SubBytesIns_Inst_Sbox_11_M50}), .b ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_12798, new_AGEMA_signal_12797, new_AGEMA_signal_12796, SubBytesIns_Inst_Sbox_11_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L14_U1 ( .a ({new_AGEMA_signal_10992, new_AGEMA_signal_10991, new_AGEMA_signal_10990, SubBytesIns_Inst_Sbox_11_M52}), .b ({new_AGEMA_signal_11004, new_AGEMA_signal_11003, new_AGEMA_signal_11002, SubBytesIns_Inst_Sbox_11_M61}), .c ({new_AGEMA_signal_11631, new_AGEMA_signal_11630, new_AGEMA_signal_11629, SubBytesIns_Inst_Sbox_11_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L15_U1 ( .a ({new_AGEMA_signal_10998, new_AGEMA_signal_10997, new_AGEMA_signal_10996, SubBytesIns_Inst_Sbox_11_M55}), .b ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, new_AGEMA_signal_11632, SubBytesIns_Inst_Sbox_11_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L16_U1 ( .a ({new_AGEMA_signal_10287, new_AGEMA_signal_10286, new_AGEMA_signal_10285, SubBytesIns_Inst_Sbox_11_M56}), .b ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}), .c ({new_AGEMA_signal_12801, new_AGEMA_signal_12800, new_AGEMA_signal_12799, SubBytesIns_Inst_Sbox_11_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L17_U1 ( .a ({new_AGEMA_signal_10290, new_AGEMA_signal_10289, new_AGEMA_signal_10288, SubBytesIns_Inst_Sbox_11_M57}), .b ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_11637, new_AGEMA_signal_11636, new_AGEMA_signal_11635, SubBytesIns_Inst_Sbox_11_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L18_U1 ( .a ({new_AGEMA_signal_11001, new_AGEMA_signal_11000, new_AGEMA_signal_10999, SubBytesIns_Inst_Sbox_11_M58}), .b ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, new_AGEMA_signal_11011, SubBytesIns_Inst_Sbox_11_L8}), .c ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, new_AGEMA_signal_11638, SubBytesIns_Inst_Sbox_11_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L19_U1 ( .a ({new_AGEMA_signal_11007, new_AGEMA_signal_11006, new_AGEMA_signal_11005, SubBytesIns_Inst_Sbox_11_M63}), .b ({new_AGEMA_signal_11625, new_AGEMA_signal_11624, new_AGEMA_signal_11623, SubBytesIns_Inst_Sbox_11_L4}), .c ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, new_AGEMA_signal_12184, SubBytesIns_Inst_Sbox_11_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L20_U1 ( .a ({new_AGEMA_signal_12168, new_AGEMA_signal_12167, new_AGEMA_signal_12166, SubBytesIns_Inst_Sbox_11_L0}), .b ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .c ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, new_AGEMA_signal_12802, SubBytesIns_Inst_Sbox_11_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L21_U1 ( .a ({new_AGEMA_signal_11010, new_AGEMA_signal_11009, new_AGEMA_signal_11008, SubBytesIns_Inst_Sbox_11_L1}), .b ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, new_AGEMA_signal_12172, SubBytesIns_Inst_Sbox_11_L7}), .c ({new_AGEMA_signal_12807, new_AGEMA_signal_12806, new_AGEMA_signal_12805, SubBytesIns_Inst_Sbox_11_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L22_U1 ( .a ({new_AGEMA_signal_11622, new_AGEMA_signal_11621, new_AGEMA_signal_11620, SubBytesIns_Inst_Sbox_11_L3}), .b ({new_AGEMA_signal_11016, new_AGEMA_signal_11015, new_AGEMA_signal_11014, SubBytesIns_Inst_Sbox_11_L12}), .c ({new_AGEMA_signal_12189, new_AGEMA_signal_12188, new_AGEMA_signal_12187, SubBytesIns_Inst_Sbox_11_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L23_U1 ( .a ({new_AGEMA_signal_11640, new_AGEMA_signal_11639, new_AGEMA_signal_11638, SubBytesIns_Inst_Sbox_11_L18}), .b ({new_AGEMA_signal_11619, new_AGEMA_signal_11618, new_AGEMA_signal_11617, SubBytesIns_Inst_Sbox_11_L2}), .c ({new_AGEMA_signal_12192, new_AGEMA_signal_12191, new_AGEMA_signal_12190, SubBytesIns_Inst_Sbox_11_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L24_U1 ( .a ({new_AGEMA_signal_11634, new_AGEMA_signal_11633, new_AGEMA_signal_11632, SubBytesIns_Inst_Sbox_11_L15}), .b ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, new_AGEMA_signal_12175, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_12810, new_AGEMA_signal_12809, new_AGEMA_signal_12808, SubBytesIns_Inst_Sbox_11_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L25_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12180, new_AGEMA_signal_12179, new_AGEMA_signal_12178, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_12813, new_AGEMA_signal_12812, new_AGEMA_signal_12811, SubBytesIns_Inst_Sbox_11_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L26_U1 ( .a ({new_AGEMA_signal_12174, new_AGEMA_signal_12173, new_AGEMA_signal_12172, SubBytesIns_Inst_Sbox_11_L7}), .b ({new_AGEMA_signal_12177, new_AGEMA_signal_12176, new_AGEMA_signal_12175, SubBytesIns_Inst_Sbox_11_L9}), .c ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, new_AGEMA_signal_12814, SubBytesIns_Inst_Sbox_11_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L27_U1 ( .a ({new_AGEMA_signal_11013, new_AGEMA_signal_11012, new_AGEMA_signal_11011, SubBytesIns_Inst_Sbox_11_L8}), .b ({new_AGEMA_signal_12180, new_AGEMA_signal_12179, new_AGEMA_signal_12178, SubBytesIns_Inst_Sbox_11_L10}), .c ({new_AGEMA_signal_12819, new_AGEMA_signal_12818, new_AGEMA_signal_12817, SubBytesIns_Inst_Sbox_11_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L28_U1 ( .a ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, new_AGEMA_signal_12181, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_11631, new_AGEMA_signal_11630, new_AGEMA_signal_11629, SubBytesIns_Inst_Sbox_11_L14}), .c ({new_AGEMA_signal_12822, new_AGEMA_signal_12821, new_AGEMA_signal_12820, SubBytesIns_Inst_Sbox_11_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_L29_U1 ( .a ({new_AGEMA_signal_12183, new_AGEMA_signal_12182, new_AGEMA_signal_12181, SubBytesIns_Inst_Sbox_11_L11}), .b ({new_AGEMA_signal_11637, new_AGEMA_signal_11636, new_AGEMA_signal_11635, SubBytesIns_Inst_Sbox_11_L17}), .c ({new_AGEMA_signal_12825, new_AGEMA_signal_12824, new_AGEMA_signal_12823, SubBytesIns_Inst_Sbox_11_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S0_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12810, new_AGEMA_signal_12809, new_AGEMA_signal_12808, SubBytesIns_Inst_Sbox_11_L24}), .c ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S1_U1 ( .a ({new_AGEMA_signal_12801, new_AGEMA_signal_12800, new_AGEMA_signal_12799, SubBytesIns_Inst_Sbox_11_L16}), .b ({new_AGEMA_signal_12816, new_AGEMA_signal_12815, new_AGEMA_signal_12814, SubBytesIns_Inst_Sbox_11_L26}), .c ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S2_U1 ( .a ({new_AGEMA_signal_12186, new_AGEMA_signal_12185, new_AGEMA_signal_12184, SubBytesIns_Inst_Sbox_11_L19}), .b ({new_AGEMA_signal_12822, new_AGEMA_signal_12821, new_AGEMA_signal_12820, SubBytesIns_Inst_Sbox_11_L28}), .c ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S3_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12807, new_AGEMA_signal_12806, new_AGEMA_signal_12805, SubBytesIns_Inst_Sbox_11_L21}), .c ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S4_U1 ( .a ({new_AGEMA_signal_12804, new_AGEMA_signal_12803, new_AGEMA_signal_12802, SubBytesIns_Inst_Sbox_11_L20}), .b ({new_AGEMA_signal_12189, new_AGEMA_signal_12188, new_AGEMA_signal_12187, SubBytesIns_Inst_Sbox_11_L22}), .c ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S5_U1 ( .a ({new_AGEMA_signal_12813, new_AGEMA_signal_12812, new_AGEMA_signal_12811, SubBytesIns_Inst_Sbox_11_L25}), .b ({new_AGEMA_signal_12825, new_AGEMA_signal_12824, new_AGEMA_signal_12823, SubBytesIns_Inst_Sbox_11_L29}), .c ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S6_U1 ( .a ({new_AGEMA_signal_12798, new_AGEMA_signal_12797, new_AGEMA_signal_12796, SubBytesIns_Inst_Sbox_11_L13}), .b ({new_AGEMA_signal_12819, new_AGEMA_signal_12818, new_AGEMA_signal_12817, SubBytesIns_Inst_Sbox_11_L27}), .c ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_11_XOR_S7_U1 ( .a ({new_AGEMA_signal_12171, new_AGEMA_signal_12170, new_AGEMA_signal_12169, SubBytesIns_Inst_Sbox_11_L6}), .b ({new_AGEMA_signal_12192, new_AGEMA_signal_12191, new_AGEMA_signal_12190, SubBytesIns_Inst_Sbox_11_L23}), .c ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M46_U1 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, new_AGEMA_signal_10306, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_6687, new_AGEMA_signal_6686, new_AGEMA_signal_6685, SubBytesIns_Inst_Sbox_12_T6}), .clk (clk), .r ({Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216]}), .c ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, new_AGEMA_signal_11020, SubBytesIns_Inst_Sbox_12_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M47_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_7407, new_AGEMA_signal_7406, new_AGEMA_signal_7405, SubBytesIns_Inst_Sbox_12_T8}), .clk (clk), .r ({Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222]}), .c ({new_AGEMA_signal_10311, new_AGEMA_signal_10310, new_AGEMA_signal_10309, SubBytesIns_Inst_Sbox_12_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M48_U1 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .b ({ciphertext_s3[96], ciphertext_s2[96], ciphertext_s1[96], ciphertext_s0[96]}), .clk (clk), .r ({Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228]}), .c ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, new_AGEMA_signal_10312, SubBytesIns_Inst_Sbox_12_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M49_U1 ( .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, new_AGEMA_signal_10303, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_6699, new_AGEMA_signal_6698, new_AGEMA_signal_6697, SubBytesIns_Inst_Sbox_12_T16}), .clk (clk), .r ({Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234]}), .c ({new_AGEMA_signal_11025, new_AGEMA_signal_11024, new_AGEMA_signal_11023, SubBytesIns_Inst_Sbox_12_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M50_U1 ( .a ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_6690, new_AGEMA_signal_6689, new_AGEMA_signal_6688, SubBytesIns_Inst_Sbox_12_T9}), .clk (clk), .r ({Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240]}), .c ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, new_AGEMA_signal_10315, SubBytesIns_Inst_Sbox_12_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M51_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_7416, new_AGEMA_signal_7415, new_AGEMA_signal_7414, SubBytesIns_Inst_Sbox_12_T17}), .clk (clk), .r ({Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246]}), .c ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, new_AGEMA_signal_10318, SubBytesIns_Inst_Sbox_12_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M52_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_6696, new_AGEMA_signal_6695, new_AGEMA_signal_6694, SubBytesIns_Inst_Sbox_12_T15}), .clk (clk), .r ({Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252]}), .c ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, new_AGEMA_signal_11026, SubBytesIns_Inst_Sbox_12_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M53_U1 ( .a ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, new_AGEMA_signal_11017, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_6708, new_AGEMA_signal_6707, new_AGEMA_signal_6706, SubBytesIns_Inst_Sbox_12_T27}), .clk (clk), .r ({Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258]}), .c ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, new_AGEMA_signal_11641, SubBytesIns_Inst_Sbox_12_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M54_U1 ( .a ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_7410, new_AGEMA_signal_7409, new_AGEMA_signal_7408, SubBytesIns_Inst_Sbox_12_T10}), .clk (clk), .r ({Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264]}), .c ({new_AGEMA_signal_11031, new_AGEMA_signal_11030, new_AGEMA_signal_11029, SubBytesIns_Inst_Sbox_12_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M55_U1 ( .a ({new_AGEMA_signal_10308, new_AGEMA_signal_10307, new_AGEMA_signal_10306, SubBytesIns_Inst_Sbox_12_M44}), .b ({new_AGEMA_signal_6693, new_AGEMA_signal_6692, new_AGEMA_signal_6691, SubBytesIns_Inst_Sbox_12_T13}), .clk (clk), .r ({Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270]}), .c ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, new_AGEMA_signal_11032, SubBytesIns_Inst_Sbox_12_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M56_U1 ( .a ({new_AGEMA_signal_9684, new_AGEMA_signal_9683, new_AGEMA_signal_9682, SubBytesIns_Inst_Sbox_12_M40}), .b ({new_AGEMA_signal_7422, new_AGEMA_signal_7421, new_AGEMA_signal_7420, SubBytesIns_Inst_Sbox_12_T23}), .clk (clk), .r ({Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276]}), .c ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, new_AGEMA_signal_10321, SubBytesIns_Inst_Sbox_12_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M57_U1 ( .a ({new_AGEMA_signal_9681, new_AGEMA_signal_9680, new_AGEMA_signal_9679, SubBytesIns_Inst_Sbox_12_M39}), .b ({new_AGEMA_signal_6702, new_AGEMA_signal_6701, new_AGEMA_signal_6700, SubBytesIns_Inst_Sbox_12_T19}), .clk (clk), .r ({Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282]}), .c ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, new_AGEMA_signal_10324, SubBytesIns_Inst_Sbox_12_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M58_U1 ( .a ({new_AGEMA_signal_10305, new_AGEMA_signal_10304, new_AGEMA_signal_10303, SubBytesIns_Inst_Sbox_12_M43}), .b ({new_AGEMA_signal_6189, new_AGEMA_signal_6188, new_AGEMA_signal_6187, SubBytesIns_Inst_Sbox_12_T3}), .clk (clk), .r ({Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288]}), .c ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, new_AGEMA_signal_11035, SubBytesIns_Inst_Sbox_12_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M59_U1 ( .a ({new_AGEMA_signal_9678, new_AGEMA_signal_9677, new_AGEMA_signal_9676, SubBytesIns_Inst_Sbox_12_M38}), .b ({new_AGEMA_signal_6705, new_AGEMA_signal_6704, new_AGEMA_signal_6703, SubBytesIns_Inst_Sbox_12_T22}), .clk (clk), .r ({Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294]}), .c ({new_AGEMA_signal_10329, new_AGEMA_signal_10328, new_AGEMA_signal_10327, SubBytesIns_Inst_Sbox_12_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M60_U1 ( .a ({new_AGEMA_signal_9675, new_AGEMA_signal_9674, new_AGEMA_signal_9673, SubBytesIns_Inst_Sbox_12_M37}), .b ({new_AGEMA_signal_7419, new_AGEMA_signal_7418, new_AGEMA_signal_7417, SubBytesIns_Inst_Sbox_12_T20}), .clk (clk), .r ({Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300]}), .c ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, new_AGEMA_signal_10330, SubBytesIns_Inst_Sbox_12_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M61_U1 ( .a ({new_AGEMA_signal_10302, new_AGEMA_signal_10301, new_AGEMA_signal_10300, SubBytesIns_Inst_Sbox_12_M42}), .b ({new_AGEMA_signal_6183, new_AGEMA_signal_6182, new_AGEMA_signal_6181, SubBytesIns_Inst_Sbox_12_T1}), .clk (clk), .r ({Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306]}), .c ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M62_U1 ( .a ({new_AGEMA_signal_11019, new_AGEMA_signal_11018, new_AGEMA_signal_11017, SubBytesIns_Inst_Sbox_12_M45}), .b ({new_AGEMA_signal_6192, new_AGEMA_signal_6191, new_AGEMA_signal_6190, SubBytesIns_Inst_Sbox_12_T4}), .clk (clk), .r ({Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312]}), .c ({new_AGEMA_signal_11646, new_AGEMA_signal_11645, new_AGEMA_signal_11644, SubBytesIns_Inst_Sbox_12_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_AND_M63_U1 ( .a ({new_AGEMA_signal_10299, new_AGEMA_signal_10298, new_AGEMA_signal_10297, SubBytesIns_Inst_Sbox_12_M41}), .b ({new_AGEMA_signal_6186, new_AGEMA_signal_6185, new_AGEMA_signal_6184, SubBytesIns_Inst_Sbox_12_T2}), .clk (clk), .r ({Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318]}), .c ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, new_AGEMA_signal_11041, SubBytesIns_Inst_Sbox_12_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L0_U1 ( .a ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}), .b ({new_AGEMA_signal_11646, new_AGEMA_signal_11645, new_AGEMA_signal_11644, SubBytesIns_Inst_Sbox_12_M62}), .c ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L1_U1 ( .a ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, new_AGEMA_signal_10315, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, new_AGEMA_signal_10321, SubBytesIns_Inst_Sbox_12_M56}), .c ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L2_U1 ( .a ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, new_AGEMA_signal_11020, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, new_AGEMA_signal_10312, SubBytesIns_Inst_Sbox_12_M48}), .c ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, new_AGEMA_signal_11647, SubBytesIns_Inst_Sbox_12_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L3_U1 ( .a ({new_AGEMA_signal_10311, new_AGEMA_signal_10310, new_AGEMA_signal_10309, SubBytesIns_Inst_Sbox_12_M47}), .b ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, new_AGEMA_signal_11032, SubBytesIns_Inst_Sbox_12_M55}), .c ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, new_AGEMA_signal_11650, SubBytesIns_Inst_Sbox_12_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L4_U1 ( .a ({new_AGEMA_signal_11031, new_AGEMA_signal_11030, new_AGEMA_signal_11029, SubBytesIns_Inst_Sbox_12_M54}), .b ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, new_AGEMA_signal_11035, SubBytesIns_Inst_Sbox_12_M58}), .c ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, new_AGEMA_signal_11653, SubBytesIns_Inst_Sbox_12_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L5_U1 ( .a ({new_AGEMA_signal_11025, new_AGEMA_signal_11024, new_AGEMA_signal_11023, SubBytesIns_Inst_Sbox_12_M49}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_11658, new_AGEMA_signal_11657, new_AGEMA_signal_11656, SubBytesIns_Inst_Sbox_12_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L6_U1 ( .a ({new_AGEMA_signal_11646, new_AGEMA_signal_11645, new_AGEMA_signal_11644, SubBytesIns_Inst_Sbox_12_M62}), .b ({new_AGEMA_signal_11658, new_AGEMA_signal_11657, new_AGEMA_signal_11656, SubBytesIns_Inst_Sbox_12_L5}), .c ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L7_U1 ( .a ({new_AGEMA_signal_11022, new_AGEMA_signal_11021, new_AGEMA_signal_11020, SubBytesIns_Inst_Sbox_12_M46}), .b ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, new_AGEMA_signal_11650, SubBytesIns_Inst_Sbox_12_L3}), .c ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, new_AGEMA_signal_12199, SubBytesIns_Inst_Sbox_12_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L8_U1 ( .a ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, new_AGEMA_signal_10318, SubBytesIns_Inst_Sbox_12_M51}), .b ({new_AGEMA_signal_10329, new_AGEMA_signal_10328, new_AGEMA_signal_10327, SubBytesIns_Inst_Sbox_12_M59}), .c ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, new_AGEMA_signal_11047, SubBytesIns_Inst_Sbox_12_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L9_U1 ( .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, new_AGEMA_signal_11026, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, new_AGEMA_signal_11641, SubBytesIns_Inst_Sbox_12_M53}), .c ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, new_AGEMA_signal_12202, SubBytesIns_Inst_Sbox_12_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L10_U1 ( .a ({new_AGEMA_signal_11643, new_AGEMA_signal_11642, new_AGEMA_signal_11641, SubBytesIns_Inst_Sbox_12_M53}), .b ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, new_AGEMA_signal_11653, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, new_AGEMA_signal_12205, SubBytesIns_Inst_Sbox_12_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L11_U1 ( .a ({new_AGEMA_signal_10332, new_AGEMA_signal_10331, new_AGEMA_signal_10330, SubBytesIns_Inst_Sbox_12_M60}), .b ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, new_AGEMA_signal_11647, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, new_AGEMA_signal_12208, SubBytesIns_Inst_Sbox_12_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L12_U1 ( .a ({new_AGEMA_signal_10314, new_AGEMA_signal_10313, new_AGEMA_signal_10312, SubBytesIns_Inst_Sbox_12_M48}), .b ({new_AGEMA_signal_10320, new_AGEMA_signal_10319, new_AGEMA_signal_10318, SubBytesIns_Inst_Sbox_12_M51}), .c ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, new_AGEMA_signal_11050, SubBytesIns_Inst_Sbox_12_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L13_U1 ( .a ({new_AGEMA_signal_10317, new_AGEMA_signal_10316, new_AGEMA_signal_10315, SubBytesIns_Inst_Sbox_12_M50}), .b ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_12831, new_AGEMA_signal_12830, new_AGEMA_signal_12829, SubBytesIns_Inst_Sbox_12_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L14_U1 ( .a ({new_AGEMA_signal_11028, new_AGEMA_signal_11027, new_AGEMA_signal_11026, SubBytesIns_Inst_Sbox_12_M52}), .b ({new_AGEMA_signal_11040, new_AGEMA_signal_11039, new_AGEMA_signal_11038, SubBytesIns_Inst_Sbox_12_M61}), .c ({new_AGEMA_signal_11661, new_AGEMA_signal_11660, new_AGEMA_signal_11659, SubBytesIns_Inst_Sbox_12_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L15_U1 ( .a ({new_AGEMA_signal_11034, new_AGEMA_signal_11033, new_AGEMA_signal_11032, SubBytesIns_Inst_Sbox_12_M55}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, new_AGEMA_signal_11662, SubBytesIns_Inst_Sbox_12_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L16_U1 ( .a ({new_AGEMA_signal_10323, new_AGEMA_signal_10322, new_AGEMA_signal_10321, SubBytesIns_Inst_Sbox_12_M56}), .b ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}), .c ({new_AGEMA_signal_12834, new_AGEMA_signal_12833, new_AGEMA_signal_12832, SubBytesIns_Inst_Sbox_12_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L17_U1 ( .a ({new_AGEMA_signal_10326, new_AGEMA_signal_10325, new_AGEMA_signal_10324, SubBytesIns_Inst_Sbox_12_M57}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_11667, new_AGEMA_signal_11666, new_AGEMA_signal_11665, SubBytesIns_Inst_Sbox_12_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L18_U1 ( .a ({new_AGEMA_signal_11037, new_AGEMA_signal_11036, new_AGEMA_signal_11035, SubBytesIns_Inst_Sbox_12_M58}), .b ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, new_AGEMA_signal_11047, SubBytesIns_Inst_Sbox_12_L8}), .c ({new_AGEMA_signal_11670, new_AGEMA_signal_11669, new_AGEMA_signal_11668, SubBytesIns_Inst_Sbox_12_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L19_U1 ( .a ({new_AGEMA_signal_11043, new_AGEMA_signal_11042, new_AGEMA_signal_11041, SubBytesIns_Inst_Sbox_12_M63}), .b ({new_AGEMA_signal_11655, new_AGEMA_signal_11654, new_AGEMA_signal_11653, SubBytesIns_Inst_Sbox_12_L4}), .c ({new_AGEMA_signal_12213, new_AGEMA_signal_12212, new_AGEMA_signal_12211, SubBytesIns_Inst_Sbox_12_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L20_U1 ( .a ({new_AGEMA_signal_12195, new_AGEMA_signal_12194, new_AGEMA_signal_12193, SubBytesIns_Inst_Sbox_12_L0}), .b ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .c ({new_AGEMA_signal_12837, new_AGEMA_signal_12836, new_AGEMA_signal_12835, SubBytesIns_Inst_Sbox_12_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L21_U1 ( .a ({new_AGEMA_signal_11046, new_AGEMA_signal_11045, new_AGEMA_signal_11044, SubBytesIns_Inst_Sbox_12_L1}), .b ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, new_AGEMA_signal_12199, SubBytesIns_Inst_Sbox_12_L7}), .c ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, new_AGEMA_signal_12838, SubBytesIns_Inst_Sbox_12_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L22_U1 ( .a ({new_AGEMA_signal_11652, new_AGEMA_signal_11651, new_AGEMA_signal_11650, SubBytesIns_Inst_Sbox_12_L3}), .b ({new_AGEMA_signal_11052, new_AGEMA_signal_11051, new_AGEMA_signal_11050, SubBytesIns_Inst_Sbox_12_L12}), .c ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, new_AGEMA_signal_12214, SubBytesIns_Inst_Sbox_12_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L23_U1 ( .a ({new_AGEMA_signal_11670, new_AGEMA_signal_11669, new_AGEMA_signal_11668, SubBytesIns_Inst_Sbox_12_L18}), .b ({new_AGEMA_signal_11649, new_AGEMA_signal_11648, new_AGEMA_signal_11647, SubBytesIns_Inst_Sbox_12_L2}), .c ({new_AGEMA_signal_12219, new_AGEMA_signal_12218, new_AGEMA_signal_12217, SubBytesIns_Inst_Sbox_12_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L24_U1 ( .a ({new_AGEMA_signal_11664, new_AGEMA_signal_11663, new_AGEMA_signal_11662, SubBytesIns_Inst_Sbox_12_L15}), .b ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, new_AGEMA_signal_12202, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_12843, new_AGEMA_signal_12842, new_AGEMA_signal_12841, SubBytesIns_Inst_Sbox_12_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L25_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, new_AGEMA_signal_12205, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_12846, new_AGEMA_signal_12845, new_AGEMA_signal_12844, SubBytesIns_Inst_Sbox_12_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L26_U1 ( .a ({new_AGEMA_signal_12201, new_AGEMA_signal_12200, new_AGEMA_signal_12199, SubBytesIns_Inst_Sbox_12_L7}), .b ({new_AGEMA_signal_12204, new_AGEMA_signal_12203, new_AGEMA_signal_12202, SubBytesIns_Inst_Sbox_12_L9}), .c ({new_AGEMA_signal_12849, new_AGEMA_signal_12848, new_AGEMA_signal_12847, SubBytesIns_Inst_Sbox_12_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L27_U1 ( .a ({new_AGEMA_signal_11049, new_AGEMA_signal_11048, new_AGEMA_signal_11047, SubBytesIns_Inst_Sbox_12_L8}), .b ({new_AGEMA_signal_12207, new_AGEMA_signal_12206, new_AGEMA_signal_12205, SubBytesIns_Inst_Sbox_12_L10}), .c ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, new_AGEMA_signal_12850, SubBytesIns_Inst_Sbox_12_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L28_U1 ( .a ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, new_AGEMA_signal_12208, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_11661, new_AGEMA_signal_11660, new_AGEMA_signal_11659, SubBytesIns_Inst_Sbox_12_L14}), .c ({new_AGEMA_signal_12855, new_AGEMA_signal_12854, new_AGEMA_signal_12853, SubBytesIns_Inst_Sbox_12_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_L29_U1 ( .a ({new_AGEMA_signal_12210, new_AGEMA_signal_12209, new_AGEMA_signal_12208, SubBytesIns_Inst_Sbox_12_L11}), .b ({new_AGEMA_signal_11667, new_AGEMA_signal_11666, new_AGEMA_signal_11665, SubBytesIns_Inst_Sbox_12_L17}), .c ({new_AGEMA_signal_12858, new_AGEMA_signal_12857, new_AGEMA_signal_12856, SubBytesIns_Inst_Sbox_12_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S0_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12843, new_AGEMA_signal_12842, new_AGEMA_signal_12841, SubBytesIns_Inst_Sbox_12_L24}), .c ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S1_U1 ( .a ({new_AGEMA_signal_12834, new_AGEMA_signal_12833, new_AGEMA_signal_12832, SubBytesIns_Inst_Sbox_12_L16}), .b ({new_AGEMA_signal_12849, new_AGEMA_signal_12848, new_AGEMA_signal_12847, SubBytesIns_Inst_Sbox_12_L26}), .c ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S2_U1 ( .a ({new_AGEMA_signal_12213, new_AGEMA_signal_12212, new_AGEMA_signal_12211, SubBytesIns_Inst_Sbox_12_L19}), .b ({new_AGEMA_signal_12855, new_AGEMA_signal_12854, new_AGEMA_signal_12853, SubBytesIns_Inst_Sbox_12_L28}), .c ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S3_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12840, new_AGEMA_signal_12839, new_AGEMA_signal_12838, SubBytesIns_Inst_Sbox_12_L21}), .c ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S4_U1 ( .a ({new_AGEMA_signal_12837, new_AGEMA_signal_12836, new_AGEMA_signal_12835, SubBytesIns_Inst_Sbox_12_L20}), .b ({new_AGEMA_signal_12216, new_AGEMA_signal_12215, new_AGEMA_signal_12214, SubBytesIns_Inst_Sbox_12_L22}), .c ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S5_U1 ( .a ({new_AGEMA_signal_12846, new_AGEMA_signal_12845, new_AGEMA_signal_12844, SubBytesIns_Inst_Sbox_12_L25}), .b ({new_AGEMA_signal_12858, new_AGEMA_signal_12857, new_AGEMA_signal_12856, SubBytesIns_Inst_Sbox_12_L29}), .c ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S6_U1 ( .a ({new_AGEMA_signal_12831, new_AGEMA_signal_12830, new_AGEMA_signal_12829, SubBytesIns_Inst_Sbox_12_L13}), .b ({new_AGEMA_signal_12852, new_AGEMA_signal_12851, new_AGEMA_signal_12850, SubBytesIns_Inst_Sbox_12_L27}), .c ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_12_XOR_S7_U1 ( .a ({new_AGEMA_signal_12198, new_AGEMA_signal_12197, new_AGEMA_signal_12196, SubBytesIns_Inst_Sbox_12_L6}), .b ({new_AGEMA_signal_12219, new_AGEMA_signal_12218, new_AGEMA_signal_12217, SubBytesIns_Inst_Sbox_12_L23}), .c ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M46_U1 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, new_AGEMA_signal_10342, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_6711, new_AGEMA_signal_6710, new_AGEMA_signal_6709, SubBytesIns_Inst_Sbox_13_T6}), .clk (clk), .r ({Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324]}), .c ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, new_AGEMA_signal_11056, SubBytesIns_Inst_Sbox_13_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M47_U1 ( .a ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_7446, new_AGEMA_signal_7445, new_AGEMA_signal_7444, SubBytesIns_Inst_Sbox_13_T8}), .clk (clk), .r ({Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330]}), .c ({new_AGEMA_signal_10347, new_AGEMA_signal_10346, new_AGEMA_signal_10345, SubBytesIns_Inst_Sbox_13_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M48_U1 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .b ({ciphertext_s3[104], ciphertext_s2[104], ciphertext_s1[104], ciphertext_s0[104]}), .clk (clk), .r ({Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336]}), .c ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, new_AGEMA_signal_10348, SubBytesIns_Inst_Sbox_13_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M49_U1 ( .a ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, new_AGEMA_signal_10339, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_6723, new_AGEMA_signal_6722, new_AGEMA_signal_6721, SubBytesIns_Inst_Sbox_13_T16}), .clk (clk), .r ({Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342]}), .c ({new_AGEMA_signal_11061, new_AGEMA_signal_11060, new_AGEMA_signal_11059, SubBytesIns_Inst_Sbox_13_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M50_U1 ( .a ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_6714, new_AGEMA_signal_6713, new_AGEMA_signal_6712, SubBytesIns_Inst_Sbox_13_T9}), .clk (clk), .r ({Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348]}), .c ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, new_AGEMA_signal_10351, SubBytesIns_Inst_Sbox_13_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M51_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_7455, new_AGEMA_signal_7454, new_AGEMA_signal_7453, SubBytesIns_Inst_Sbox_13_T17}), .clk (clk), .r ({Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354]}), .c ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, new_AGEMA_signal_10354, SubBytesIns_Inst_Sbox_13_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M52_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_6720, new_AGEMA_signal_6719, new_AGEMA_signal_6718, SubBytesIns_Inst_Sbox_13_T15}), .clk (clk), .r ({Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360]}), .c ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, new_AGEMA_signal_11062, SubBytesIns_Inst_Sbox_13_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M53_U1 ( .a ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, new_AGEMA_signal_11053, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_6732, new_AGEMA_signal_6731, new_AGEMA_signal_6730, SubBytesIns_Inst_Sbox_13_T27}), .clk (clk), .r ({Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366]}), .c ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, new_AGEMA_signal_11671, SubBytesIns_Inst_Sbox_13_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M54_U1 ( .a ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_7449, new_AGEMA_signal_7448, new_AGEMA_signal_7447, SubBytesIns_Inst_Sbox_13_T10}), .clk (clk), .r ({Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372]}), .c ({new_AGEMA_signal_11067, new_AGEMA_signal_11066, new_AGEMA_signal_11065, SubBytesIns_Inst_Sbox_13_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M55_U1 ( .a ({new_AGEMA_signal_10344, new_AGEMA_signal_10343, new_AGEMA_signal_10342, SubBytesIns_Inst_Sbox_13_M44}), .b ({new_AGEMA_signal_6717, new_AGEMA_signal_6716, new_AGEMA_signal_6715, SubBytesIns_Inst_Sbox_13_T13}), .clk (clk), .r ({Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378]}), .c ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, new_AGEMA_signal_11068, SubBytesIns_Inst_Sbox_13_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M56_U1 ( .a ({new_AGEMA_signal_9696, new_AGEMA_signal_9695, new_AGEMA_signal_9694, SubBytesIns_Inst_Sbox_13_M40}), .b ({new_AGEMA_signal_7461, new_AGEMA_signal_7460, new_AGEMA_signal_7459, SubBytesIns_Inst_Sbox_13_T23}), .clk (clk), .r ({Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384]}), .c ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, new_AGEMA_signal_10357, SubBytesIns_Inst_Sbox_13_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M57_U1 ( .a ({new_AGEMA_signal_9693, new_AGEMA_signal_9692, new_AGEMA_signal_9691, SubBytesIns_Inst_Sbox_13_M39}), .b ({new_AGEMA_signal_6726, new_AGEMA_signal_6725, new_AGEMA_signal_6724, SubBytesIns_Inst_Sbox_13_T19}), .clk (clk), .r ({Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390]}), .c ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, new_AGEMA_signal_10360, SubBytesIns_Inst_Sbox_13_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M58_U1 ( .a ({new_AGEMA_signal_10341, new_AGEMA_signal_10340, new_AGEMA_signal_10339, SubBytesIns_Inst_Sbox_13_M43}), .b ({new_AGEMA_signal_6219, new_AGEMA_signal_6218, new_AGEMA_signal_6217, SubBytesIns_Inst_Sbox_13_T3}), .clk (clk), .r ({Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396]}), .c ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, new_AGEMA_signal_11071, SubBytesIns_Inst_Sbox_13_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M59_U1 ( .a ({new_AGEMA_signal_9690, new_AGEMA_signal_9689, new_AGEMA_signal_9688, SubBytesIns_Inst_Sbox_13_M38}), .b ({new_AGEMA_signal_6729, new_AGEMA_signal_6728, new_AGEMA_signal_6727, SubBytesIns_Inst_Sbox_13_T22}), .clk (clk), .r ({Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402]}), .c ({new_AGEMA_signal_10365, new_AGEMA_signal_10364, new_AGEMA_signal_10363, SubBytesIns_Inst_Sbox_13_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M60_U1 ( .a ({new_AGEMA_signal_9687, new_AGEMA_signal_9686, new_AGEMA_signal_9685, SubBytesIns_Inst_Sbox_13_M37}), .b ({new_AGEMA_signal_7458, new_AGEMA_signal_7457, new_AGEMA_signal_7456, SubBytesIns_Inst_Sbox_13_T20}), .clk (clk), .r ({Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408]}), .c ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, new_AGEMA_signal_10366, SubBytesIns_Inst_Sbox_13_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M61_U1 ( .a ({new_AGEMA_signal_10338, new_AGEMA_signal_10337, new_AGEMA_signal_10336, SubBytesIns_Inst_Sbox_13_M42}), .b ({new_AGEMA_signal_6213, new_AGEMA_signal_6212, new_AGEMA_signal_6211, SubBytesIns_Inst_Sbox_13_T1}), .clk (clk), .r ({Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414]}), .c ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M62_U1 ( .a ({new_AGEMA_signal_11055, new_AGEMA_signal_11054, new_AGEMA_signal_11053, SubBytesIns_Inst_Sbox_13_M45}), .b ({new_AGEMA_signal_6222, new_AGEMA_signal_6221, new_AGEMA_signal_6220, SubBytesIns_Inst_Sbox_13_T4}), .clk (clk), .r ({Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420]}), .c ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, new_AGEMA_signal_11674, SubBytesIns_Inst_Sbox_13_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_AND_M63_U1 ( .a ({new_AGEMA_signal_10335, new_AGEMA_signal_10334, new_AGEMA_signal_10333, SubBytesIns_Inst_Sbox_13_M41}), .b ({new_AGEMA_signal_6216, new_AGEMA_signal_6215, new_AGEMA_signal_6214, SubBytesIns_Inst_Sbox_13_T2}), .clk (clk), .r ({Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426]}), .c ({new_AGEMA_signal_11079, new_AGEMA_signal_11078, new_AGEMA_signal_11077, SubBytesIns_Inst_Sbox_13_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L0_U1 ( .a ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}), .b ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, new_AGEMA_signal_11674, SubBytesIns_Inst_Sbox_13_M62}), .c ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L1_U1 ( .a ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, new_AGEMA_signal_10351, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, new_AGEMA_signal_10357, SubBytesIns_Inst_Sbox_13_M56}), .c ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L2_U1 ( .a ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, new_AGEMA_signal_11056, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, new_AGEMA_signal_10348, SubBytesIns_Inst_Sbox_13_M48}), .c ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, new_AGEMA_signal_11677, SubBytesIns_Inst_Sbox_13_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L3_U1 ( .a ({new_AGEMA_signal_10347, new_AGEMA_signal_10346, new_AGEMA_signal_10345, SubBytesIns_Inst_Sbox_13_M47}), .b ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, new_AGEMA_signal_11068, SubBytesIns_Inst_Sbox_13_M55}), .c ({new_AGEMA_signal_11682, new_AGEMA_signal_11681, new_AGEMA_signal_11680, SubBytesIns_Inst_Sbox_13_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L4_U1 ( .a ({new_AGEMA_signal_11067, new_AGEMA_signal_11066, new_AGEMA_signal_11065, SubBytesIns_Inst_Sbox_13_M54}), .b ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, new_AGEMA_signal_11071, SubBytesIns_Inst_Sbox_13_M58}), .c ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, new_AGEMA_signal_11683, SubBytesIns_Inst_Sbox_13_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L5_U1 ( .a ({new_AGEMA_signal_11061, new_AGEMA_signal_11060, new_AGEMA_signal_11059, SubBytesIns_Inst_Sbox_13_M49}), .b ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, new_AGEMA_signal_11686, SubBytesIns_Inst_Sbox_13_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L6_U1 ( .a ({new_AGEMA_signal_11676, new_AGEMA_signal_11675, new_AGEMA_signal_11674, SubBytesIns_Inst_Sbox_13_M62}), .b ({new_AGEMA_signal_11688, new_AGEMA_signal_11687, new_AGEMA_signal_11686, SubBytesIns_Inst_Sbox_13_L5}), .c ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L7_U1 ( .a ({new_AGEMA_signal_11058, new_AGEMA_signal_11057, new_AGEMA_signal_11056, SubBytesIns_Inst_Sbox_13_M46}), .b ({new_AGEMA_signal_11682, new_AGEMA_signal_11681, new_AGEMA_signal_11680, SubBytesIns_Inst_Sbox_13_L3}), .c ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, new_AGEMA_signal_12226, SubBytesIns_Inst_Sbox_13_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L8_U1 ( .a ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, new_AGEMA_signal_10354, SubBytesIns_Inst_Sbox_13_M51}), .b ({new_AGEMA_signal_10365, new_AGEMA_signal_10364, new_AGEMA_signal_10363, SubBytesIns_Inst_Sbox_13_M59}), .c ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, new_AGEMA_signal_11083, SubBytesIns_Inst_Sbox_13_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L9_U1 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, new_AGEMA_signal_11062, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, new_AGEMA_signal_11671, SubBytesIns_Inst_Sbox_13_M53}), .c ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, new_AGEMA_signal_12229, SubBytesIns_Inst_Sbox_13_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L10_U1 ( .a ({new_AGEMA_signal_11673, new_AGEMA_signal_11672, new_AGEMA_signal_11671, SubBytesIns_Inst_Sbox_13_M53}), .b ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, new_AGEMA_signal_11683, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, new_AGEMA_signal_12232, SubBytesIns_Inst_Sbox_13_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L11_U1 ( .a ({new_AGEMA_signal_10368, new_AGEMA_signal_10367, new_AGEMA_signal_10366, SubBytesIns_Inst_Sbox_13_M60}), .b ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, new_AGEMA_signal_11677, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, new_AGEMA_signal_12235, SubBytesIns_Inst_Sbox_13_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L12_U1 ( .a ({new_AGEMA_signal_10350, new_AGEMA_signal_10349, new_AGEMA_signal_10348, SubBytesIns_Inst_Sbox_13_M48}), .b ({new_AGEMA_signal_10356, new_AGEMA_signal_10355, new_AGEMA_signal_10354, SubBytesIns_Inst_Sbox_13_M51}), .c ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, new_AGEMA_signal_11086, SubBytesIns_Inst_Sbox_13_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L13_U1 ( .a ({new_AGEMA_signal_10353, new_AGEMA_signal_10352, new_AGEMA_signal_10351, SubBytesIns_Inst_Sbox_13_M50}), .b ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_12864, new_AGEMA_signal_12863, new_AGEMA_signal_12862, SubBytesIns_Inst_Sbox_13_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L14_U1 ( .a ({new_AGEMA_signal_11064, new_AGEMA_signal_11063, new_AGEMA_signal_11062, SubBytesIns_Inst_Sbox_13_M52}), .b ({new_AGEMA_signal_11076, new_AGEMA_signal_11075, new_AGEMA_signal_11074, SubBytesIns_Inst_Sbox_13_M61}), .c ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, new_AGEMA_signal_11689, SubBytesIns_Inst_Sbox_13_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L15_U1 ( .a ({new_AGEMA_signal_11070, new_AGEMA_signal_11069, new_AGEMA_signal_11068, SubBytesIns_Inst_Sbox_13_M55}), .b ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_11694, new_AGEMA_signal_11693, new_AGEMA_signal_11692, SubBytesIns_Inst_Sbox_13_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L16_U1 ( .a ({new_AGEMA_signal_10359, new_AGEMA_signal_10358, new_AGEMA_signal_10357, SubBytesIns_Inst_Sbox_13_M56}), .b ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}), .c ({new_AGEMA_signal_12867, new_AGEMA_signal_12866, new_AGEMA_signal_12865, SubBytesIns_Inst_Sbox_13_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L17_U1 ( .a ({new_AGEMA_signal_10362, new_AGEMA_signal_10361, new_AGEMA_signal_10360, SubBytesIns_Inst_Sbox_13_M57}), .b ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_11697, new_AGEMA_signal_11696, new_AGEMA_signal_11695, SubBytesIns_Inst_Sbox_13_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L18_U1 ( .a ({new_AGEMA_signal_11073, new_AGEMA_signal_11072, new_AGEMA_signal_11071, SubBytesIns_Inst_Sbox_13_M58}), .b ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, new_AGEMA_signal_11083, SubBytesIns_Inst_Sbox_13_L8}), .c ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, new_AGEMA_signal_11698, SubBytesIns_Inst_Sbox_13_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L19_U1 ( .a ({new_AGEMA_signal_11079, new_AGEMA_signal_11078, new_AGEMA_signal_11077, SubBytesIns_Inst_Sbox_13_M63}), .b ({new_AGEMA_signal_11685, new_AGEMA_signal_11684, new_AGEMA_signal_11683, SubBytesIns_Inst_Sbox_13_L4}), .c ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, new_AGEMA_signal_12238, SubBytesIns_Inst_Sbox_13_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L20_U1 ( .a ({new_AGEMA_signal_12222, new_AGEMA_signal_12221, new_AGEMA_signal_12220, SubBytesIns_Inst_Sbox_13_L0}), .b ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .c ({new_AGEMA_signal_12870, new_AGEMA_signal_12869, new_AGEMA_signal_12868, SubBytesIns_Inst_Sbox_13_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L21_U1 ( .a ({new_AGEMA_signal_11082, new_AGEMA_signal_11081, new_AGEMA_signal_11080, SubBytesIns_Inst_Sbox_13_L1}), .b ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, new_AGEMA_signal_12226, SubBytesIns_Inst_Sbox_13_L7}), .c ({new_AGEMA_signal_12873, new_AGEMA_signal_12872, new_AGEMA_signal_12871, SubBytesIns_Inst_Sbox_13_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L22_U1 ( .a ({new_AGEMA_signal_11682, new_AGEMA_signal_11681, new_AGEMA_signal_11680, SubBytesIns_Inst_Sbox_13_L3}), .b ({new_AGEMA_signal_11088, new_AGEMA_signal_11087, new_AGEMA_signal_11086, SubBytesIns_Inst_Sbox_13_L12}), .c ({new_AGEMA_signal_12243, new_AGEMA_signal_12242, new_AGEMA_signal_12241, SubBytesIns_Inst_Sbox_13_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L23_U1 ( .a ({new_AGEMA_signal_11700, new_AGEMA_signal_11699, new_AGEMA_signal_11698, SubBytesIns_Inst_Sbox_13_L18}), .b ({new_AGEMA_signal_11679, new_AGEMA_signal_11678, new_AGEMA_signal_11677, SubBytesIns_Inst_Sbox_13_L2}), .c ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, new_AGEMA_signal_12244, SubBytesIns_Inst_Sbox_13_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L24_U1 ( .a ({new_AGEMA_signal_11694, new_AGEMA_signal_11693, new_AGEMA_signal_11692, SubBytesIns_Inst_Sbox_13_L15}), .b ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, new_AGEMA_signal_12229, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_12876, new_AGEMA_signal_12875, new_AGEMA_signal_12874, SubBytesIns_Inst_Sbox_13_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L25_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, new_AGEMA_signal_12232, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_12879, new_AGEMA_signal_12878, new_AGEMA_signal_12877, SubBytesIns_Inst_Sbox_13_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L26_U1 ( .a ({new_AGEMA_signal_12228, new_AGEMA_signal_12227, new_AGEMA_signal_12226, SubBytesIns_Inst_Sbox_13_L7}), .b ({new_AGEMA_signal_12231, new_AGEMA_signal_12230, new_AGEMA_signal_12229, SubBytesIns_Inst_Sbox_13_L9}), .c ({new_AGEMA_signal_12882, new_AGEMA_signal_12881, new_AGEMA_signal_12880, SubBytesIns_Inst_Sbox_13_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L27_U1 ( .a ({new_AGEMA_signal_11085, new_AGEMA_signal_11084, new_AGEMA_signal_11083, SubBytesIns_Inst_Sbox_13_L8}), .b ({new_AGEMA_signal_12234, new_AGEMA_signal_12233, new_AGEMA_signal_12232, SubBytesIns_Inst_Sbox_13_L10}), .c ({new_AGEMA_signal_12885, new_AGEMA_signal_12884, new_AGEMA_signal_12883, SubBytesIns_Inst_Sbox_13_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L28_U1 ( .a ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, new_AGEMA_signal_12235, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_11691, new_AGEMA_signal_11690, new_AGEMA_signal_11689, SubBytesIns_Inst_Sbox_13_L14}), .c ({new_AGEMA_signal_12888, new_AGEMA_signal_12887, new_AGEMA_signal_12886, SubBytesIns_Inst_Sbox_13_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_L29_U1 ( .a ({new_AGEMA_signal_12237, new_AGEMA_signal_12236, new_AGEMA_signal_12235, SubBytesIns_Inst_Sbox_13_L11}), .b ({new_AGEMA_signal_11697, new_AGEMA_signal_11696, new_AGEMA_signal_11695, SubBytesIns_Inst_Sbox_13_L17}), .c ({new_AGEMA_signal_12891, new_AGEMA_signal_12890, new_AGEMA_signal_12889, SubBytesIns_Inst_Sbox_13_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S0_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12876, new_AGEMA_signal_12875, new_AGEMA_signal_12874, SubBytesIns_Inst_Sbox_13_L24}), .c ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S1_U1 ( .a ({new_AGEMA_signal_12867, new_AGEMA_signal_12866, new_AGEMA_signal_12865, SubBytesIns_Inst_Sbox_13_L16}), .b ({new_AGEMA_signal_12882, new_AGEMA_signal_12881, new_AGEMA_signal_12880, SubBytesIns_Inst_Sbox_13_L26}), .c ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S2_U1 ( .a ({new_AGEMA_signal_12240, new_AGEMA_signal_12239, new_AGEMA_signal_12238, SubBytesIns_Inst_Sbox_13_L19}), .b ({new_AGEMA_signal_12888, new_AGEMA_signal_12887, new_AGEMA_signal_12886, SubBytesIns_Inst_Sbox_13_L28}), .c ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S3_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12873, new_AGEMA_signal_12872, new_AGEMA_signal_12871, SubBytesIns_Inst_Sbox_13_L21}), .c ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S4_U1 ( .a ({new_AGEMA_signal_12870, new_AGEMA_signal_12869, new_AGEMA_signal_12868, SubBytesIns_Inst_Sbox_13_L20}), .b ({new_AGEMA_signal_12243, new_AGEMA_signal_12242, new_AGEMA_signal_12241, SubBytesIns_Inst_Sbox_13_L22}), .c ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S5_U1 ( .a ({new_AGEMA_signal_12879, new_AGEMA_signal_12878, new_AGEMA_signal_12877, SubBytesIns_Inst_Sbox_13_L25}), .b ({new_AGEMA_signal_12891, new_AGEMA_signal_12890, new_AGEMA_signal_12889, SubBytesIns_Inst_Sbox_13_L29}), .c ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S6_U1 ( .a ({new_AGEMA_signal_12864, new_AGEMA_signal_12863, new_AGEMA_signal_12862, SubBytesIns_Inst_Sbox_13_L13}), .b ({new_AGEMA_signal_12885, new_AGEMA_signal_12884, new_AGEMA_signal_12883, SubBytesIns_Inst_Sbox_13_L27}), .c ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_13_XOR_S7_U1 ( .a ({new_AGEMA_signal_12225, new_AGEMA_signal_12224, new_AGEMA_signal_12223, SubBytesIns_Inst_Sbox_13_L6}), .b ({new_AGEMA_signal_12246, new_AGEMA_signal_12245, new_AGEMA_signal_12244, SubBytesIns_Inst_Sbox_13_L23}), .c ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M46_U1 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, new_AGEMA_signal_10378, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_6735, new_AGEMA_signal_6734, new_AGEMA_signal_6733, SubBytesIns_Inst_Sbox_14_T6}), .clk (clk), .r ({Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432]}), .c ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, new_AGEMA_signal_11092, SubBytesIns_Inst_Sbox_14_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M47_U1 ( .a ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_7485, new_AGEMA_signal_7484, new_AGEMA_signal_7483, SubBytesIns_Inst_Sbox_14_T8}), .clk (clk), .r ({Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438]}), .c ({new_AGEMA_signal_10383, new_AGEMA_signal_10382, new_AGEMA_signal_10381, SubBytesIns_Inst_Sbox_14_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M48_U1 ( .a ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .b ({ciphertext_s3[112], ciphertext_s2[112], ciphertext_s1[112], ciphertext_s0[112]}), .clk (clk), .r ({Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444]}), .c ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, new_AGEMA_signal_10384, SubBytesIns_Inst_Sbox_14_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M49_U1 ( .a ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, new_AGEMA_signal_10375, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_6747, new_AGEMA_signal_6746, new_AGEMA_signal_6745, SubBytesIns_Inst_Sbox_14_T16}), .clk (clk), .r ({Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450]}), .c ({new_AGEMA_signal_11097, new_AGEMA_signal_11096, new_AGEMA_signal_11095, SubBytesIns_Inst_Sbox_14_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M50_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_6738, new_AGEMA_signal_6737, new_AGEMA_signal_6736, SubBytesIns_Inst_Sbox_14_T9}), .clk (clk), .r ({Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456]}), .c ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, new_AGEMA_signal_10387, SubBytesIns_Inst_Sbox_14_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M51_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_7494, new_AGEMA_signal_7493, new_AGEMA_signal_7492, SubBytesIns_Inst_Sbox_14_T17}), .clk (clk), .r ({Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462]}), .c ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, new_AGEMA_signal_10390, SubBytesIns_Inst_Sbox_14_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M52_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_6744, new_AGEMA_signal_6743, new_AGEMA_signal_6742, SubBytesIns_Inst_Sbox_14_T15}), .clk (clk), .r ({Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468]}), .c ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, new_AGEMA_signal_11098, SubBytesIns_Inst_Sbox_14_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M53_U1 ( .a ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, new_AGEMA_signal_11089, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_6756, new_AGEMA_signal_6755, new_AGEMA_signal_6754, SubBytesIns_Inst_Sbox_14_T27}), .clk (clk), .r ({Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474]}), .c ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, new_AGEMA_signal_11701, SubBytesIns_Inst_Sbox_14_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M54_U1 ( .a ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_7488, new_AGEMA_signal_7487, new_AGEMA_signal_7486, SubBytesIns_Inst_Sbox_14_T10}), .clk (clk), .r ({Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480]}), .c ({new_AGEMA_signal_11103, new_AGEMA_signal_11102, new_AGEMA_signal_11101, SubBytesIns_Inst_Sbox_14_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M55_U1 ( .a ({new_AGEMA_signal_10380, new_AGEMA_signal_10379, new_AGEMA_signal_10378, SubBytesIns_Inst_Sbox_14_M44}), .b ({new_AGEMA_signal_6741, new_AGEMA_signal_6740, new_AGEMA_signal_6739, SubBytesIns_Inst_Sbox_14_T13}), .clk (clk), .r ({Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486]}), .c ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, new_AGEMA_signal_11104, SubBytesIns_Inst_Sbox_14_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M56_U1 ( .a ({new_AGEMA_signal_9708, new_AGEMA_signal_9707, new_AGEMA_signal_9706, SubBytesIns_Inst_Sbox_14_M40}), .b ({new_AGEMA_signal_7500, new_AGEMA_signal_7499, new_AGEMA_signal_7498, SubBytesIns_Inst_Sbox_14_T23}), .clk (clk), .r ({Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492]}), .c ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, new_AGEMA_signal_10393, SubBytesIns_Inst_Sbox_14_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M57_U1 ( .a ({new_AGEMA_signal_9705, new_AGEMA_signal_9704, new_AGEMA_signal_9703, SubBytesIns_Inst_Sbox_14_M39}), .b ({new_AGEMA_signal_6750, new_AGEMA_signal_6749, new_AGEMA_signal_6748, SubBytesIns_Inst_Sbox_14_T19}), .clk (clk), .r ({Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498]}), .c ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, new_AGEMA_signal_10396, SubBytesIns_Inst_Sbox_14_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M58_U1 ( .a ({new_AGEMA_signal_10377, new_AGEMA_signal_10376, new_AGEMA_signal_10375, SubBytesIns_Inst_Sbox_14_M43}), .b ({new_AGEMA_signal_6249, new_AGEMA_signal_6248, new_AGEMA_signal_6247, SubBytesIns_Inst_Sbox_14_T3}), .clk (clk), .r ({Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504]}), .c ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, new_AGEMA_signal_11107, SubBytesIns_Inst_Sbox_14_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M59_U1 ( .a ({new_AGEMA_signal_9702, new_AGEMA_signal_9701, new_AGEMA_signal_9700, SubBytesIns_Inst_Sbox_14_M38}), .b ({new_AGEMA_signal_6753, new_AGEMA_signal_6752, new_AGEMA_signal_6751, SubBytesIns_Inst_Sbox_14_T22}), .clk (clk), .r ({Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510]}), .c ({new_AGEMA_signal_10401, new_AGEMA_signal_10400, new_AGEMA_signal_10399, SubBytesIns_Inst_Sbox_14_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M60_U1 ( .a ({new_AGEMA_signal_9699, new_AGEMA_signal_9698, new_AGEMA_signal_9697, SubBytesIns_Inst_Sbox_14_M37}), .b ({new_AGEMA_signal_7497, new_AGEMA_signal_7496, new_AGEMA_signal_7495, SubBytesIns_Inst_Sbox_14_T20}), .clk (clk), .r ({Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516]}), .c ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, new_AGEMA_signal_10402, SubBytesIns_Inst_Sbox_14_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M61_U1 ( .a ({new_AGEMA_signal_10374, new_AGEMA_signal_10373, new_AGEMA_signal_10372, SubBytesIns_Inst_Sbox_14_M42}), .b ({new_AGEMA_signal_6243, new_AGEMA_signal_6242, new_AGEMA_signal_6241, SubBytesIns_Inst_Sbox_14_T1}), .clk (clk), .r ({Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522]}), .c ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M62_U1 ( .a ({new_AGEMA_signal_11091, new_AGEMA_signal_11090, new_AGEMA_signal_11089, SubBytesIns_Inst_Sbox_14_M45}), .b ({new_AGEMA_signal_6252, new_AGEMA_signal_6251, new_AGEMA_signal_6250, SubBytesIns_Inst_Sbox_14_T4}), .clk (clk), .r ({Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528]}), .c ({new_AGEMA_signal_11706, new_AGEMA_signal_11705, new_AGEMA_signal_11704, SubBytesIns_Inst_Sbox_14_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_AND_M63_U1 ( .a ({new_AGEMA_signal_10371, new_AGEMA_signal_10370, new_AGEMA_signal_10369, SubBytesIns_Inst_Sbox_14_M41}), .b ({new_AGEMA_signal_6246, new_AGEMA_signal_6245, new_AGEMA_signal_6244, SubBytesIns_Inst_Sbox_14_T2}), .clk (clk), .r ({Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534]}), .c ({new_AGEMA_signal_11115, new_AGEMA_signal_11114, new_AGEMA_signal_11113, SubBytesIns_Inst_Sbox_14_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L0_U1 ( .a ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}), .b ({new_AGEMA_signal_11706, new_AGEMA_signal_11705, new_AGEMA_signal_11704, SubBytesIns_Inst_Sbox_14_M62}), .c ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L1_U1 ( .a ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, new_AGEMA_signal_10387, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, new_AGEMA_signal_10393, SubBytesIns_Inst_Sbox_14_M56}), .c ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L2_U1 ( .a ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, new_AGEMA_signal_11092, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, new_AGEMA_signal_10384, SubBytesIns_Inst_Sbox_14_M48}), .c ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, new_AGEMA_signal_11707, SubBytesIns_Inst_Sbox_14_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L3_U1 ( .a ({new_AGEMA_signal_10383, new_AGEMA_signal_10382, new_AGEMA_signal_10381, SubBytesIns_Inst_Sbox_14_M47}), .b ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, new_AGEMA_signal_11104, SubBytesIns_Inst_Sbox_14_M55}), .c ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, new_AGEMA_signal_11710, SubBytesIns_Inst_Sbox_14_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L4_U1 ( .a ({new_AGEMA_signal_11103, new_AGEMA_signal_11102, new_AGEMA_signal_11101, SubBytesIns_Inst_Sbox_14_M54}), .b ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, new_AGEMA_signal_11107, SubBytesIns_Inst_Sbox_14_M58}), .c ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, new_AGEMA_signal_11713, SubBytesIns_Inst_Sbox_14_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L5_U1 ( .a ({new_AGEMA_signal_11097, new_AGEMA_signal_11096, new_AGEMA_signal_11095, SubBytesIns_Inst_Sbox_14_M49}), .b ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_11718, new_AGEMA_signal_11717, new_AGEMA_signal_11716, SubBytesIns_Inst_Sbox_14_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L6_U1 ( .a ({new_AGEMA_signal_11706, new_AGEMA_signal_11705, new_AGEMA_signal_11704, SubBytesIns_Inst_Sbox_14_M62}), .b ({new_AGEMA_signal_11718, new_AGEMA_signal_11717, new_AGEMA_signal_11716, SubBytesIns_Inst_Sbox_14_L5}), .c ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L7_U1 ( .a ({new_AGEMA_signal_11094, new_AGEMA_signal_11093, new_AGEMA_signal_11092, SubBytesIns_Inst_Sbox_14_M46}), .b ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, new_AGEMA_signal_11710, SubBytesIns_Inst_Sbox_14_L3}), .c ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, new_AGEMA_signal_12253, SubBytesIns_Inst_Sbox_14_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L8_U1 ( .a ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, new_AGEMA_signal_10390, SubBytesIns_Inst_Sbox_14_M51}), .b ({new_AGEMA_signal_10401, new_AGEMA_signal_10400, new_AGEMA_signal_10399, SubBytesIns_Inst_Sbox_14_M59}), .c ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, new_AGEMA_signal_11119, SubBytesIns_Inst_Sbox_14_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L9_U1 ( .a ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, new_AGEMA_signal_11098, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, new_AGEMA_signal_11701, SubBytesIns_Inst_Sbox_14_M53}), .c ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, new_AGEMA_signal_12256, SubBytesIns_Inst_Sbox_14_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L10_U1 ( .a ({new_AGEMA_signal_11703, new_AGEMA_signal_11702, new_AGEMA_signal_11701, SubBytesIns_Inst_Sbox_14_M53}), .b ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, new_AGEMA_signal_11713, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, new_AGEMA_signal_12259, SubBytesIns_Inst_Sbox_14_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L11_U1 ( .a ({new_AGEMA_signal_10404, new_AGEMA_signal_10403, new_AGEMA_signal_10402, SubBytesIns_Inst_Sbox_14_M60}), .b ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, new_AGEMA_signal_11707, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, new_AGEMA_signal_12262, SubBytesIns_Inst_Sbox_14_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L12_U1 ( .a ({new_AGEMA_signal_10386, new_AGEMA_signal_10385, new_AGEMA_signal_10384, SubBytesIns_Inst_Sbox_14_M48}), .b ({new_AGEMA_signal_10392, new_AGEMA_signal_10391, new_AGEMA_signal_10390, SubBytesIns_Inst_Sbox_14_M51}), .c ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, new_AGEMA_signal_11122, SubBytesIns_Inst_Sbox_14_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L13_U1 ( .a ({new_AGEMA_signal_10389, new_AGEMA_signal_10388, new_AGEMA_signal_10387, SubBytesIns_Inst_Sbox_14_M50}), .b ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_12897, new_AGEMA_signal_12896, new_AGEMA_signal_12895, SubBytesIns_Inst_Sbox_14_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L14_U1 ( .a ({new_AGEMA_signal_11100, new_AGEMA_signal_11099, new_AGEMA_signal_11098, SubBytesIns_Inst_Sbox_14_M52}), .b ({new_AGEMA_signal_11112, new_AGEMA_signal_11111, new_AGEMA_signal_11110, SubBytesIns_Inst_Sbox_14_M61}), .c ({new_AGEMA_signal_11721, new_AGEMA_signal_11720, new_AGEMA_signal_11719, SubBytesIns_Inst_Sbox_14_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L15_U1 ( .a ({new_AGEMA_signal_11106, new_AGEMA_signal_11105, new_AGEMA_signal_11104, SubBytesIns_Inst_Sbox_14_M55}), .b ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, new_AGEMA_signal_11722, SubBytesIns_Inst_Sbox_14_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L16_U1 ( .a ({new_AGEMA_signal_10395, new_AGEMA_signal_10394, new_AGEMA_signal_10393, SubBytesIns_Inst_Sbox_14_M56}), .b ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}), .c ({new_AGEMA_signal_12900, new_AGEMA_signal_12899, new_AGEMA_signal_12898, SubBytesIns_Inst_Sbox_14_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L17_U1 ( .a ({new_AGEMA_signal_10398, new_AGEMA_signal_10397, new_AGEMA_signal_10396, SubBytesIns_Inst_Sbox_14_M57}), .b ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_11727, new_AGEMA_signal_11726, new_AGEMA_signal_11725, SubBytesIns_Inst_Sbox_14_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L18_U1 ( .a ({new_AGEMA_signal_11109, new_AGEMA_signal_11108, new_AGEMA_signal_11107, SubBytesIns_Inst_Sbox_14_M58}), .b ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, new_AGEMA_signal_11119, SubBytesIns_Inst_Sbox_14_L8}), .c ({new_AGEMA_signal_11730, new_AGEMA_signal_11729, new_AGEMA_signal_11728, SubBytesIns_Inst_Sbox_14_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L19_U1 ( .a ({new_AGEMA_signal_11115, new_AGEMA_signal_11114, new_AGEMA_signal_11113, SubBytesIns_Inst_Sbox_14_M63}), .b ({new_AGEMA_signal_11715, new_AGEMA_signal_11714, new_AGEMA_signal_11713, SubBytesIns_Inst_Sbox_14_L4}), .c ({new_AGEMA_signal_12267, new_AGEMA_signal_12266, new_AGEMA_signal_12265, SubBytesIns_Inst_Sbox_14_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L20_U1 ( .a ({new_AGEMA_signal_12249, new_AGEMA_signal_12248, new_AGEMA_signal_12247, SubBytesIns_Inst_Sbox_14_L0}), .b ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .c ({new_AGEMA_signal_12903, new_AGEMA_signal_12902, new_AGEMA_signal_12901, SubBytesIns_Inst_Sbox_14_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L21_U1 ( .a ({new_AGEMA_signal_11118, new_AGEMA_signal_11117, new_AGEMA_signal_11116, SubBytesIns_Inst_Sbox_14_L1}), .b ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, new_AGEMA_signal_12253, SubBytesIns_Inst_Sbox_14_L7}), .c ({new_AGEMA_signal_12906, new_AGEMA_signal_12905, new_AGEMA_signal_12904, SubBytesIns_Inst_Sbox_14_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L22_U1 ( .a ({new_AGEMA_signal_11712, new_AGEMA_signal_11711, new_AGEMA_signal_11710, SubBytesIns_Inst_Sbox_14_L3}), .b ({new_AGEMA_signal_11124, new_AGEMA_signal_11123, new_AGEMA_signal_11122, SubBytesIns_Inst_Sbox_14_L12}), .c ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, new_AGEMA_signal_12268, SubBytesIns_Inst_Sbox_14_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L23_U1 ( .a ({new_AGEMA_signal_11730, new_AGEMA_signal_11729, new_AGEMA_signal_11728, SubBytesIns_Inst_Sbox_14_L18}), .b ({new_AGEMA_signal_11709, new_AGEMA_signal_11708, new_AGEMA_signal_11707, SubBytesIns_Inst_Sbox_14_L2}), .c ({new_AGEMA_signal_12273, new_AGEMA_signal_12272, new_AGEMA_signal_12271, SubBytesIns_Inst_Sbox_14_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L24_U1 ( .a ({new_AGEMA_signal_11724, new_AGEMA_signal_11723, new_AGEMA_signal_11722, SubBytesIns_Inst_Sbox_14_L15}), .b ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, new_AGEMA_signal_12256, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_12909, new_AGEMA_signal_12908, new_AGEMA_signal_12907, SubBytesIns_Inst_Sbox_14_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L25_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, new_AGEMA_signal_12259, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_12912, new_AGEMA_signal_12911, new_AGEMA_signal_12910, SubBytesIns_Inst_Sbox_14_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L26_U1 ( .a ({new_AGEMA_signal_12255, new_AGEMA_signal_12254, new_AGEMA_signal_12253, SubBytesIns_Inst_Sbox_14_L7}), .b ({new_AGEMA_signal_12258, new_AGEMA_signal_12257, new_AGEMA_signal_12256, SubBytesIns_Inst_Sbox_14_L9}), .c ({new_AGEMA_signal_12915, new_AGEMA_signal_12914, new_AGEMA_signal_12913, SubBytesIns_Inst_Sbox_14_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L27_U1 ( .a ({new_AGEMA_signal_11121, new_AGEMA_signal_11120, new_AGEMA_signal_11119, SubBytesIns_Inst_Sbox_14_L8}), .b ({new_AGEMA_signal_12261, new_AGEMA_signal_12260, new_AGEMA_signal_12259, SubBytesIns_Inst_Sbox_14_L10}), .c ({new_AGEMA_signal_12918, new_AGEMA_signal_12917, new_AGEMA_signal_12916, SubBytesIns_Inst_Sbox_14_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L28_U1 ( .a ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, new_AGEMA_signal_12262, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_11721, new_AGEMA_signal_11720, new_AGEMA_signal_11719, SubBytesIns_Inst_Sbox_14_L14}), .c ({new_AGEMA_signal_12921, new_AGEMA_signal_12920, new_AGEMA_signal_12919, SubBytesIns_Inst_Sbox_14_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_L29_U1 ( .a ({new_AGEMA_signal_12264, new_AGEMA_signal_12263, new_AGEMA_signal_12262, SubBytesIns_Inst_Sbox_14_L11}), .b ({new_AGEMA_signal_11727, new_AGEMA_signal_11726, new_AGEMA_signal_11725, SubBytesIns_Inst_Sbox_14_L17}), .c ({new_AGEMA_signal_12924, new_AGEMA_signal_12923, new_AGEMA_signal_12922, SubBytesIns_Inst_Sbox_14_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S0_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12909, new_AGEMA_signal_12908, new_AGEMA_signal_12907, SubBytesIns_Inst_Sbox_14_L24}), .c ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S1_U1 ( .a ({new_AGEMA_signal_12900, new_AGEMA_signal_12899, new_AGEMA_signal_12898, SubBytesIns_Inst_Sbox_14_L16}), .b ({new_AGEMA_signal_12915, new_AGEMA_signal_12914, new_AGEMA_signal_12913, SubBytesIns_Inst_Sbox_14_L26}), .c ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S2_U1 ( .a ({new_AGEMA_signal_12267, new_AGEMA_signal_12266, new_AGEMA_signal_12265, SubBytesIns_Inst_Sbox_14_L19}), .b ({new_AGEMA_signal_12921, new_AGEMA_signal_12920, new_AGEMA_signal_12919, SubBytesIns_Inst_Sbox_14_L28}), .c ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S3_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12906, new_AGEMA_signal_12905, new_AGEMA_signal_12904, SubBytesIns_Inst_Sbox_14_L21}), .c ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S4_U1 ( .a ({new_AGEMA_signal_12903, new_AGEMA_signal_12902, new_AGEMA_signal_12901, SubBytesIns_Inst_Sbox_14_L20}), .b ({new_AGEMA_signal_12270, new_AGEMA_signal_12269, new_AGEMA_signal_12268, SubBytesIns_Inst_Sbox_14_L22}), .c ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S5_U1 ( .a ({new_AGEMA_signal_12912, new_AGEMA_signal_12911, new_AGEMA_signal_12910, SubBytesIns_Inst_Sbox_14_L25}), .b ({new_AGEMA_signal_12924, new_AGEMA_signal_12923, new_AGEMA_signal_12922, SubBytesIns_Inst_Sbox_14_L29}), .c ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S6_U1 ( .a ({new_AGEMA_signal_12897, new_AGEMA_signal_12896, new_AGEMA_signal_12895, SubBytesIns_Inst_Sbox_14_L13}), .b ({new_AGEMA_signal_12918, new_AGEMA_signal_12917, new_AGEMA_signal_12916, SubBytesIns_Inst_Sbox_14_L27}), .c ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_14_XOR_S7_U1 ( .a ({new_AGEMA_signal_12252, new_AGEMA_signal_12251, new_AGEMA_signal_12250, SubBytesIns_Inst_Sbox_14_L6}), .b ({new_AGEMA_signal_12273, new_AGEMA_signal_12272, new_AGEMA_signal_12271, SubBytesIns_Inst_Sbox_14_L23}), .c ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M46_U1 ( .a ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, new_AGEMA_signal_10414, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_6759, new_AGEMA_signal_6758, new_AGEMA_signal_6757, SubBytesIns_Inst_Sbox_15_T6}), .clk (clk), .r ({Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540]}), .c ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, new_AGEMA_signal_11128, SubBytesIns_Inst_Sbox_15_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M47_U1 ( .a ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_7524, new_AGEMA_signal_7523, new_AGEMA_signal_7522, SubBytesIns_Inst_Sbox_15_T8}), .clk (clk), .r ({Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546]}), .c ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, new_AGEMA_signal_10417, SubBytesIns_Inst_Sbox_15_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M48_U1 ( .a ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .b ({ciphertext_s3[120], ciphertext_s2[120], ciphertext_s1[120], ciphertext_s0[120]}), .clk (clk), .r ({Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552]}), .c ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, new_AGEMA_signal_10420, SubBytesIns_Inst_Sbox_15_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M49_U1 ( .a ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, new_AGEMA_signal_10411, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_6771, new_AGEMA_signal_6770, new_AGEMA_signal_6769, SubBytesIns_Inst_Sbox_15_T16}), .clk (clk), .r ({Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558]}), .c ({new_AGEMA_signal_11133, new_AGEMA_signal_11132, new_AGEMA_signal_11131, SubBytesIns_Inst_Sbox_15_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M50_U1 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_6762, new_AGEMA_signal_6761, new_AGEMA_signal_6760, SubBytesIns_Inst_Sbox_15_T9}), .clk (clk), .r ({Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564]}), .c ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, new_AGEMA_signal_10423, SubBytesIns_Inst_Sbox_15_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M51_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_7533, new_AGEMA_signal_7532, new_AGEMA_signal_7531, SubBytesIns_Inst_Sbox_15_T17}), .clk (clk), .r ({Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570]}), .c ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, new_AGEMA_signal_10426, SubBytesIns_Inst_Sbox_15_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M52_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_6768, new_AGEMA_signal_6767, new_AGEMA_signal_6766, SubBytesIns_Inst_Sbox_15_T15}), .clk (clk), .r ({Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576]}), .c ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, new_AGEMA_signal_11134, SubBytesIns_Inst_Sbox_15_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M53_U1 ( .a ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, new_AGEMA_signal_11125, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_6780, new_AGEMA_signal_6779, new_AGEMA_signal_6778, SubBytesIns_Inst_Sbox_15_T27}), .clk (clk), .r ({Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582]}), .c ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, new_AGEMA_signal_11731, SubBytesIns_Inst_Sbox_15_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M54_U1 ( .a ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_7527, new_AGEMA_signal_7526, new_AGEMA_signal_7525, SubBytesIns_Inst_Sbox_15_T10}), .clk (clk), .r ({Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588]}), .c ({new_AGEMA_signal_11139, new_AGEMA_signal_11138, new_AGEMA_signal_11137, SubBytesIns_Inst_Sbox_15_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M55_U1 ( .a ({new_AGEMA_signal_10416, new_AGEMA_signal_10415, new_AGEMA_signal_10414, SubBytesIns_Inst_Sbox_15_M44}), .b ({new_AGEMA_signal_6765, new_AGEMA_signal_6764, new_AGEMA_signal_6763, SubBytesIns_Inst_Sbox_15_T13}), .clk (clk), .r ({Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594]}), .c ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, new_AGEMA_signal_11140, SubBytesIns_Inst_Sbox_15_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M56_U1 ( .a ({new_AGEMA_signal_9720, new_AGEMA_signal_9719, new_AGEMA_signal_9718, SubBytesIns_Inst_Sbox_15_M40}), .b ({new_AGEMA_signal_7539, new_AGEMA_signal_7538, new_AGEMA_signal_7537, SubBytesIns_Inst_Sbox_15_T23}), .clk (clk), .r ({Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600]}), .c ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, new_AGEMA_signal_10429, SubBytesIns_Inst_Sbox_15_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M57_U1 ( .a ({new_AGEMA_signal_9717, new_AGEMA_signal_9716, new_AGEMA_signal_9715, SubBytesIns_Inst_Sbox_15_M39}), .b ({new_AGEMA_signal_6774, new_AGEMA_signal_6773, new_AGEMA_signal_6772, SubBytesIns_Inst_Sbox_15_T19}), .clk (clk), .r ({Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606]}), .c ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, new_AGEMA_signal_10432, SubBytesIns_Inst_Sbox_15_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M58_U1 ( .a ({new_AGEMA_signal_10413, new_AGEMA_signal_10412, new_AGEMA_signal_10411, SubBytesIns_Inst_Sbox_15_M43}), .b ({new_AGEMA_signal_6279, new_AGEMA_signal_6278, new_AGEMA_signal_6277, SubBytesIns_Inst_Sbox_15_T3}), .clk (clk), .r ({Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612]}), .c ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, new_AGEMA_signal_11143, SubBytesIns_Inst_Sbox_15_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M59_U1 ( .a ({new_AGEMA_signal_9714, new_AGEMA_signal_9713, new_AGEMA_signal_9712, SubBytesIns_Inst_Sbox_15_M38}), .b ({new_AGEMA_signal_6777, new_AGEMA_signal_6776, new_AGEMA_signal_6775, SubBytesIns_Inst_Sbox_15_T22}), .clk (clk), .r ({Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618]}), .c ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, new_AGEMA_signal_10435, SubBytesIns_Inst_Sbox_15_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M60_U1 ( .a ({new_AGEMA_signal_9711, new_AGEMA_signal_9710, new_AGEMA_signal_9709, SubBytesIns_Inst_Sbox_15_M37}), .b ({new_AGEMA_signal_7536, new_AGEMA_signal_7535, new_AGEMA_signal_7534, SubBytesIns_Inst_Sbox_15_T20}), .clk (clk), .r ({Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624]}), .c ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, new_AGEMA_signal_10438, SubBytesIns_Inst_Sbox_15_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M61_U1 ( .a ({new_AGEMA_signal_10410, new_AGEMA_signal_10409, new_AGEMA_signal_10408, SubBytesIns_Inst_Sbox_15_M42}), .b ({new_AGEMA_signal_6273, new_AGEMA_signal_6272, new_AGEMA_signal_6271, SubBytesIns_Inst_Sbox_15_T1}), .clk (clk), .r ({Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630]}), .c ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M62_U1 ( .a ({new_AGEMA_signal_11127, new_AGEMA_signal_11126, new_AGEMA_signal_11125, SubBytesIns_Inst_Sbox_15_M45}), .b ({new_AGEMA_signal_6282, new_AGEMA_signal_6281, new_AGEMA_signal_6280, SubBytesIns_Inst_Sbox_15_T4}), .clk (clk), .r ({Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636]}), .c ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, new_AGEMA_signal_11734, SubBytesIns_Inst_Sbox_15_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_AND_M63_U1 ( .a ({new_AGEMA_signal_10407, new_AGEMA_signal_10406, new_AGEMA_signal_10405, SubBytesIns_Inst_Sbox_15_M41}), .b ({new_AGEMA_signal_6276, new_AGEMA_signal_6275, new_AGEMA_signal_6274, SubBytesIns_Inst_Sbox_15_T2}), .clk (clk), .r ({Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642]}), .c ({new_AGEMA_signal_11151, new_AGEMA_signal_11150, new_AGEMA_signal_11149, SubBytesIns_Inst_Sbox_15_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L0_U1 ( .a ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}), .b ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, new_AGEMA_signal_11734, SubBytesIns_Inst_Sbox_15_M62}), .c ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L1_U1 ( .a ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, new_AGEMA_signal_10423, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, new_AGEMA_signal_10429, SubBytesIns_Inst_Sbox_15_M56}), .c ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L2_U1 ( .a ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, new_AGEMA_signal_11128, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, new_AGEMA_signal_10420, SubBytesIns_Inst_Sbox_15_M48}), .c ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, new_AGEMA_signal_11737, SubBytesIns_Inst_Sbox_15_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L3_U1 ( .a ({new_AGEMA_signal_10419, new_AGEMA_signal_10418, new_AGEMA_signal_10417, SubBytesIns_Inst_Sbox_15_M47}), .b ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, new_AGEMA_signal_11140, SubBytesIns_Inst_Sbox_15_M55}), .c ({new_AGEMA_signal_11742, new_AGEMA_signal_11741, new_AGEMA_signal_11740, SubBytesIns_Inst_Sbox_15_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L4_U1 ( .a ({new_AGEMA_signal_11139, new_AGEMA_signal_11138, new_AGEMA_signal_11137, SubBytesIns_Inst_Sbox_15_M54}), .b ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, new_AGEMA_signal_11143, SubBytesIns_Inst_Sbox_15_M58}), .c ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, new_AGEMA_signal_11743, SubBytesIns_Inst_Sbox_15_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L5_U1 ( .a ({new_AGEMA_signal_11133, new_AGEMA_signal_11132, new_AGEMA_signal_11131, SubBytesIns_Inst_Sbox_15_M49}), .b ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, new_AGEMA_signal_11746, SubBytesIns_Inst_Sbox_15_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L6_U1 ( .a ({new_AGEMA_signal_11736, new_AGEMA_signal_11735, new_AGEMA_signal_11734, SubBytesIns_Inst_Sbox_15_M62}), .b ({new_AGEMA_signal_11748, new_AGEMA_signal_11747, new_AGEMA_signal_11746, SubBytesIns_Inst_Sbox_15_L5}), .c ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L7_U1 ( .a ({new_AGEMA_signal_11130, new_AGEMA_signal_11129, new_AGEMA_signal_11128, SubBytesIns_Inst_Sbox_15_M46}), .b ({new_AGEMA_signal_11742, new_AGEMA_signal_11741, new_AGEMA_signal_11740, SubBytesIns_Inst_Sbox_15_L3}), .c ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, new_AGEMA_signal_12280, SubBytesIns_Inst_Sbox_15_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L8_U1 ( .a ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, new_AGEMA_signal_10426, SubBytesIns_Inst_Sbox_15_M51}), .b ({new_AGEMA_signal_10437, new_AGEMA_signal_10436, new_AGEMA_signal_10435, SubBytesIns_Inst_Sbox_15_M59}), .c ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, new_AGEMA_signal_11155, SubBytesIns_Inst_Sbox_15_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L9_U1 ( .a ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, new_AGEMA_signal_11134, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, new_AGEMA_signal_11731, SubBytesIns_Inst_Sbox_15_M53}), .c ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, new_AGEMA_signal_12283, SubBytesIns_Inst_Sbox_15_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L10_U1 ( .a ({new_AGEMA_signal_11733, new_AGEMA_signal_11732, new_AGEMA_signal_11731, SubBytesIns_Inst_Sbox_15_M53}), .b ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, new_AGEMA_signal_11743, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, new_AGEMA_signal_12286, SubBytesIns_Inst_Sbox_15_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L11_U1 ( .a ({new_AGEMA_signal_10440, new_AGEMA_signal_10439, new_AGEMA_signal_10438, SubBytesIns_Inst_Sbox_15_M60}), .b ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, new_AGEMA_signal_11737, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, new_AGEMA_signal_12289, SubBytesIns_Inst_Sbox_15_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L12_U1 ( .a ({new_AGEMA_signal_10422, new_AGEMA_signal_10421, new_AGEMA_signal_10420, SubBytesIns_Inst_Sbox_15_M48}), .b ({new_AGEMA_signal_10428, new_AGEMA_signal_10427, new_AGEMA_signal_10426, SubBytesIns_Inst_Sbox_15_M51}), .c ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, new_AGEMA_signal_11158, SubBytesIns_Inst_Sbox_15_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L13_U1 ( .a ({new_AGEMA_signal_10425, new_AGEMA_signal_10424, new_AGEMA_signal_10423, SubBytesIns_Inst_Sbox_15_M50}), .b ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_12930, new_AGEMA_signal_12929, new_AGEMA_signal_12928, SubBytesIns_Inst_Sbox_15_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L14_U1 ( .a ({new_AGEMA_signal_11136, new_AGEMA_signal_11135, new_AGEMA_signal_11134, SubBytesIns_Inst_Sbox_15_M52}), .b ({new_AGEMA_signal_11148, new_AGEMA_signal_11147, new_AGEMA_signal_11146, SubBytesIns_Inst_Sbox_15_M61}), .c ({new_AGEMA_signal_11751, new_AGEMA_signal_11750, new_AGEMA_signal_11749, SubBytesIns_Inst_Sbox_15_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L15_U1 ( .a ({new_AGEMA_signal_11142, new_AGEMA_signal_11141, new_AGEMA_signal_11140, SubBytesIns_Inst_Sbox_15_M55}), .b ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_11754, new_AGEMA_signal_11753, new_AGEMA_signal_11752, SubBytesIns_Inst_Sbox_15_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L16_U1 ( .a ({new_AGEMA_signal_10431, new_AGEMA_signal_10430, new_AGEMA_signal_10429, SubBytesIns_Inst_Sbox_15_M56}), .b ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}), .c ({new_AGEMA_signal_12933, new_AGEMA_signal_12932, new_AGEMA_signal_12931, SubBytesIns_Inst_Sbox_15_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L17_U1 ( .a ({new_AGEMA_signal_10434, new_AGEMA_signal_10433, new_AGEMA_signal_10432, SubBytesIns_Inst_Sbox_15_M57}), .b ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_11757, new_AGEMA_signal_11756, new_AGEMA_signal_11755, SubBytesIns_Inst_Sbox_15_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L18_U1 ( .a ({new_AGEMA_signal_11145, new_AGEMA_signal_11144, new_AGEMA_signal_11143, SubBytesIns_Inst_Sbox_15_M58}), .b ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, new_AGEMA_signal_11155, SubBytesIns_Inst_Sbox_15_L8}), .c ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, new_AGEMA_signal_11758, SubBytesIns_Inst_Sbox_15_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L19_U1 ( .a ({new_AGEMA_signal_11151, new_AGEMA_signal_11150, new_AGEMA_signal_11149, SubBytesIns_Inst_Sbox_15_M63}), .b ({new_AGEMA_signal_11745, new_AGEMA_signal_11744, new_AGEMA_signal_11743, SubBytesIns_Inst_Sbox_15_L4}), .c ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, new_AGEMA_signal_12292, SubBytesIns_Inst_Sbox_15_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L20_U1 ( .a ({new_AGEMA_signal_12276, new_AGEMA_signal_12275, new_AGEMA_signal_12274, SubBytesIns_Inst_Sbox_15_L0}), .b ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .c ({new_AGEMA_signal_12936, new_AGEMA_signal_12935, new_AGEMA_signal_12934, SubBytesIns_Inst_Sbox_15_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L21_U1 ( .a ({new_AGEMA_signal_11154, new_AGEMA_signal_11153, new_AGEMA_signal_11152, SubBytesIns_Inst_Sbox_15_L1}), .b ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, new_AGEMA_signal_12280, SubBytesIns_Inst_Sbox_15_L7}), .c ({new_AGEMA_signal_12939, new_AGEMA_signal_12938, new_AGEMA_signal_12937, SubBytesIns_Inst_Sbox_15_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L22_U1 ( .a ({new_AGEMA_signal_11742, new_AGEMA_signal_11741, new_AGEMA_signal_11740, SubBytesIns_Inst_Sbox_15_L3}), .b ({new_AGEMA_signal_11160, new_AGEMA_signal_11159, new_AGEMA_signal_11158, SubBytesIns_Inst_Sbox_15_L12}), .c ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, new_AGEMA_signal_12295, SubBytesIns_Inst_Sbox_15_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L23_U1 ( .a ({new_AGEMA_signal_11760, new_AGEMA_signal_11759, new_AGEMA_signal_11758, SubBytesIns_Inst_Sbox_15_L18}), .b ({new_AGEMA_signal_11739, new_AGEMA_signal_11738, new_AGEMA_signal_11737, SubBytesIns_Inst_Sbox_15_L2}), .c ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, new_AGEMA_signal_12298, SubBytesIns_Inst_Sbox_15_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L24_U1 ( .a ({new_AGEMA_signal_11754, new_AGEMA_signal_11753, new_AGEMA_signal_11752, SubBytesIns_Inst_Sbox_15_L15}), .b ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, new_AGEMA_signal_12283, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_12942, new_AGEMA_signal_12941, new_AGEMA_signal_12940, SubBytesIns_Inst_Sbox_15_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L25_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, new_AGEMA_signal_12286, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_12945, new_AGEMA_signal_12944, new_AGEMA_signal_12943, SubBytesIns_Inst_Sbox_15_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L26_U1 ( .a ({new_AGEMA_signal_12282, new_AGEMA_signal_12281, new_AGEMA_signal_12280, SubBytesIns_Inst_Sbox_15_L7}), .b ({new_AGEMA_signal_12285, new_AGEMA_signal_12284, new_AGEMA_signal_12283, SubBytesIns_Inst_Sbox_15_L9}), .c ({new_AGEMA_signal_12948, new_AGEMA_signal_12947, new_AGEMA_signal_12946, SubBytesIns_Inst_Sbox_15_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L27_U1 ( .a ({new_AGEMA_signal_11157, new_AGEMA_signal_11156, new_AGEMA_signal_11155, SubBytesIns_Inst_Sbox_15_L8}), .b ({new_AGEMA_signal_12288, new_AGEMA_signal_12287, new_AGEMA_signal_12286, SubBytesIns_Inst_Sbox_15_L10}), .c ({new_AGEMA_signal_12951, new_AGEMA_signal_12950, new_AGEMA_signal_12949, SubBytesIns_Inst_Sbox_15_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L28_U1 ( .a ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, new_AGEMA_signal_12289, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_11751, new_AGEMA_signal_11750, new_AGEMA_signal_11749, SubBytesIns_Inst_Sbox_15_L14}), .c ({new_AGEMA_signal_12954, new_AGEMA_signal_12953, new_AGEMA_signal_12952, SubBytesIns_Inst_Sbox_15_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_L29_U1 ( .a ({new_AGEMA_signal_12291, new_AGEMA_signal_12290, new_AGEMA_signal_12289, SubBytesIns_Inst_Sbox_15_L11}), .b ({new_AGEMA_signal_11757, new_AGEMA_signal_11756, new_AGEMA_signal_11755, SubBytesIns_Inst_Sbox_15_L17}), .c ({new_AGEMA_signal_12957, new_AGEMA_signal_12956, new_AGEMA_signal_12955, SubBytesIns_Inst_Sbox_15_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S0_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12942, new_AGEMA_signal_12941, new_AGEMA_signal_12940, SubBytesIns_Inst_Sbox_15_L24}), .c ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S1_U1 ( .a ({new_AGEMA_signal_12933, new_AGEMA_signal_12932, new_AGEMA_signal_12931, SubBytesIns_Inst_Sbox_15_L16}), .b ({new_AGEMA_signal_12948, new_AGEMA_signal_12947, new_AGEMA_signal_12946, SubBytesIns_Inst_Sbox_15_L26}), .c ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S2_U1 ( .a ({new_AGEMA_signal_12294, new_AGEMA_signal_12293, new_AGEMA_signal_12292, SubBytesIns_Inst_Sbox_15_L19}), .b ({new_AGEMA_signal_12954, new_AGEMA_signal_12953, new_AGEMA_signal_12952, SubBytesIns_Inst_Sbox_15_L28}), .c ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S3_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12939, new_AGEMA_signal_12938, new_AGEMA_signal_12937, SubBytesIns_Inst_Sbox_15_L21}), .c ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S4_U1 ( .a ({new_AGEMA_signal_12936, new_AGEMA_signal_12935, new_AGEMA_signal_12934, SubBytesIns_Inst_Sbox_15_L20}), .b ({new_AGEMA_signal_12297, new_AGEMA_signal_12296, new_AGEMA_signal_12295, SubBytesIns_Inst_Sbox_15_L22}), .c ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S5_U1 ( .a ({new_AGEMA_signal_12945, new_AGEMA_signal_12944, new_AGEMA_signal_12943, SubBytesIns_Inst_Sbox_15_L25}), .b ({new_AGEMA_signal_12957, new_AGEMA_signal_12956, new_AGEMA_signal_12955, SubBytesIns_Inst_Sbox_15_L29}), .c ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S6_U1 ( .a ({new_AGEMA_signal_12930, new_AGEMA_signal_12929, new_AGEMA_signal_12928, SubBytesIns_Inst_Sbox_15_L13}), .b ({new_AGEMA_signal_12951, new_AGEMA_signal_12950, new_AGEMA_signal_12949, SubBytesIns_Inst_Sbox_15_L27}), .c ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) SubBytesIns_Inst_Sbox_15_XOR_S7_U1 ( .a ({new_AGEMA_signal_12279, new_AGEMA_signal_12278, new_AGEMA_signal_12277, SubBytesIns_Inst_Sbox_15_L6}), .b ({new_AGEMA_signal_12300, new_AGEMA_signal_12299, new_AGEMA_signal_12298, SubBytesIns_Inst_Sbox_15_L23}), .c ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U96 ( .a ({new_AGEMA_signal_14811, new_AGEMA_signal_14810, new_AGEMA_signal_14809, MixColumnsIns_MixOneColumnInst_0_n64}), .b ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_15714, new_AGEMA_signal_15713, new_AGEMA_signal_15712, MixColumnsOutput[105]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U95 ( .a ({new_AGEMA_signal_14202, new_AGEMA_signal_14201, new_AGEMA_signal_14200, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_14190, new_AGEMA_signal_14189, new_AGEMA_signal_14188, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_14811, new_AGEMA_signal_14810, new_AGEMA_signal_14809, MixColumnsIns_MixOneColumnInst_0_n64}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U94 ( .a ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, new_AGEMA_signal_14137, MixColumnsIns_MixOneColumnInst_0_n61}), .b ({new_AGEMA_signal_13536, new_AGEMA_signal_13535, new_AGEMA_signal_13534, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_14814, new_AGEMA_signal_14813, new_AGEMA_signal_14812, MixColumnsOutput[104]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U93 ( .a ({new_AGEMA_signal_13566, new_AGEMA_signal_13565, new_AGEMA_signal_13564, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .c ({new_AGEMA_signal_14139, new_AGEMA_signal_14138, new_AGEMA_signal_14137, MixColumnsIns_MixOneColumnInst_0_n61}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U92 ( .a ({new_AGEMA_signal_14142, new_AGEMA_signal_14141, new_AGEMA_signal_14140, MixColumnsIns_MixOneColumnInst_0_n58}), .b ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, new_AGEMA_signal_13507, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_14817, new_AGEMA_signal_14816, new_AGEMA_signal_14815, MixColumnsOutput[103]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U91 ( .a ({new_AGEMA_signal_13542, new_AGEMA_signal_13541, new_AGEMA_signal_13540, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .c ({new_AGEMA_signal_14142, new_AGEMA_signal_14141, new_AGEMA_signal_14140, MixColumnsIns_MixOneColumnInst_0_n58}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U90 ( .a ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, new_AGEMA_signal_14143, MixColumnsIns_MixOneColumnInst_0_n55}), .b ({new_AGEMA_signal_13512, new_AGEMA_signal_13511, new_AGEMA_signal_13510, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_14820, new_AGEMA_signal_14819, new_AGEMA_signal_14818, MixColumnsOutput[102]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U89 ( .a ({new_AGEMA_signal_13548, new_AGEMA_signal_13547, new_AGEMA_signal_13546, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_14145, new_AGEMA_signal_14144, new_AGEMA_signal_14143, MixColumnsIns_MixOneColumnInst_0_n55}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U88 ( .a ({new_AGEMA_signal_14148, new_AGEMA_signal_14147, new_AGEMA_signal_14146, MixColumnsIns_MixOneColumnInst_0_n52}), .b ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, new_AGEMA_signal_13513, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_14823, new_AGEMA_signal_14822, new_AGEMA_signal_14821, MixColumnsOutput[101]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U87 ( .a ({new_AGEMA_signal_13554, new_AGEMA_signal_13553, new_AGEMA_signal_13552, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_14148, new_AGEMA_signal_14147, new_AGEMA_signal_14146, MixColumnsIns_MixOneColumnInst_0_n52}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U86 ( .a ({new_AGEMA_signal_14826, new_AGEMA_signal_14825, new_AGEMA_signal_14824, MixColumnsIns_MixOneColumnInst_0_n49}), .b ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, new_AGEMA_signal_14161, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_15717, new_AGEMA_signal_15716, new_AGEMA_signal_15715, MixColumnsOutput[100]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U85 ( .a ({new_AGEMA_signal_14220, new_AGEMA_signal_14219, new_AGEMA_signal_14218, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_14826, new_AGEMA_signal_14825, new_AGEMA_signal_14824, MixColumnsIns_MixOneColumnInst_0_n49}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U84 ( .a ({new_AGEMA_signal_14829, new_AGEMA_signal_14828, new_AGEMA_signal_14827, MixColumnsIns_MixOneColumnInst_0_n46}), .b ({new_AGEMA_signal_14166, new_AGEMA_signal_14165, new_AGEMA_signal_14164, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_15720, new_AGEMA_signal_15719, new_AGEMA_signal_15718, MixColumnsOutput[99]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U83 ( .a ({new_AGEMA_signal_14226, new_AGEMA_signal_14225, new_AGEMA_signal_14224, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .c ({new_AGEMA_signal_14829, new_AGEMA_signal_14828, new_AGEMA_signal_14827, MixColumnsIns_MixOneColumnInst_0_n46}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U82 ( .a ({new_AGEMA_signal_14151, new_AGEMA_signal_14150, new_AGEMA_signal_14149, MixColumnsIns_MixOneColumnInst_0_n43}), .b ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, new_AGEMA_signal_13507, MixColumnsIns_MixOneColumnInst_0_n57}), .c ({new_AGEMA_signal_14832, new_AGEMA_signal_14831, new_AGEMA_signal_14830, MixColumnsOutput[127]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U81 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_13509, new_AGEMA_signal_13508, new_AGEMA_signal_13507, MixColumnsIns_MixOneColumnInst_0_n57}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U80 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, new_AGEMA_signal_13519, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_14151, new_AGEMA_signal_14150, new_AGEMA_signal_14149, MixColumnsIns_MixOneColumnInst_0_n43}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U79 ( .a ({new_AGEMA_signal_14154, new_AGEMA_signal_14153, new_AGEMA_signal_14152, MixColumnsIns_MixOneColumnInst_0_n41}), .b ({new_AGEMA_signal_13512, new_AGEMA_signal_13511, new_AGEMA_signal_13510, MixColumnsIns_MixOneColumnInst_0_n54}), .c ({new_AGEMA_signal_14835, new_AGEMA_signal_14834, new_AGEMA_signal_14833, MixColumnsOutput[126]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U78 ( .a ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .b ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_13512, new_AGEMA_signal_13511, new_AGEMA_signal_13510, MixColumnsIns_MixOneColumnInst_0_n54}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U77 ( .a ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_13524, new_AGEMA_signal_13523, new_AGEMA_signal_13522, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_14154, new_AGEMA_signal_14153, new_AGEMA_signal_14152, MixColumnsIns_MixOneColumnInst_0_n41}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U76 ( .a ({new_AGEMA_signal_14157, new_AGEMA_signal_14156, new_AGEMA_signal_14155, MixColumnsIns_MixOneColumnInst_0_n39}), .b ({new_AGEMA_signal_13518, new_AGEMA_signal_13517, new_AGEMA_signal_13516, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_14838, new_AGEMA_signal_14837, new_AGEMA_signal_14836, MixColumnsOutput[98]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U75 ( .a ({new_AGEMA_signal_13560, new_AGEMA_signal_13559, new_AGEMA_signal_13558, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .c ({new_AGEMA_signal_14157, new_AGEMA_signal_14156, new_AGEMA_signal_14155, MixColumnsIns_MixOneColumnInst_0_n39}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U74 ( .a ({new_AGEMA_signal_14160, new_AGEMA_signal_14159, new_AGEMA_signal_14158, MixColumnsIns_MixOneColumnInst_0_n36}), .b ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, new_AGEMA_signal_13513, MixColumnsIns_MixOneColumnInst_0_n51}), .c ({new_AGEMA_signal_14841, new_AGEMA_signal_14840, new_AGEMA_signal_14839, MixColumnsOutput[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U73 ( .a ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_13515, new_AGEMA_signal_13514, new_AGEMA_signal_13513, MixColumnsIns_MixOneColumnInst_0_n51}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U72 ( .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, new_AGEMA_signal_13525, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_14160, new_AGEMA_signal_14159, new_AGEMA_signal_14158, MixColumnsIns_MixOneColumnInst_0_n36}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U71 ( .a ({new_AGEMA_signal_14844, new_AGEMA_signal_14843, new_AGEMA_signal_14842, MixColumnsIns_MixOneColumnInst_0_n34}), .b ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, new_AGEMA_signal_14161, MixColumnsIns_MixOneColumnInst_0_n48}), .c ({new_AGEMA_signal_15723, new_AGEMA_signal_15722, new_AGEMA_signal_15721, MixColumnsOutput[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U70 ( .a ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .b ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, new_AGEMA_signal_13567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}), .c ({new_AGEMA_signal_14163, new_AGEMA_signal_14162, new_AGEMA_signal_14161, MixColumnsIns_MixOneColumnInst_0_n48}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U69 ( .a ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_14184, new_AGEMA_signal_14183, new_AGEMA_signal_14182, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_14844, new_AGEMA_signal_14843, new_AGEMA_signal_14842, MixColumnsIns_MixOneColumnInst_0_n34}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U68 ( .a ({new_AGEMA_signal_14847, new_AGEMA_signal_14846, new_AGEMA_signal_14845, MixColumnsIns_MixOneColumnInst_0_n32}), .b ({new_AGEMA_signal_14166, new_AGEMA_signal_14165, new_AGEMA_signal_14164, MixColumnsIns_MixOneColumnInst_0_n45}), .c ({new_AGEMA_signal_15726, new_AGEMA_signal_15725, new_AGEMA_signal_15724, MixColumnsOutput[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U67 ( .a ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .b ({new_AGEMA_signal_13572, new_AGEMA_signal_13571, new_AGEMA_signal_13570, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}), .c ({new_AGEMA_signal_14166, new_AGEMA_signal_14165, new_AGEMA_signal_14164, MixColumnsIns_MixOneColumnInst_0_n45}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U66 ( .a ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .b ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, new_AGEMA_signal_14191, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_14847, new_AGEMA_signal_14846, new_AGEMA_signal_14845, MixColumnsIns_MixOneColumnInst_0_n32}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U65 ( .a ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, new_AGEMA_signal_14167, MixColumnsIns_MixOneColumnInst_0_n30}), .b ({new_AGEMA_signal_13518, new_AGEMA_signal_13517, new_AGEMA_signal_13516, MixColumnsIns_MixOneColumnInst_0_n38}), .c ({new_AGEMA_signal_14850, new_AGEMA_signal_14849, new_AGEMA_signal_14848, MixColumnsOutput[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U64 ( .a ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .b ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_13518, new_AGEMA_signal_13517, new_AGEMA_signal_13516, MixColumnsIns_MixOneColumnInst_0_n38}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U63 ( .a ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .b ({new_AGEMA_signal_13530, new_AGEMA_signal_13529, new_AGEMA_signal_13528, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_14169, new_AGEMA_signal_14168, new_AGEMA_signal_14167, MixColumnsIns_MixOneColumnInst_0_n30}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U62 ( .a ({new_AGEMA_signal_14853, new_AGEMA_signal_14852, new_AGEMA_signal_14851, MixColumnsIns_MixOneColumnInst_0_n28}), .b ({new_AGEMA_signal_14187, new_AGEMA_signal_14186, new_AGEMA_signal_14185, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_15729, new_AGEMA_signal_15728, new_AGEMA_signal_15727, MixColumnsOutput[121]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U61 ( .a ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, new_AGEMA_signal_14197, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_14853, new_AGEMA_signal_14852, new_AGEMA_signal_14851, MixColumnsIns_MixOneColumnInst_0_n28}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U60 ( .a ({new_AGEMA_signal_14172, new_AGEMA_signal_14171, new_AGEMA_signal_14170, MixColumnsIns_MixOneColumnInst_0_n25}), .b ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, new_AGEMA_signal_13531, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_14856, new_AGEMA_signal_14855, new_AGEMA_signal_14854, MixColumnsOutput[120]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U59 ( .a ({new_AGEMA_signal_13563, new_AGEMA_signal_13562, new_AGEMA_signal_13561, MixColumnsIns_MixOneColumnInst_0_n23}), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .c ({new_AGEMA_signal_14172, new_AGEMA_signal_14171, new_AGEMA_signal_14170, MixColumnsIns_MixOneColumnInst_0_n25}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U58 ( .a ({new_AGEMA_signal_14175, new_AGEMA_signal_14174, new_AGEMA_signal_14173, MixColumnsIns_MixOneColumnInst_0_n22}), .b ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, new_AGEMA_signal_13519, MixColumnsIns_MixOneColumnInst_0_n42}), .c ({new_AGEMA_signal_14859, new_AGEMA_signal_14858, new_AGEMA_signal_14857, MixColumnsOutput[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U57 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_13521, new_AGEMA_signal_13520, new_AGEMA_signal_13519, MixColumnsIns_MixOneColumnInst_0_n42}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U56 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, new_AGEMA_signal_13537, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_14175, new_AGEMA_signal_14174, new_AGEMA_signal_14173, MixColumnsIns_MixOneColumnInst_0_n22}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U55 ( .a ({new_AGEMA_signal_14178, new_AGEMA_signal_14177, new_AGEMA_signal_14176, MixColumnsIns_MixOneColumnInst_0_n20}), .b ({new_AGEMA_signal_13524, new_AGEMA_signal_13523, new_AGEMA_signal_13522, MixColumnsIns_MixOneColumnInst_0_n40}), .c ({new_AGEMA_signal_14862, new_AGEMA_signal_14861, new_AGEMA_signal_14860, MixColumnsOutput[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U54 ( .a ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .b ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_13524, new_AGEMA_signal_13523, new_AGEMA_signal_13522, MixColumnsIns_MixOneColumnInst_0_n40}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U53 ( .a ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .b ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, new_AGEMA_signal_13543, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_14178, new_AGEMA_signal_14177, new_AGEMA_signal_14176, MixColumnsIns_MixOneColumnInst_0_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U52 ( .a ({new_AGEMA_signal_14181, new_AGEMA_signal_14180, new_AGEMA_signal_14179, MixColumnsIns_MixOneColumnInst_0_n18}), .b ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, new_AGEMA_signal_13525, MixColumnsIns_MixOneColumnInst_0_n35}), .c ({new_AGEMA_signal_14865, new_AGEMA_signal_14864, new_AGEMA_signal_14863, MixColumnsOutput[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U51 ( .a ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .b ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_13527, new_AGEMA_signal_13526, new_AGEMA_signal_13525, MixColumnsIns_MixOneColumnInst_0_n35}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U50 ( .a ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .b ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, new_AGEMA_signal_13549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_14181, new_AGEMA_signal_14180, new_AGEMA_signal_14179, MixColumnsIns_MixOneColumnInst_0_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U49 ( .a ({new_AGEMA_signal_14868, new_AGEMA_signal_14867, new_AGEMA_signal_14866, MixColumnsIns_MixOneColumnInst_0_n16}), .b ({new_AGEMA_signal_14184, new_AGEMA_signal_14183, new_AGEMA_signal_14182, MixColumnsIns_MixOneColumnInst_0_n33}), .c ({new_AGEMA_signal_15732, new_AGEMA_signal_15731, new_AGEMA_signal_15730, MixColumnsOutput[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U48 ( .a ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .b ({new_AGEMA_signal_13578, new_AGEMA_signal_13577, new_AGEMA_signal_13576, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}), .c ({new_AGEMA_signal_14184, new_AGEMA_signal_14183, new_AGEMA_signal_14182, MixColumnsIns_MixOneColumnInst_0_n33}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U47 ( .a ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .b ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, new_AGEMA_signal_14215, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_14868, new_AGEMA_signal_14867, new_AGEMA_signal_14866, MixColumnsIns_MixOneColumnInst_0_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U46 ( .a ({new_AGEMA_signal_14871, new_AGEMA_signal_14870, new_AGEMA_signal_14869, MixColumnsIns_MixOneColumnInst_0_n14}), .b ({new_AGEMA_signal_14187, new_AGEMA_signal_14186, new_AGEMA_signal_14185, MixColumnsIns_MixOneColumnInst_0_n27}), .c ({new_AGEMA_signal_15735, new_AGEMA_signal_15734, new_AGEMA_signal_15733, MixColumnsOutput[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U45 ( .a ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .b ({new_AGEMA_signal_13575, new_AGEMA_signal_13574, new_AGEMA_signal_13573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}), .c ({new_AGEMA_signal_14187, new_AGEMA_signal_14186, new_AGEMA_signal_14185, MixColumnsIns_MixOneColumnInst_0_n27}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U44 ( .a ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .b ({new_AGEMA_signal_14190, new_AGEMA_signal_14189, new_AGEMA_signal_14188, MixColumnsIns_MixOneColumnInst_0_n62}), .c ({new_AGEMA_signal_14871, new_AGEMA_signal_14870, new_AGEMA_signal_14869, MixColumnsIns_MixOneColumnInst_0_n14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U43 ( .a ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .b ({new_AGEMA_signal_13602, new_AGEMA_signal_13601, new_AGEMA_signal_13600, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}), .c ({new_AGEMA_signal_14190, new_AGEMA_signal_14189, new_AGEMA_signal_14188, MixColumnsIns_MixOneColumnInst_0_n62}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U42 ( .a ({new_AGEMA_signal_14874, new_AGEMA_signal_14873, new_AGEMA_signal_14872, MixColumnsIns_MixOneColumnInst_0_n13}), .b ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, new_AGEMA_signal_14191, MixColumnsIns_MixOneColumnInst_0_n31}), .c ({new_AGEMA_signal_15738, new_AGEMA_signal_15737, new_AGEMA_signal_15736, MixColumnsOutput[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U41 ( .a ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .b ({new_AGEMA_signal_13581, new_AGEMA_signal_13580, new_AGEMA_signal_13579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}), .c ({new_AGEMA_signal_14193, new_AGEMA_signal_14192, new_AGEMA_signal_14191, MixColumnsIns_MixOneColumnInst_0_n31}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U40 ( .a ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .b ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, new_AGEMA_signal_14221, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_14874, new_AGEMA_signal_14873, new_AGEMA_signal_14872, MixColumnsIns_MixOneColumnInst_0_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U39 ( .a ({new_AGEMA_signal_14196, new_AGEMA_signal_14195, new_AGEMA_signal_14194, MixColumnsIns_MixOneColumnInst_0_n11}), .b ({new_AGEMA_signal_13530, new_AGEMA_signal_13529, new_AGEMA_signal_13528, MixColumnsIns_MixOneColumnInst_0_n29}), .c ({new_AGEMA_signal_14877, new_AGEMA_signal_14876, new_AGEMA_signal_14875, MixColumnsOutput[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U38 ( .a ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .b ({new_AGEMA_signal_13287, new_AGEMA_signal_13286, new_AGEMA_signal_13285, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[18]}), .c ({new_AGEMA_signal_13530, new_AGEMA_signal_13529, new_AGEMA_signal_13528, MixColumnsIns_MixOneColumnInst_0_n29}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U37 ( .a ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .b ({new_AGEMA_signal_13557, new_AGEMA_signal_13556, new_AGEMA_signal_13555, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_14196, new_AGEMA_signal_14195, new_AGEMA_signal_14194, MixColumnsIns_MixOneColumnInst_0_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U36 ( .a ({new_AGEMA_signal_14880, new_AGEMA_signal_14879, new_AGEMA_signal_14878, MixColumnsIns_MixOneColumnInst_0_n9}), .b ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, new_AGEMA_signal_14197, MixColumnsIns_MixOneColumnInst_0_n26}), .c ({new_AGEMA_signal_15741, new_AGEMA_signal_15740, new_AGEMA_signal_15739, MixColumnsOutput[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U35 ( .a ({new_AGEMA_signal_13584, new_AGEMA_signal_13583, new_AGEMA_signal_13582, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}), .b ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_14199, new_AGEMA_signal_14198, new_AGEMA_signal_14197, MixColumnsIns_MixOneColumnInst_0_n26}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U34 ( .a ({new_AGEMA_signal_14202, new_AGEMA_signal_14201, new_AGEMA_signal_14200, MixColumnsIns_MixOneColumnInst_0_n63}), .b ({new_AGEMA_signal_13392, new_AGEMA_signal_13391, new_AGEMA_signal_13390, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[26]}), .c ({new_AGEMA_signal_14880, new_AGEMA_signal_14879, new_AGEMA_signal_14878, MixColumnsIns_MixOneColumnInst_0_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U33 ( .a ({new_AGEMA_signal_13593, new_AGEMA_signal_13592, new_AGEMA_signal_13591, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}), .b ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .c ({new_AGEMA_signal_14202, new_AGEMA_signal_14201, new_AGEMA_signal_14200, MixColumnsIns_MixOneColumnInst_0_n63}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U32 ( .a ({new_AGEMA_signal_14205, new_AGEMA_signal_14204, new_AGEMA_signal_14203, MixColumnsIns_MixOneColumnInst_0_n8}), .b ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, new_AGEMA_signal_13531, MixColumnsIns_MixOneColumnInst_0_n24}), .c ({new_AGEMA_signal_14883, new_AGEMA_signal_14882, new_AGEMA_signal_14881, MixColumnsOutput[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U31 ( .a ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .b ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_13533, new_AGEMA_signal_13532, new_AGEMA_signal_13531, MixColumnsIns_MixOneColumnInst_0_n24}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U30 ( .a ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .b ({new_AGEMA_signal_13536, new_AGEMA_signal_13535, new_AGEMA_signal_13534, MixColumnsIns_MixOneColumnInst_0_n60}), .c ({new_AGEMA_signal_14205, new_AGEMA_signal_14204, new_AGEMA_signal_14203, MixColumnsIns_MixOneColumnInst_0_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U29 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .c ({new_AGEMA_signal_13536, new_AGEMA_signal_13535, new_AGEMA_signal_13534, MixColumnsIns_MixOneColumnInst_0_n60}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U28 ( .a ({new_AGEMA_signal_14208, new_AGEMA_signal_14207, new_AGEMA_signal_14206, MixColumnsIns_MixOneColumnInst_0_n7}), .b ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, new_AGEMA_signal_13537, MixColumnsIns_MixOneColumnInst_0_n21}), .c ({new_AGEMA_signal_14886, new_AGEMA_signal_14885, new_AGEMA_signal_14884, MixColumnsOutput[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U27 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13167, new_AGEMA_signal_13166, new_AGEMA_signal_13165, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[15]}), .c ({new_AGEMA_signal_13539, new_AGEMA_signal_13538, new_AGEMA_signal_13537, MixColumnsIns_MixOneColumnInst_0_n21}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U26 ( .a ({new_AGEMA_signal_13542, new_AGEMA_signal_13541, new_AGEMA_signal_13540, MixColumnsIns_MixOneColumnInst_0_n56}), .b ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .c ({new_AGEMA_signal_14208, new_AGEMA_signal_14207, new_AGEMA_signal_14206, MixColumnsIns_MixOneColumnInst_0_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U25 ( .a ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_13542, new_AGEMA_signal_13541, new_AGEMA_signal_13540, MixColumnsIns_MixOneColumnInst_0_n56}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U24 ( .a ({new_AGEMA_signal_14211, new_AGEMA_signal_14210, new_AGEMA_signal_14209, MixColumnsIns_MixOneColumnInst_0_n6}), .b ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, new_AGEMA_signal_13543, MixColumnsIns_MixOneColumnInst_0_n19}), .c ({new_AGEMA_signal_14889, new_AGEMA_signal_14888, new_AGEMA_signal_14887, MixColumnsOutput[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U23 ( .a ({new_AGEMA_signal_13062, new_AGEMA_signal_13061, new_AGEMA_signal_13060, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[7]}), .b ({new_AGEMA_signal_13170, new_AGEMA_signal_13169, new_AGEMA_signal_13168, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[14]}), .c ({new_AGEMA_signal_13545, new_AGEMA_signal_13544, new_AGEMA_signal_13543, MixColumnsIns_MixOneColumnInst_0_n19}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U22 ( .a ({new_AGEMA_signal_13548, new_AGEMA_signal_13547, new_AGEMA_signal_13546, MixColumnsIns_MixOneColumnInst_0_n53}), .b ({new_AGEMA_signal_13272, new_AGEMA_signal_13271, new_AGEMA_signal_13270, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[23]}), .c ({new_AGEMA_signal_14211, new_AGEMA_signal_14210, new_AGEMA_signal_14209, MixColumnsIns_MixOneColumnInst_0_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U21 ( .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_13377, new_AGEMA_signal_13376, new_AGEMA_signal_13375, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[31]}), .c ({new_AGEMA_signal_13548, new_AGEMA_signal_13547, new_AGEMA_signal_13546, MixColumnsIns_MixOneColumnInst_0_n53}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U20 ( .a ({new_AGEMA_signal_14214, new_AGEMA_signal_14213, new_AGEMA_signal_14212, MixColumnsIns_MixOneColumnInst_0_n5}), .b ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, new_AGEMA_signal_13549, MixColumnsIns_MixOneColumnInst_0_n17}), .c ({new_AGEMA_signal_14892, new_AGEMA_signal_14891, new_AGEMA_signal_14890, MixColumnsOutput[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U19 ( .a ({new_AGEMA_signal_13065, new_AGEMA_signal_13064, new_AGEMA_signal_13063, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[6]}), .b ({new_AGEMA_signal_13173, new_AGEMA_signal_13172, new_AGEMA_signal_13171, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[13]}), .c ({new_AGEMA_signal_13551, new_AGEMA_signal_13550, new_AGEMA_signal_13549, MixColumnsIns_MixOneColumnInst_0_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U18 ( .a ({new_AGEMA_signal_13554, new_AGEMA_signal_13553, new_AGEMA_signal_13552, MixColumnsIns_MixOneColumnInst_0_n50}), .b ({new_AGEMA_signal_13275, new_AGEMA_signal_13274, new_AGEMA_signal_13273, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[22]}), .c ({new_AGEMA_signal_14214, new_AGEMA_signal_14213, new_AGEMA_signal_14212, MixColumnsIns_MixOneColumnInst_0_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U17 ( .a ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_13380, new_AGEMA_signal_13379, new_AGEMA_signal_13378, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[30]}), .c ({new_AGEMA_signal_13554, new_AGEMA_signal_13553, new_AGEMA_signal_13552, MixColumnsIns_MixOneColumnInst_0_n50}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U16 ( .a ({new_AGEMA_signal_14895, new_AGEMA_signal_14894, new_AGEMA_signal_14893, MixColumnsIns_MixOneColumnInst_0_n4}), .b ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, new_AGEMA_signal_14215, MixColumnsIns_MixOneColumnInst_0_n15}), .c ({new_AGEMA_signal_15744, new_AGEMA_signal_15743, new_AGEMA_signal_15742, MixColumnsOutput[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U15 ( .a ({new_AGEMA_signal_13068, new_AGEMA_signal_13067, new_AGEMA_signal_13066, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[5]}), .b ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, new_AGEMA_signal_13585, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}), .c ({new_AGEMA_signal_14217, new_AGEMA_signal_14216, new_AGEMA_signal_14215, MixColumnsIns_MixOneColumnInst_0_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U14 ( .a ({new_AGEMA_signal_14220, new_AGEMA_signal_14219, new_AGEMA_signal_14218, MixColumnsIns_MixOneColumnInst_0_n47}), .b ({new_AGEMA_signal_13278, new_AGEMA_signal_13277, new_AGEMA_signal_13276, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[21]}), .c ({new_AGEMA_signal_14895, new_AGEMA_signal_14894, new_AGEMA_signal_14893, MixColumnsIns_MixOneColumnInst_0_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U13 ( .a ({new_AGEMA_signal_13596, new_AGEMA_signal_13595, new_AGEMA_signal_13594, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}), .b ({new_AGEMA_signal_13383, new_AGEMA_signal_13382, new_AGEMA_signal_13381, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[29]}), .c ({new_AGEMA_signal_14220, new_AGEMA_signal_14219, new_AGEMA_signal_14218, MixColumnsIns_MixOneColumnInst_0_n47}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U12 ( .a ({new_AGEMA_signal_14898, new_AGEMA_signal_14897, new_AGEMA_signal_14896, MixColumnsIns_MixOneColumnInst_0_n3}), .b ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, new_AGEMA_signal_14221, MixColumnsIns_MixOneColumnInst_0_n12}), .c ({new_AGEMA_signal_15747, new_AGEMA_signal_15746, new_AGEMA_signal_15745, MixColumnsOutput[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U11 ( .a ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .b ({new_AGEMA_signal_13590, new_AGEMA_signal_13589, new_AGEMA_signal_13588, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}), .c ({new_AGEMA_signal_14223, new_AGEMA_signal_14222, new_AGEMA_signal_14221, MixColumnsIns_MixOneColumnInst_0_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U10 ( .a ({new_AGEMA_signal_14226, new_AGEMA_signal_14225, new_AGEMA_signal_14224, MixColumnsIns_MixOneColumnInst_0_n44}), .b ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .c ({new_AGEMA_signal_14898, new_AGEMA_signal_14897, new_AGEMA_signal_14896, MixColumnsIns_MixOneColumnInst_0_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U9 ( .a ({new_AGEMA_signal_13599, new_AGEMA_signal_13598, new_AGEMA_signal_13597, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .c ({new_AGEMA_signal_14226, new_AGEMA_signal_14225, new_AGEMA_signal_14224, MixColumnsIns_MixOneColumnInst_0_n44}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U8 ( .a ({new_AGEMA_signal_14229, new_AGEMA_signal_14228, new_AGEMA_signal_14227, MixColumnsIns_MixOneColumnInst_0_n2}), .b ({new_AGEMA_signal_13557, new_AGEMA_signal_13556, new_AGEMA_signal_13555, MixColumnsIns_MixOneColumnInst_0_n10}), .c ({new_AGEMA_signal_14901, new_AGEMA_signal_14900, new_AGEMA_signal_14899, MixColumnsOutput[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U7 ( .a ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .b ({new_AGEMA_signal_13182, new_AGEMA_signal_13181, new_AGEMA_signal_13180, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[10]}), .c ({new_AGEMA_signal_13557, new_AGEMA_signal_13556, new_AGEMA_signal_13555, MixColumnsIns_MixOneColumnInst_0_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U6 ( .a ({new_AGEMA_signal_13560, new_AGEMA_signal_13559, new_AGEMA_signal_13558, MixColumnsIns_MixOneColumnInst_0_n37}), .b ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .c ({new_AGEMA_signal_14229, new_AGEMA_signal_14228, new_AGEMA_signal_14227, MixColumnsIns_MixOneColumnInst_0_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U5 ( .a ({new_AGEMA_signal_13077, new_AGEMA_signal_13076, new_AGEMA_signal_13075, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[2]}), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .c ({new_AGEMA_signal_13560, new_AGEMA_signal_13559, new_AGEMA_signal_13558, MixColumnsIns_MixOneColumnInst_0_n37}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U4 ( .a ({new_AGEMA_signal_14232, new_AGEMA_signal_14231, new_AGEMA_signal_14230, MixColumnsIns_MixOneColumnInst_0_n1}), .b ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .c ({new_AGEMA_signal_14904, new_AGEMA_signal_14903, new_AGEMA_signal_14902, MixColumnsOutput[96]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U3 ( .a ({new_AGEMA_signal_13566, new_AGEMA_signal_13565, new_AGEMA_signal_13564, MixColumnsIns_MixOneColumnInst_0_n59}), .b ({new_AGEMA_signal_13563, new_AGEMA_signal_13562, new_AGEMA_signal_13561, MixColumnsIns_MixOneColumnInst_0_n23}), .c ({new_AGEMA_signal_14232, new_AGEMA_signal_14231, new_AGEMA_signal_14230, MixColumnsIns_MixOneColumnInst_0_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U2 ( .a ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .b ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .c ({new_AGEMA_signal_13563, new_AGEMA_signal_13562, new_AGEMA_signal_13561, MixColumnsIns_MixOneColumnInst_0_n23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_U1 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .c ({new_AGEMA_signal_13566, new_AGEMA_signal_13565, new_AGEMA_signal_13564, MixColumnsIns_MixOneColumnInst_0_n59}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_13386, new_AGEMA_signal_13385, new_AGEMA_signal_13384, MixColumnsInput[123]}), .c ({new_AGEMA_signal_13569, new_AGEMA_signal_13568, new_AGEMA_signal_13567, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_13389, new_AGEMA_signal_13388, new_AGEMA_signal_13387, MixColumnsInput[122]}), .c ({new_AGEMA_signal_13572, new_AGEMA_signal_13571, new_AGEMA_signal_13570, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13374, new_AGEMA_signal_13373, new_AGEMA_signal_13372, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[24]}), .b ({new_AGEMA_signal_12960, new_AGEMA_signal_12959, new_AGEMA_signal_12958, MixColumnsInput[120]}), .c ({new_AGEMA_signal_13575, new_AGEMA_signal_13574, new_AGEMA_signal_13573, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_13281, new_AGEMA_signal_13280, new_AGEMA_signal_13279, MixColumnsInput[115]}), .c ({new_AGEMA_signal_13578, new_AGEMA_signal_13577, new_AGEMA_signal_13576, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_13284, new_AGEMA_signal_13283, new_AGEMA_signal_13282, MixColumnsInput[114]}), .c ({new_AGEMA_signal_13581, new_AGEMA_signal_13580, new_AGEMA_signal_13579, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13269, new_AGEMA_signal_13268, new_AGEMA_signal_13267, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[16]}), .b ({new_AGEMA_signal_12795, new_AGEMA_signal_12794, new_AGEMA_signal_12793, MixColumnsInput[112]}), .c ({new_AGEMA_signal_13584, new_AGEMA_signal_13583, new_AGEMA_signal_13582, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_13176, new_AGEMA_signal_13175, new_AGEMA_signal_13174, MixColumnsInput[107]}), .c ({new_AGEMA_signal_13587, new_AGEMA_signal_13586, new_AGEMA_signal_13585, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_13179, new_AGEMA_signal_13178, new_AGEMA_signal_13177, MixColumnsInput[106]}), .c ({new_AGEMA_signal_13590, new_AGEMA_signal_13589, new_AGEMA_signal_13588, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13164, new_AGEMA_signal_13163, new_AGEMA_signal_13162, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[8]}), .b ({new_AGEMA_signal_12630, new_AGEMA_signal_12629, new_AGEMA_signal_12628, MixColumnsInput[104]}), .c ({new_AGEMA_signal_13593, new_AGEMA_signal_13592, new_AGEMA_signal_13591, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13071, new_AGEMA_signal_13070, new_AGEMA_signal_13069, MixColumnsInput[99]}), .c ({new_AGEMA_signal_13596, new_AGEMA_signal_13595, new_AGEMA_signal_13594, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_13074, new_AGEMA_signal_13073, new_AGEMA_signal_13072, MixColumnsInput[98]}), .c ({new_AGEMA_signal_13599, new_AGEMA_signal_13598, new_AGEMA_signal_13597, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_0_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13059, new_AGEMA_signal_13058, new_AGEMA_signal_13057, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[0]}), .b ({new_AGEMA_signal_12465, new_AGEMA_signal_12464, new_AGEMA_signal_12463, MixColumnsInput[96]}), .c ({new_AGEMA_signal_13602, new_AGEMA_signal_13601, new_AGEMA_signal_13600, MixColumnsIns_MixOneColumnInst_0_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U96 ( .a ({new_AGEMA_signal_14907, new_AGEMA_signal_14906, new_AGEMA_signal_14905, MixColumnsIns_MixOneColumnInst_1_n64}), .b ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_15750, new_AGEMA_signal_15749, new_AGEMA_signal_15748, MixColumnsOutput[73]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U95 ( .a ({new_AGEMA_signal_14298, new_AGEMA_signal_14297, new_AGEMA_signal_14296, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_14286, new_AGEMA_signal_14285, new_AGEMA_signal_14284, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_14907, new_AGEMA_signal_14906, new_AGEMA_signal_14905, MixColumnsIns_MixOneColumnInst_1_n64}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U94 ( .a ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, new_AGEMA_signal_14233, MixColumnsIns_MixOneColumnInst_1_n61}), .b ({new_AGEMA_signal_13632, new_AGEMA_signal_13631, new_AGEMA_signal_13630, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_14910, new_AGEMA_signal_14909, new_AGEMA_signal_14908, MixColumnsOutput[72]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U93 ( .a ({new_AGEMA_signal_13662, new_AGEMA_signal_13661, new_AGEMA_signal_13660, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .c ({new_AGEMA_signal_14235, new_AGEMA_signal_14234, new_AGEMA_signal_14233, MixColumnsIns_MixOneColumnInst_1_n61}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U92 ( .a ({new_AGEMA_signal_14238, new_AGEMA_signal_14237, new_AGEMA_signal_14236, MixColumnsIns_MixOneColumnInst_1_n58}), .b ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, new_AGEMA_signal_13603, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_14913, new_AGEMA_signal_14912, new_AGEMA_signal_14911, MixColumnsOutput[71]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U91 ( .a ({new_AGEMA_signal_13638, new_AGEMA_signal_13637, new_AGEMA_signal_13636, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .c ({new_AGEMA_signal_14238, new_AGEMA_signal_14237, new_AGEMA_signal_14236, MixColumnsIns_MixOneColumnInst_1_n58}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U90 ( .a ({new_AGEMA_signal_14241, new_AGEMA_signal_14240, new_AGEMA_signal_14239, MixColumnsIns_MixOneColumnInst_1_n55}), .b ({new_AGEMA_signal_13608, new_AGEMA_signal_13607, new_AGEMA_signal_13606, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_14916, new_AGEMA_signal_14915, new_AGEMA_signal_14914, MixColumnsOutput[70]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U89 ( .a ({new_AGEMA_signal_13644, new_AGEMA_signal_13643, new_AGEMA_signal_13642, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_14241, new_AGEMA_signal_14240, new_AGEMA_signal_14239, MixColumnsIns_MixOneColumnInst_1_n55}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U88 ( .a ({new_AGEMA_signal_14244, new_AGEMA_signal_14243, new_AGEMA_signal_14242, MixColumnsIns_MixOneColumnInst_1_n52}), .b ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, new_AGEMA_signal_13609, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_14919, new_AGEMA_signal_14918, new_AGEMA_signal_14917, MixColumnsOutput[69]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U87 ( .a ({new_AGEMA_signal_13650, new_AGEMA_signal_13649, new_AGEMA_signal_13648, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_14244, new_AGEMA_signal_14243, new_AGEMA_signal_14242, MixColumnsIns_MixOneColumnInst_1_n52}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U86 ( .a ({new_AGEMA_signal_14922, new_AGEMA_signal_14921, new_AGEMA_signal_14920, MixColumnsIns_MixOneColumnInst_1_n49}), .b ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, new_AGEMA_signal_14257, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_15753, new_AGEMA_signal_15752, new_AGEMA_signal_15751, MixColumnsOutput[68]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U85 ( .a ({new_AGEMA_signal_14316, new_AGEMA_signal_14315, new_AGEMA_signal_14314, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_14922, new_AGEMA_signal_14921, new_AGEMA_signal_14920, MixColumnsIns_MixOneColumnInst_1_n49}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U84 ( .a ({new_AGEMA_signal_14925, new_AGEMA_signal_14924, new_AGEMA_signal_14923, MixColumnsIns_MixOneColumnInst_1_n46}), .b ({new_AGEMA_signal_14262, new_AGEMA_signal_14261, new_AGEMA_signal_14260, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_15756, new_AGEMA_signal_15755, new_AGEMA_signal_15754, MixColumnsOutput[67]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U83 ( .a ({new_AGEMA_signal_14322, new_AGEMA_signal_14321, new_AGEMA_signal_14320, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .c ({new_AGEMA_signal_14925, new_AGEMA_signal_14924, new_AGEMA_signal_14923, MixColumnsIns_MixOneColumnInst_1_n46}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U82 ( .a ({new_AGEMA_signal_14247, new_AGEMA_signal_14246, new_AGEMA_signal_14245, MixColumnsIns_MixOneColumnInst_1_n43}), .b ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, new_AGEMA_signal_13603, MixColumnsIns_MixOneColumnInst_1_n57}), .c ({new_AGEMA_signal_14928, new_AGEMA_signal_14927, new_AGEMA_signal_14926, MixColumnsOutput[95]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U81 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_13605, new_AGEMA_signal_13604, new_AGEMA_signal_13603, MixColumnsIns_MixOneColumnInst_1_n57}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U80 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, new_AGEMA_signal_13615, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_14247, new_AGEMA_signal_14246, new_AGEMA_signal_14245, MixColumnsIns_MixOneColumnInst_1_n43}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U79 ( .a ({new_AGEMA_signal_14250, new_AGEMA_signal_14249, new_AGEMA_signal_14248, MixColumnsIns_MixOneColumnInst_1_n41}), .b ({new_AGEMA_signal_13608, new_AGEMA_signal_13607, new_AGEMA_signal_13606, MixColumnsIns_MixOneColumnInst_1_n54}), .c ({new_AGEMA_signal_14931, new_AGEMA_signal_14930, new_AGEMA_signal_14929, MixColumnsOutput[94]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U78 ( .a ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .b ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_13608, new_AGEMA_signal_13607, new_AGEMA_signal_13606, MixColumnsIns_MixOneColumnInst_1_n54}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U77 ( .a ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_13620, new_AGEMA_signal_13619, new_AGEMA_signal_13618, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_14250, new_AGEMA_signal_14249, new_AGEMA_signal_14248, MixColumnsIns_MixOneColumnInst_1_n41}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U76 ( .a ({new_AGEMA_signal_14253, new_AGEMA_signal_14252, new_AGEMA_signal_14251, MixColumnsIns_MixOneColumnInst_1_n39}), .b ({new_AGEMA_signal_13614, new_AGEMA_signal_13613, new_AGEMA_signal_13612, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_14934, new_AGEMA_signal_14933, new_AGEMA_signal_14932, MixColumnsOutput[66]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U75 ( .a ({new_AGEMA_signal_13656, new_AGEMA_signal_13655, new_AGEMA_signal_13654, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .c ({new_AGEMA_signal_14253, new_AGEMA_signal_14252, new_AGEMA_signal_14251, MixColumnsIns_MixOneColumnInst_1_n39}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U74 ( .a ({new_AGEMA_signal_14256, new_AGEMA_signal_14255, new_AGEMA_signal_14254, MixColumnsIns_MixOneColumnInst_1_n36}), .b ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, new_AGEMA_signal_13609, MixColumnsIns_MixOneColumnInst_1_n51}), .c ({new_AGEMA_signal_14937, new_AGEMA_signal_14936, new_AGEMA_signal_14935, MixColumnsOutput[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U73 ( .a ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_13611, new_AGEMA_signal_13610, new_AGEMA_signal_13609, MixColumnsIns_MixOneColumnInst_1_n51}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U72 ( .a ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, new_AGEMA_signal_13621, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_14256, new_AGEMA_signal_14255, new_AGEMA_signal_14254, MixColumnsIns_MixOneColumnInst_1_n36}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U71 ( .a ({new_AGEMA_signal_14940, new_AGEMA_signal_14939, new_AGEMA_signal_14938, MixColumnsIns_MixOneColumnInst_1_n34}), .b ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, new_AGEMA_signal_14257, MixColumnsIns_MixOneColumnInst_1_n48}), .c ({new_AGEMA_signal_15759, new_AGEMA_signal_15758, new_AGEMA_signal_15757, MixColumnsOutput[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U70 ( .a ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .b ({new_AGEMA_signal_13665, new_AGEMA_signal_13664, new_AGEMA_signal_13663, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}), .c ({new_AGEMA_signal_14259, new_AGEMA_signal_14258, new_AGEMA_signal_14257, MixColumnsIns_MixOneColumnInst_1_n48}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U69 ( .a ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_14280, new_AGEMA_signal_14279, new_AGEMA_signal_14278, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_14940, new_AGEMA_signal_14939, new_AGEMA_signal_14938, MixColumnsIns_MixOneColumnInst_1_n34}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U68 ( .a ({new_AGEMA_signal_14943, new_AGEMA_signal_14942, new_AGEMA_signal_14941, MixColumnsIns_MixOneColumnInst_1_n32}), .b ({new_AGEMA_signal_14262, new_AGEMA_signal_14261, new_AGEMA_signal_14260, MixColumnsIns_MixOneColumnInst_1_n45}), .c ({new_AGEMA_signal_15762, new_AGEMA_signal_15761, new_AGEMA_signal_15760, MixColumnsOutput[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U67 ( .a ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .b ({new_AGEMA_signal_13668, new_AGEMA_signal_13667, new_AGEMA_signal_13666, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}), .c ({new_AGEMA_signal_14262, new_AGEMA_signal_14261, new_AGEMA_signal_14260, MixColumnsIns_MixOneColumnInst_1_n45}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U66 ( .a ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .b ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, new_AGEMA_signal_14287, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_14943, new_AGEMA_signal_14942, new_AGEMA_signal_14941, MixColumnsIns_MixOneColumnInst_1_n32}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U65 ( .a ({new_AGEMA_signal_14265, new_AGEMA_signal_14264, new_AGEMA_signal_14263, MixColumnsIns_MixOneColumnInst_1_n30}), .b ({new_AGEMA_signal_13614, new_AGEMA_signal_13613, new_AGEMA_signal_13612, MixColumnsIns_MixOneColumnInst_1_n38}), .c ({new_AGEMA_signal_14946, new_AGEMA_signal_14945, new_AGEMA_signal_14944, MixColumnsOutput[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U64 ( .a ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .b ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_13614, new_AGEMA_signal_13613, new_AGEMA_signal_13612, MixColumnsIns_MixOneColumnInst_1_n38}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U63 ( .a ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .b ({new_AGEMA_signal_13626, new_AGEMA_signal_13625, new_AGEMA_signal_13624, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_14265, new_AGEMA_signal_14264, new_AGEMA_signal_14263, MixColumnsIns_MixOneColumnInst_1_n30}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U62 ( .a ({new_AGEMA_signal_14949, new_AGEMA_signal_14948, new_AGEMA_signal_14947, MixColumnsIns_MixOneColumnInst_1_n28}), .b ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, new_AGEMA_signal_14281, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_15765, new_AGEMA_signal_15764, new_AGEMA_signal_15763, MixColumnsOutput[89]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U61 ( .a ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, new_AGEMA_signal_14293, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_14949, new_AGEMA_signal_14948, new_AGEMA_signal_14947, MixColumnsIns_MixOneColumnInst_1_n28}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U60 ( .a ({new_AGEMA_signal_14268, new_AGEMA_signal_14267, new_AGEMA_signal_14266, MixColumnsIns_MixOneColumnInst_1_n25}), .b ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, new_AGEMA_signal_13627, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_14952, new_AGEMA_signal_14951, new_AGEMA_signal_14950, MixColumnsOutput[88]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U59 ( .a ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, new_AGEMA_signal_13657, MixColumnsIns_MixOneColumnInst_1_n23}), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .c ({new_AGEMA_signal_14268, new_AGEMA_signal_14267, new_AGEMA_signal_14266, MixColumnsIns_MixOneColumnInst_1_n25}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U58 ( .a ({new_AGEMA_signal_14271, new_AGEMA_signal_14270, new_AGEMA_signal_14269, MixColumnsIns_MixOneColumnInst_1_n22}), .b ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, new_AGEMA_signal_13615, MixColumnsIns_MixOneColumnInst_1_n42}), .c ({new_AGEMA_signal_14955, new_AGEMA_signal_14954, new_AGEMA_signal_14953, MixColumnsOutput[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U57 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_13617, new_AGEMA_signal_13616, new_AGEMA_signal_13615, MixColumnsIns_MixOneColumnInst_1_n42}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U56 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, new_AGEMA_signal_13633, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_14271, new_AGEMA_signal_14270, new_AGEMA_signal_14269, MixColumnsIns_MixOneColumnInst_1_n22}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U55 ( .a ({new_AGEMA_signal_14274, new_AGEMA_signal_14273, new_AGEMA_signal_14272, MixColumnsIns_MixOneColumnInst_1_n20}), .b ({new_AGEMA_signal_13620, new_AGEMA_signal_13619, new_AGEMA_signal_13618, MixColumnsIns_MixOneColumnInst_1_n40}), .c ({new_AGEMA_signal_14958, new_AGEMA_signal_14957, new_AGEMA_signal_14956, MixColumnsOutput[86]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U54 ( .a ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .b ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_13620, new_AGEMA_signal_13619, new_AGEMA_signal_13618, MixColumnsIns_MixOneColumnInst_1_n40}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U53 ( .a ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .b ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, new_AGEMA_signal_13639, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_14274, new_AGEMA_signal_14273, new_AGEMA_signal_14272, MixColumnsIns_MixOneColumnInst_1_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U52 ( .a ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, new_AGEMA_signal_14275, MixColumnsIns_MixOneColumnInst_1_n18}), .b ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, new_AGEMA_signal_13621, MixColumnsIns_MixOneColumnInst_1_n35}), .c ({new_AGEMA_signal_14961, new_AGEMA_signal_14960, new_AGEMA_signal_14959, MixColumnsOutput[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U51 ( .a ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_13623, new_AGEMA_signal_13622, new_AGEMA_signal_13621, MixColumnsIns_MixOneColumnInst_1_n35}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U50 ( .a ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .b ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, new_AGEMA_signal_13645, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_14277, new_AGEMA_signal_14276, new_AGEMA_signal_14275, MixColumnsIns_MixOneColumnInst_1_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U49 ( .a ({new_AGEMA_signal_14964, new_AGEMA_signal_14963, new_AGEMA_signal_14962, MixColumnsIns_MixOneColumnInst_1_n16}), .b ({new_AGEMA_signal_14280, new_AGEMA_signal_14279, new_AGEMA_signal_14278, MixColumnsIns_MixOneColumnInst_1_n33}), .c ({new_AGEMA_signal_15768, new_AGEMA_signal_15767, new_AGEMA_signal_15766, MixColumnsOutput[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U48 ( .a ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .b ({new_AGEMA_signal_13674, new_AGEMA_signal_13673, new_AGEMA_signal_13672, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}), .c ({new_AGEMA_signal_14280, new_AGEMA_signal_14279, new_AGEMA_signal_14278, MixColumnsIns_MixOneColumnInst_1_n33}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U47 ( .a ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .b ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, new_AGEMA_signal_14311, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_14964, new_AGEMA_signal_14963, new_AGEMA_signal_14962, MixColumnsIns_MixOneColumnInst_1_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U46 ( .a ({new_AGEMA_signal_14967, new_AGEMA_signal_14966, new_AGEMA_signal_14965, MixColumnsIns_MixOneColumnInst_1_n14}), .b ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, new_AGEMA_signal_14281, MixColumnsIns_MixOneColumnInst_1_n27}), .c ({new_AGEMA_signal_15771, new_AGEMA_signal_15770, new_AGEMA_signal_15769, MixColumnsOutput[65]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U45 ( .a ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .b ({new_AGEMA_signal_13671, new_AGEMA_signal_13670, new_AGEMA_signal_13669, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}), .c ({new_AGEMA_signal_14283, new_AGEMA_signal_14282, new_AGEMA_signal_14281, MixColumnsIns_MixOneColumnInst_1_n27}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U44 ( .a ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .b ({new_AGEMA_signal_14286, new_AGEMA_signal_14285, new_AGEMA_signal_14284, MixColumnsIns_MixOneColumnInst_1_n62}), .c ({new_AGEMA_signal_14967, new_AGEMA_signal_14966, new_AGEMA_signal_14965, MixColumnsIns_MixOneColumnInst_1_n14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U43 ( .a ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .b ({new_AGEMA_signal_13698, new_AGEMA_signal_13697, new_AGEMA_signal_13696, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}), .c ({new_AGEMA_signal_14286, new_AGEMA_signal_14285, new_AGEMA_signal_14284, MixColumnsIns_MixOneColumnInst_1_n62}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U42 ( .a ({new_AGEMA_signal_14970, new_AGEMA_signal_14969, new_AGEMA_signal_14968, MixColumnsIns_MixOneColumnInst_1_n13}), .b ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, new_AGEMA_signal_14287, MixColumnsIns_MixOneColumnInst_1_n31}), .c ({new_AGEMA_signal_15774, new_AGEMA_signal_15773, new_AGEMA_signal_15772, MixColumnsOutput[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U41 ( .a ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .b ({new_AGEMA_signal_13677, new_AGEMA_signal_13676, new_AGEMA_signal_13675, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}), .c ({new_AGEMA_signal_14289, new_AGEMA_signal_14288, new_AGEMA_signal_14287, MixColumnsIns_MixOneColumnInst_1_n31}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U40 ( .a ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .b ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, new_AGEMA_signal_14317, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_14970, new_AGEMA_signal_14969, new_AGEMA_signal_14968, MixColumnsIns_MixOneColumnInst_1_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U39 ( .a ({new_AGEMA_signal_14292, new_AGEMA_signal_14291, new_AGEMA_signal_14290, MixColumnsIns_MixOneColumnInst_1_n11}), .b ({new_AGEMA_signal_13626, new_AGEMA_signal_13625, new_AGEMA_signal_13624, MixColumnsIns_MixOneColumnInst_1_n29}), .c ({new_AGEMA_signal_14973, new_AGEMA_signal_14972, new_AGEMA_signal_14971, MixColumnsOutput[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U38 ( .a ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .b ({new_AGEMA_signal_13203, new_AGEMA_signal_13202, new_AGEMA_signal_13201, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[18]}), .c ({new_AGEMA_signal_13626, new_AGEMA_signal_13625, new_AGEMA_signal_13624, MixColumnsIns_MixOneColumnInst_1_n29}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U37 ( .a ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .b ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, new_AGEMA_signal_13651, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_14292, new_AGEMA_signal_14291, new_AGEMA_signal_14290, MixColumnsIns_MixOneColumnInst_1_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U36 ( .a ({new_AGEMA_signal_14976, new_AGEMA_signal_14975, new_AGEMA_signal_14974, MixColumnsIns_MixOneColumnInst_1_n9}), .b ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, new_AGEMA_signal_14293, MixColumnsIns_MixOneColumnInst_1_n26}), .c ({new_AGEMA_signal_15777, new_AGEMA_signal_15776, new_AGEMA_signal_15775, MixColumnsOutput[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U35 ( .a ({new_AGEMA_signal_13680, new_AGEMA_signal_13679, new_AGEMA_signal_13678, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}), .b ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_14295, new_AGEMA_signal_14294, new_AGEMA_signal_14293, MixColumnsIns_MixOneColumnInst_1_n26}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U34 ( .a ({new_AGEMA_signal_14298, new_AGEMA_signal_14297, new_AGEMA_signal_14296, MixColumnsIns_MixOneColumnInst_1_n63}), .b ({new_AGEMA_signal_13308, new_AGEMA_signal_13307, new_AGEMA_signal_13306, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[26]}), .c ({new_AGEMA_signal_14976, new_AGEMA_signal_14975, new_AGEMA_signal_14974, MixColumnsIns_MixOneColumnInst_1_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U33 ( .a ({new_AGEMA_signal_13689, new_AGEMA_signal_13688, new_AGEMA_signal_13687, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}), .b ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .c ({new_AGEMA_signal_14298, new_AGEMA_signal_14297, new_AGEMA_signal_14296, MixColumnsIns_MixOneColumnInst_1_n63}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U32 ( .a ({new_AGEMA_signal_14301, new_AGEMA_signal_14300, new_AGEMA_signal_14299, MixColumnsIns_MixOneColumnInst_1_n8}), .b ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, new_AGEMA_signal_13627, MixColumnsIns_MixOneColumnInst_1_n24}), .c ({new_AGEMA_signal_14979, new_AGEMA_signal_14978, new_AGEMA_signal_14977, MixColumnsOutput[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U31 ( .a ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_13629, new_AGEMA_signal_13628, new_AGEMA_signal_13627, MixColumnsIns_MixOneColumnInst_1_n24}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U30 ( .a ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .b ({new_AGEMA_signal_13632, new_AGEMA_signal_13631, new_AGEMA_signal_13630, MixColumnsIns_MixOneColumnInst_1_n60}), .c ({new_AGEMA_signal_14301, new_AGEMA_signal_14300, new_AGEMA_signal_14299, MixColumnsIns_MixOneColumnInst_1_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U29 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .c ({new_AGEMA_signal_13632, new_AGEMA_signal_13631, new_AGEMA_signal_13630, MixColumnsIns_MixOneColumnInst_1_n60}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U28 ( .a ({new_AGEMA_signal_14304, new_AGEMA_signal_14303, new_AGEMA_signal_14302, MixColumnsIns_MixOneColumnInst_1_n7}), .b ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, new_AGEMA_signal_13633, MixColumnsIns_MixOneColumnInst_1_n21}), .c ({new_AGEMA_signal_14982, new_AGEMA_signal_14981, new_AGEMA_signal_14980, MixColumnsOutput[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U27 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13083, new_AGEMA_signal_13082, new_AGEMA_signal_13081, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[15]}), .c ({new_AGEMA_signal_13635, new_AGEMA_signal_13634, new_AGEMA_signal_13633, MixColumnsIns_MixOneColumnInst_1_n21}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U26 ( .a ({new_AGEMA_signal_13638, new_AGEMA_signal_13637, new_AGEMA_signal_13636, MixColumnsIns_MixOneColumnInst_1_n56}), .b ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .c ({new_AGEMA_signal_14304, new_AGEMA_signal_14303, new_AGEMA_signal_14302, MixColumnsIns_MixOneColumnInst_1_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U25 ( .a ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_13638, new_AGEMA_signal_13637, new_AGEMA_signal_13636, MixColumnsIns_MixOneColumnInst_1_n56}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U24 ( .a ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, new_AGEMA_signal_14305, MixColumnsIns_MixOneColumnInst_1_n6}), .b ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, new_AGEMA_signal_13639, MixColumnsIns_MixOneColumnInst_1_n19}), .c ({new_AGEMA_signal_14985, new_AGEMA_signal_14984, new_AGEMA_signal_14983, MixColumnsOutput[78]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U23 ( .a ({new_AGEMA_signal_13314, new_AGEMA_signal_13313, new_AGEMA_signal_13312, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[7]}), .b ({new_AGEMA_signal_13086, new_AGEMA_signal_13085, new_AGEMA_signal_13084, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[14]}), .c ({new_AGEMA_signal_13641, new_AGEMA_signal_13640, new_AGEMA_signal_13639, MixColumnsIns_MixOneColumnInst_1_n19}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U22 ( .a ({new_AGEMA_signal_13644, new_AGEMA_signal_13643, new_AGEMA_signal_13642, MixColumnsIns_MixOneColumnInst_1_n53}), .b ({new_AGEMA_signal_13188, new_AGEMA_signal_13187, new_AGEMA_signal_13186, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[23]}), .c ({new_AGEMA_signal_14307, new_AGEMA_signal_14306, new_AGEMA_signal_14305, MixColumnsIns_MixOneColumnInst_1_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U21 ( .a ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_13293, new_AGEMA_signal_13292, new_AGEMA_signal_13291, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[31]}), .c ({new_AGEMA_signal_13644, new_AGEMA_signal_13643, new_AGEMA_signal_13642, MixColumnsIns_MixOneColumnInst_1_n53}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U20 ( .a ({new_AGEMA_signal_14310, new_AGEMA_signal_14309, new_AGEMA_signal_14308, MixColumnsIns_MixOneColumnInst_1_n5}), .b ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, new_AGEMA_signal_13645, MixColumnsIns_MixOneColumnInst_1_n17}), .c ({new_AGEMA_signal_14988, new_AGEMA_signal_14987, new_AGEMA_signal_14986, MixColumnsOutput[77]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U19 ( .a ({new_AGEMA_signal_13317, new_AGEMA_signal_13316, new_AGEMA_signal_13315, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[6]}), .b ({new_AGEMA_signal_13089, new_AGEMA_signal_13088, new_AGEMA_signal_13087, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[13]}), .c ({new_AGEMA_signal_13647, new_AGEMA_signal_13646, new_AGEMA_signal_13645, MixColumnsIns_MixOneColumnInst_1_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U18 ( .a ({new_AGEMA_signal_13650, new_AGEMA_signal_13649, new_AGEMA_signal_13648, MixColumnsIns_MixOneColumnInst_1_n50}), .b ({new_AGEMA_signal_13191, new_AGEMA_signal_13190, new_AGEMA_signal_13189, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[22]}), .c ({new_AGEMA_signal_14310, new_AGEMA_signal_14309, new_AGEMA_signal_14308, MixColumnsIns_MixOneColumnInst_1_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U17 ( .a ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_13296, new_AGEMA_signal_13295, new_AGEMA_signal_13294, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[30]}), .c ({new_AGEMA_signal_13650, new_AGEMA_signal_13649, new_AGEMA_signal_13648, MixColumnsIns_MixOneColumnInst_1_n50}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U16 ( .a ({new_AGEMA_signal_14991, new_AGEMA_signal_14990, new_AGEMA_signal_14989, MixColumnsIns_MixOneColumnInst_1_n4}), .b ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, new_AGEMA_signal_14311, MixColumnsIns_MixOneColumnInst_1_n15}), .c ({new_AGEMA_signal_15780, new_AGEMA_signal_15779, new_AGEMA_signal_15778, MixColumnsOutput[76]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U15 ( .a ({new_AGEMA_signal_13320, new_AGEMA_signal_13319, new_AGEMA_signal_13318, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[5]}), .b ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, new_AGEMA_signal_13681, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}), .c ({new_AGEMA_signal_14313, new_AGEMA_signal_14312, new_AGEMA_signal_14311, MixColumnsIns_MixOneColumnInst_1_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U14 ( .a ({new_AGEMA_signal_14316, new_AGEMA_signal_14315, new_AGEMA_signal_14314, MixColumnsIns_MixOneColumnInst_1_n47}), .b ({new_AGEMA_signal_13194, new_AGEMA_signal_13193, new_AGEMA_signal_13192, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[21]}), .c ({new_AGEMA_signal_14991, new_AGEMA_signal_14990, new_AGEMA_signal_14989, MixColumnsIns_MixOneColumnInst_1_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U13 ( .a ({new_AGEMA_signal_13692, new_AGEMA_signal_13691, new_AGEMA_signal_13690, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}), .b ({new_AGEMA_signal_13299, new_AGEMA_signal_13298, new_AGEMA_signal_13297, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[29]}), .c ({new_AGEMA_signal_14316, new_AGEMA_signal_14315, new_AGEMA_signal_14314, MixColumnsIns_MixOneColumnInst_1_n47}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U12 ( .a ({new_AGEMA_signal_14994, new_AGEMA_signal_14993, new_AGEMA_signal_14992, MixColumnsIns_MixOneColumnInst_1_n3}), .b ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, new_AGEMA_signal_14317, MixColumnsIns_MixOneColumnInst_1_n12}), .c ({new_AGEMA_signal_15783, new_AGEMA_signal_15782, new_AGEMA_signal_15781, MixColumnsOutput[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U11 ( .a ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .b ({new_AGEMA_signal_13686, new_AGEMA_signal_13685, new_AGEMA_signal_13684, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}), .c ({new_AGEMA_signal_14319, new_AGEMA_signal_14318, new_AGEMA_signal_14317, MixColumnsIns_MixOneColumnInst_1_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U10 ( .a ({new_AGEMA_signal_14322, new_AGEMA_signal_14321, new_AGEMA_signal_14320, MixColumnsIns_MixOneColumnInst_1_n44}), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .c ({new_AGEMA_signal_14994, new_AGEMA_signal_14993, new_AGEMA_signal_14992, MixColumnsIns_MixOneColumnInst_1_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U9 ( .a ({new_AGEMA_signal_13695, new_AGEMA_signal_13694, new_AGEMA_signal_13693, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}), .b ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .c ({new_AGEMA_signal_14322, new_AGEMA_signal_14321, new_AGEMA_signal_14320, MixColumnsIns_MixOneColumnInst_1_n44}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U8 ( .a ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, new_AGEMA_signal_14323, MixColumnsIns_MixOneColumnInst_1_n2}), .b ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, new_AGEMA_signal_13651, MixColumnsIns_MixOneColumnInst_1_n10}), .c ({new_AGEMA_signal_14997, new_AGEMA_signal_14996, new_AGEMA_signal_14995, MixColumnsOutput[74]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U7 ( .a ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .b ({new_AGEMA_signal_13098, new_AGEMA_signal_13097, new_AGEMA_signal_13096, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[10]}), .c ({new_AGEMA_signal_13653, new_AGEMA_signal_13652, new_AGEMA_signal_13651, MixColumnsIns_MixOneColumnInst_1_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U6 ( .a ({new_AGEMA_signal_13656, new_AGEMA_signal_13655, new_AGEMA_signal_13654, MixColumnsIns_MixOneColumnInst_1_n37}), .b ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .c ({new_AGEMA_signal_14325, new_AGEMA_signal_14324, new_AGEMA_signal_14323, MixColumnsIns_MixOneColumnInst_1_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U5 ( .a ({new_AGEMA_signal_13329, new_AGEMA_signal_13328, new_AGEMA_signal_13327, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[2]}), .b ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .c ({new_AGEMA_signal_13656, new_AGEMA_signal_13655, new_AGEMA_signal_13654, MixColumnsIns_MixOneColumnInst_1_n37}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U4 ( .a ({new_AGEMA_signal_14328, new_AGEMA_signal_14327, new_AGEMA_signal_14326, MixColumnsIns_MixOneColumnInst_1_n1}), .b ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .c ({new_AGEMA_signal_15000, new_AGEMA_signal_14999, new_AGEMA_signal_14998, MixColumnsOutput[64]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U3 ( .a ({new_AGEMA_signal_13662, new_AGEMA_signal_13661, new_AGEMA_signal_13660, MixColumnsIns_MixOneColumnInst_1_n59}), .b ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, new_AGEMA_signal_13657, MixColumnsIns_MixOneColumnInst_1_n23}), .c ({new_AGEMA_signal_14328, new_AGEMA_signal_14327, new_AGEMA_signal_14326, MixColumnsIns_MixOneColumnInst_1_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U2 ( .a ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .b ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .c ({new_AGEMA_signal_13659, new_AGEMA_signal_13658, new_AGEMA_signal_13657, MixColumnsIns_MixOneColumnInst_1_n23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_U1 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .c ({new_AGEMA_signal_13662, new_AGEMA_signal_13661, new_AGEMA_signal_13660, MixColumnsIns_MixOneColumnInst_1_n59}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_13302, new_AGEMA_signal_13301, new_AGEMA_signal_13300, MixColumnsInput[91]}), .c ({new_AGEMA_signal_13665, new_AGEMA_signal_13664, new_AGEMA_signal_13663, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_13305, new_AGEMA_signal_13304, new_AGEMA_signal_13303, MixColumnsInput[90]}), .c ({new_AGEMA_signal_13668, new_AGEMA_signal_13667, new_AGEMA_signal_13666, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13290, new_AGEMA_signal_13289, new_AGEMA_signal_13288, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[24]}), .b ({new_AGEMA_signal_12828, new_AGEMA_signal_12827, new_AGEMA_signal_12826, MixColumnsInput[88]}), .c ({new_AGEMA_signal_13671, new_AGEMA_signal_13670, new_AGEMA_signal_13669, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_13197, new_AGEMA_signal_13196, new_AGEMA_signal_13195, MixColumnsInput[83]}), .c ({new_AGEMA_signal_13674, new_AGEMA_signal_13673, new_AGEMA_signal_13672, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_13200, new_AGEMA_signal_13199, new_AGEMA_signal_13198, MixColumnsInput[82]}), .c ({new_AGEMA_signal_13677, new_AGEMA_signal_13676, new_AGEMA_signal_13675, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13185, new_AGEMA_signal_13184, new_AGEMA_signal_13183, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[16]}), .b ({new_AGEMA_signal_12663, new_AGEMA_signal_12662, new_AGEMA_signal_12661, MixColumnsInput[80]}), .c ({new_AGEMA_signal_13680, new_AGEMA_signal_13679, new_AGEMA_signal_13678, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_13092, new_AGEMA_signal_13091, new_AGEMA_signal_13090, MixColumnsInput[75]}), .c ({new_AGEMA_signal_13683, new_AGEMA_signal_13682, new_AGEMA_signal_13681, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_13095, new_AGEMA_signal_13094, new_AGEMA_signal_13093, MixColumnsInput[74]}), .c ({new_AGEMA_signal_13686, new_AGEMA_signal_13685, new_AGEMA_signal_13684, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13080, new_AGEMA_signal_13079, new_AGEMA_signal_13078, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[8]}), .b ({new_AGEMA_signal_12498, new_AGEMA_signal_12497, new_AGEMA_signal_12496, MixColumnsInput[72]}), .c ({new_AGEMA_signal_13689, new_AGEMA_signal_13688, new_AGEMA_signal_13687, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13323, new_AGEMA_signal_13322, new_AGEMA_signal_13321, MixColumnsInput[67]}), .c ({new_AGEMA_signal_13692, new_AGEMA_signal_13691, new_AGEMA_signal_13690, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_13326, new_AGEMA_signal_13325, new_AGEMA_signal_13324, MixColumnsInput[66]}), .c ({new_AGEMA_signal_13695, new_AGEMA_signal_13694, new_AGEMA_signal_13693, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_1_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13311, new_AGEMA_signal_13310, new_AGEMA_signal_13309, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[0]}), .b ({new_AGEMA_signal_12861, new_AGEMA_signal_12860, new_AGEMA_signal_12859, MixColumnsInput[64]}), .c ({new_AGEMA_signal_13698, new_AGEMA_signal_13697, new_AGEMA_signal_13696, MixColumnsIns_MixOneColumnInst_1_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U96 ( .a ({new_AGEMA_signal_15003, new_AGEMA_signal_15002, new_AGEMA_signal_15001, MixColumnsIns_MixOneColumnInst_2_n64}), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_15786, new_AGEMA_signal_15785, new_AGEMA_signal_15784, MixColumnsOutput[41]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U95 ( .a ({new_AGEMA_signal_14394, new_AGEMA_signal_14393, new_AGEMA_signal_14392, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_14382, new_AGEMA_signal_14381, new_AGEMA_signal_14380, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_15003, new_AGEMA_signal_15002, new_AGEMA_signal_15001, MixColumnsIns_MixOneColumnInst_2_n64}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U94 ( .a ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, new_AGEMA_signal_14329, MixColumnsIns_MixOneColumnInst_2_n61}), .b ({new_AGEMA_signal_13728, new_AGEMA_signal_13727, new_AGEMA_signal_13726, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_15006, new_AGEMA_signal_15005, new_AGEMA_signal_15004, MixColumnsOutput[40]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U93 ( .a ({new_AGEMA_signal_13758, new_AGEMA_signal_13757, new_AGEMA_signal_13756, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .c ({new_AGEMA_signal_14331, new_AGEMA_signal_14330, new_AGEMA_signal_14329, MixColumnsIns_MixOneColumnInst_2_n61}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U92 ( .a ({new_AGEMA_signal_14334, new_AGEMA_signal_14333, new_AGEMA_signal_14332, MixColumnsIns_MixOneColumnInst_2_n58}), .b ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, new_AGEMA_signal_13699, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_15009, new_AGEMA_signal_15008, new_AGEMA_signal_15007, MixColumnsOutput[39]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U91 ( .a ({new_AGEMA_signal_13734, new_AGEMA_signal_13733, new_AGEMA_signal_13732, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .c ({new_AGEMA_signal_14334, new_AGEMA_signal_14333, new_AGEMA_signal_14332, MixColumnsIns_MixOneColumnInst_2_n58}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U90 ( .a ({new_AGEMA_signal_14337, new_AGEMA_signal_14336, new_AGEMA_signal_14335, MixColumnsIns_MixOneColumnInst_2_n55}), .b ({new_AGEMA_signal_13704, new_AGEMA_signal_13703, new_AGEMA_signal_13702, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_15012, new_AGEMA_signal_15011, new_AGEMA_signal_15010, MixColumnsOutput[38]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U89 ( .a ({new_AGEMA_signal_13740, new_AGEMA_signal_13739, new_AGEMA_signal_13738, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_14337, new_AGEMA_signal_14336, new_AGEMA_signal_14335, MixColumnsIns_MixOneColumnInst_2_n55}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U88 ( .a ({new_AGEMA_signal_14340, new_AGEMA_signal_14339, new_AGEMA_signal_14338, MixColumnsIns_MixOneColumnInst_2_n52}), .b ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, new_AGEMA_signal_13705, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_15015, new_AGEMA_signal_15014, new_AGEMA_signal_15013, MixColumnsOutput[37]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U87 ( .a ({new_AGEMA_signal_13746, new_AGEMA_signal_13745, new_AGEMA_signal_13744, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_14340, new_AGEMA_signal_14339, new_AGEMA_signal_14338, MixColumnsIns_MixOneColumnInst_2_n52}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U86 ( .a ({new_AGEMA_signal_15018, new_AGEMA_signal_15017, new_AGEMA_signal_15016, MixColumnsIns_MixOneColumnInst_2_n49}), .b ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, new_AGEMA_signal_14353, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_15789, new_AGEMA_signal_15788, new_AGEMA_signal_15787, MixColumnsOutput[36]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U85 ( .a ({new_AGEMA_signal_14412, new_AGEMA_signal_14411, new_AGEMA_signal_14410, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_15018, new_AGEMA_signal_15017, new_AGEMA_signal_15016, MixColumnsIns_MixOneColumnInst_2_n49}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U84 ( .a ({new_AGEMA_signal_15021, new_AGEMA_signal_15020, new_AGEMA_signal_15019, MixColumnsIns_MixOneColumnInst_2_n46}), .b ({new_AGEMA_signal_14358, new_AGEMA_signal_14357, new_AGEMA_signal_14356, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_15792, new_AGEMA_signal_15791, new_AGEMA_signal_15790, MixColumnsOutput[35]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U83 ( .a ({new_AGEMA_signal_14418, new_AGEMA_signal_14417, new_AGEMA_signal_14416, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .c ({new_AGEMA_signal_15021, new_AGEMA_signal_15020, new_AGEMA_signal_15019, MixColumnsIns_MixOneColumnInst_2_n46}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U82 ( .a ({new_AGEMA_signal_14343, new_AGEMA_signal_14342, new_AGEMA_signal_14341, MixColumnsIns_MixOneColumnInst_2_n43}), .b ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, new_AGEMA_signal_13699, MixColumnsIns_MixOneColumnInst_2_n57}), .c ({new_AGEMA_signal_15024, new_AGEMA_signal_15023, new_AGEMA_signal_15022, MixColumnsOutput[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U81 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_13701, new_AGEMA_signal_13700, new_AGEMA_signal_13699, MixColumnsIns_MixOneColumnInst_2_n57}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U80 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, new_AGEMA_signal_13711, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_14343, new_AGEMA_signal_14342, new_AGEMA_signal_14341, MixColumnsIns_MixOneColumnInst_2_n43}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U79 ( .a ({new_AGEMA_signal_14346, new_AGEMA_signal_14345, new_AGEMA_signal_14344, MixColumnsIns_MixOneColumnInst_2_n41}), .b ({new_AGEMA_signal_13704, new_AGEMA_signal_13703, new_AGEMA_signal_13702, MixColumnsIns_MixOneColumnInst_2_n54}), .c ({new_AGEMA_signal_15027, new_AGEMA_signal_15026, new_AGEMA_signal_15025, MixColumnsOutput[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U78 ( .a ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .b ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_13704, new_AGEMA_signal_13703, new_AGEMA_signal_13702, MixColumnsIns_MixOneColumnInst_2_n54}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U77 ( .a ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_13716, new_AGEMA_signal_13715, new_AGEMA_signal_13714, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_14346, new_AGEMA_signal_14345, new_AGEMA_signal_14344, MixColumnsIns_MixOneColumnInst_2_n41}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U76 ( .a ({new_AGEMA_signal_14349, new_AGEMA_signal_14348, new_AGEMA_signal_14347, MixColumnsIns_MixOneColumnInst_2_n39}), .b ({new_AGEMA_signal_13710, new_AGEMA_signal_13709, new_AGEMA_signal_13708, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_15030, new_AGEMA_signal_15029, new_AGEMA_signal_15028, MixColumnsOutput[34]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U75 ( .a ({new_AGEMA_signal_13752, new_AGEMA_signal_13751, new_AGEMA_signal_13750, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .c ({new_AGEMA_signal_14349, new_AGEMA_signal_14348, new_AGEMA_signal_14347, MixColumnsIns_MixOneColumnInst_2_n39}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U74 ( .a ({new_AGEMA_signal_14352, new_AGEMA_signal_14351, new_AGEMA_signal_14350, MixColumnsIns_MixOneColumnInst_2_n36}), .b ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, new_AGEMA_signal_13705, MixColumnsIns_MixOneColumnInst_2_n51}), .c ({new_AGEMA_signal_15033, new_AGEMA_signal_15032, new_AGEMA_signal_15031, MixColumnsOutput[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U73 ( .a ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_13707, new_AGEMA_signal_13706, new_AGEMA_signal_13705, MixColumnsIns_MixOneColumnInst_2_n51}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U72 ( .a ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, new_AGEMA_signal_13717, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_14352, new_AGEMA_signal_14351, new_AGEMA_signal_14350, MixColumnsIns_MixOneColumnInst_2_n36}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U71 ( .a ({new_AGEMA_signal_15036, new_AGEMA_signal_15035, new_AGEMA_signal_15034, MixColumnsIns_MixOneColumnInst_2_n34}), .b ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, new_AGEMA_signal_14353, MixColumnsIns_MixOneColumnInst_2_n48}), .c ({new_AGEMA_signal_15795, new_AGEMA_signal_15794, new_AGEMA_signal_15793, MixColumnsOutput[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U70 ( .a ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .b ({new_AGEMA_signal_13761, new_AGEMA_signal_13760, new_AGEMA_signal_13759, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}), .c ({new_AGEMA_signal_14355, new_AGEMA_signal_14354, new_AGEMA_signal_14353, MixColumnsIns_MixOneColumnInst_2_n48}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U69 ( .a ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_14376, new_AGEMA_signal_14375, new_AGEMA_signal_14374, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_15036, new_AGEMA_signal_15035, new_AGEMA_signal_15034, MixColumnsIns_MixOneColumnInst_2_n34}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U68 ( .a ({new_AGEMA_signal_15039, new_AGEMA_signal_15038, new_AGEMA_signal_15037, MixColumnsIns_MixOneColumnInst_2_n32}), .b ({new_AGEMA_signal_14358, new_AGEMA_signal_14357, new_AGEMA_signal_14356, MixColumnsIns_MixOneColumnInst_2_n45}), .c ({new_AGEMA_signal_15798, new_AGEMA_signal_15797, new_AGEMA_signal_15796, MixColumnsOutput[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U67 ( .a ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .b ({new_AGEMA_signal_13764, new_AGEMA_signal_13763, new_AGEMA_signal_13762, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}), .c ({new_AGEMA_signal_14358, new_AGEMA_signal_14357, new_AGEMA_signal_14356, MixColumnsIns_MixOneColumnInst_2_n45}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U66 ( .a ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .b ({new_AGEMA_signal_14385, new_AGEMA_signal_14384, new_AGEMA_signal_14383, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_15039, new_AGEMA_signal_15038, new_AGEMA_signal_15037, MixColumnsIns_MixOneColumnInst_2_n32}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U65 ( .a ({new_AGEMA_signal_14361, new_AGEMA_signal_14360, new_AGEMA_signal_14359, MixColumnsIns_MixOneColumnInst_2_n30}), .b ({new_AGEMA_signal_13710, new_AGEMA_signal_13709, new_AGEMA_signal_13708, MixColumnsIns_MixOneColumnInst_2_n38}), .c ({new_AGEMA_signal_15042, new_AGEMA_signal_15041, new_AGEMA_signal_15040, MixColumnsOutput[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U64 ( .a ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .b ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_13710, new_AGEMA_signal_13709, new_AGEMA_signal_13708, MixColumnsIns_MixOneColumnInst_2_n38}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U63 ( .a ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .b ({new_AGEMA_signal_13722, new_AGEMA_signal_13721, new_AGEMA_signal_13720, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_14361, new_AGEMA_signal_14360, new_AGEMA_signal_14359, MixColumnsIns_MixOneColumnInst_2_n30}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U62 ( .a ({new_AGEMA_signal_15045, new_AGEMA_signal_15044, new_AGEMA_signal_15043, MixColumnsIns_MixOneColumnInst_2_n28}), .b ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, new_AGEMA_signal_14377, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_15801, new_AGEMA_signal_15800, new_AGEMA_signal_15799, MixColumnsOutput[57]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U61 ( .a ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_14391, new_AGEMA_signal_14390, new_AGEMA_signal_14389, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_15045, new_AGEMA_signal_15044, new_AGEMA_signal_15043, MixColumnsIns_MixOneColumnInst_2_n28}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U60 ( .a ({new_AGEMA_signal_14364, new_AGEMA_signal_14363, new_AGEMA_signal_14362, MixColumnsIns_MixOneColumnInst_2_n25}), .b ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, new_AGEMA_signal_13723, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_15048, new_AGEMA_signal_15047, new_AGEMA_signal_15046, MixColumnsOutput[56]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U59 ( .a ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, new_AGEMA_signal_13753, MixColumnsIns_MixOneColumnInst_2_n23}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .c ({new_AGEMA_signal_14364, new_AGEMA_signal_14363, new_AGEMA_signal_14362, MixColumnsIns_MixOneColumnInst_2_n25}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U58 ( .a ({new_AGEMA_signal_14367, new_AGEMA_signal_14366, new_AGEMA_signal_14365, MixColumnsIns_MixOneColumnInst_2_n22}), .b ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, new_AGEMA_signal_13711, MixColumnsIns_MixOneColumnInst_2_n42}), .c ({new_AGEMA_signal_15051, new_AGEMA_signal_15050, new_AGEMA_signal_15049, MixColumnsOutput[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U57 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_13713, new_AGEMA_signal_13712, new_AGEMA_signal_13711, MixColumnsIns_MixOneColumnInst_2_n42}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U56 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, new_AGEMA_signal_13729, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_14367, new_AGEMA_signal_14366, new_AGEMA_signal_14365, MixColumnsIns_MixOneColumnInst_2_n22}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U55 ( .a ({new_AGEMA_signal_14370, new_AGEMA_signal_14369, new_AGEMA_signal_14368, MixColumnsIns_MixOneColumnInst_2_n20}), .b ({new_AGEMA_signal_13716, new_AGEMA_signal_13715, new_AGEMA_signal_13714, MixColumnsIns_MixOneColumnInst_2_n40}), .c ({new_AGEMA_signal_15054, new_AGEMA_signal_15053, new_AGEMA_signal_15052, MixColumnsOutput[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U54 ( .a ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_13716, new_AGEMA_signal_13715, new_AGEMA_signal_13714, MixColumnsIns_MixOneColumnInst_2_n40}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U53 ( .a ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .b ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, new_AGEMA_signal_13735, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_14370, new_AGEMA_signal_14369, new_AGEMA_signal_14368, MixColumnsIns_MixOneColumnInst_2_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U52 ( .a ({new_AGEMA_signal_14373, new_AGEMA_signal_14372, new_AGEMA_signal_14371, MixColumnsIns_MixOneColumnInst_2_n18}), .b ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, new_AGEMA_signal_13717, MixColumnsIns_MixOneColumnInst_2_n35}), .c ({new_AGEMA_signal_15057, new_AGEMA_signal_15056, new_AGEMA_signal_15055, MixColumnsOutput[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U51 ( .a ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .b ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_13719, new_AGEMA_signal_13718, new_AGEMA_signal_13717, MixColumnsIns_MixOneColumnInst_2_n35}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U50 ( .a ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .b ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, new_AGEMA_signal_13741, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_14373, new_AGEMA_signal_14372, new_AGEMA_signal_14371, MixColumnsIns_MixOneColumnInst_2_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U49 ( .a ({new_AGEMA_signal_15060, new_AGEMA_signal_15059, new_AGEMA_signal_15058, MixColumnsIns_MixOneColumnInst_2_n16}), .b ({new_AGEMA_signal_14376, new_AGEMA_signal_14375, new_AGEMA_signal_14374, MixColumnsIns_MixOneColumnInst_2_n33}), .c ({new_AGEMA_signal_15804, new_AGEMA_signal_15803, new_AGEMA_signal_15802, MixColumnsOutput[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U48 ( .a ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .b ({new_AGEMA_signal_13770, new_AGEMA_signal_13769, new_AGEMA_signal_13768, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}), .c ({new_AGEMA_signal_14376, new_AGEMA_signal_14375, new_AGEMA_signal_14374, MixColumnsIns_MixOneColumnInst_2_n33}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U47 ( .a ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .b ({new_AGEMA_signal_14409, new_AGEMA_signal_14408, new_AGEMA_signal_14407, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_15060, new_AGEMA_signal_15059, new_AGEMA_signal_15058, MixColumnsIns_MixOneColumnInst_2_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U46 ( .a ({new_AGEMA_signal_15063, new_AGEMA_signal_15062, new_AGEMA_signal_15061, MixColumnsIns_MixOneColumnInst_2_n14}), .b ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, new_AGEMA_signal_14377, MixColumnsIns_MixOneColumnInst_2_n27}), .c ({new_AGEMA_signal_15807, new_AGEMA_signal_15806, new_AGEMA_signal_15805, MixColumnsOutput[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U45 ( .a ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .b ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, new_AGEMA_signal_13765, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}), .c ({new_AGEMA_signal_14379, new_AGEMA_signal_14378, new_AGEMA_signal_14377, MixColumnsIns_MixOneColumnInst_2_n27}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U44 ( .a ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .b ({new_AGEMA_signal_14382, new_AGEMA_signal_14381, new_AGEMA_signal_14380, MixColumnsIns_MixOneColumnInst_2_n62}), .c ({new_AGEMA_signal_15063, new_AGEMA_signal_15062, new_AGEMA_signal_15061, MixColumnsIns_MixOneColumnInst_2_n14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U43 ( .a ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .b ({new_AGEMA_signal_13794, new_AGEMA_signal_13793, new_AGEMA_signal_13792, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}), .c ({new_AGEMA_signal_14382, new_AGEMA_signal_14381, new_AGEMA_signal_14380, MixColumnsIns_MixOneColumnInst_2_n62}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U42 ( .a ({new_AGEMA_signal_15066, new_AGEMA_signal_15065, new_AGEMA_signal_15064, MixColumnsIns_MixOneColumnInst_2_n13}), .b ({new_AGEMA_signal_14385, new_AGEMA_signal_14384, new_AGEMA_signal_14383, MixColumnsIns_MixOneColumnInst_2_n31}), .c ({new_AGEMA_signal_15810, new_AGEMA_signal_15809, new_AGEMA_signal_15808, MixColumnsOutput[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U41 ( .a ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .b ({new_AGEMA_signal_13773, new_AGEMA_signal_13772, new_AGEMA_signal_13771, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}), .c ({new_AGEMA_signal_14385, new_AGEMA_signal_14384, new_AGEMA_signal_14383, MixColumnsIns_MixOneColumnInst_2_n31}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U40 ( .a ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .b ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, new_AGEMA_signal_14413, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_15066, new_AGEMA_signal_15065, new_AGEMA_signal_15064, MixColumnsIns_MixOneColumnInst_2_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U39 ( .a ({new_AGEMA_signal_14388, new_AGEMA_signal_14387, new_AGEMA_signal_14386, MixColumnsIns_MixOneColumnInst_2_n11}), .b ({new_AGEMA_signal_13722, new_AGEMA_signal_13721, new_AGEMA_signal_13720, MixColumnsIns_MixOneColumnInst_2_n29}), .c ({new_AGEMA_signal_15069, new_AGEMA_signal_15068, new_AGEMA_signal_15067, MixColumnsOutput[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U38 ( .a ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .b ({new_AGEMA_signal_13119, new_AGEMA_signal_13118, new_AGEMA_signal_13117, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[18]}), .c ({new_AGEMA_signal_13722, new_AGEMA_signal_13721, new_AGEMA_signal_13720, MixColumnsIns_MixOneColumnInst_2_n29}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U37 ( .a ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .b ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, new_AGEMA_signal_13747, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_14388, new_AGEMA_signal_14387, new_AGEMA_signal_14386, MixColumnsIns_MixOneColumnInst_2_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U36 ( .a ({new_AGEMA_signal_15072, new_AGEMA_signal_15071, new_AGEMA_signal_15070, MixColumnsIns_MixOneColumnInst_2_n9}), .b ({new_AGEMA_signal_14391, new_AGEMA_signal_14390, new_AGEMA_signal_14389, MixColumnsIns_MixOneColumnInst_2_n26}), .c ({new_AGEMA_signal_15813, new_AGEMA_signal_15812, new_AGEMA_signal_15811, MixColumnsOutput[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U35 ( .a ({new_AGEMA_signal_13776, new_AGEMA_signal_13775, new_AGEMA_signal_13774, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}), .b ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_14391, new_AGEMA_signal_14390, new_AGEMA_signal_14389, MixColumnsIns_MixOneColumnInst_2_n26}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U34 ( .a ({new_AGEMA_signal_14394, new_AGEMA_signal_14393, new_AGEMA_signal_14392, MixColumnsIns_MixOneColumnInst_2_n63}), .b ({new_AGEMA_signal_13224, new_AGEMA_signal_13223, new_AGEMA_signal_13222, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[26]}), .c ({new_AGEMA_signal_15072, new_AGEMA_signal_15071, new_AGEMA_signal_15070, MixColumnsIns_MixOneColumnInst_2_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U33 ( .a ({new_AGEMA_signal_13785, new_AGEMA_signal_13784, new_AGEMA_signal_13783, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}), .b ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .c ({new_AGEMA_signal_14394, new_AGEMA_signal_14393, new_AGEMA_signal_14392, MixColumnsIns_MixOneColumnInst_2_n63}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U32 ( .a ({new_AGEMA_signal_14397, new_AGEMA_signal_14396, new_AGEMA_signal_14395, MixColumnsIns_MixOneColumnInst_2_n8}), .b ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, new_AGEMA_signal_13723, MixColumnsIns_MixOneColumnInst_2_n24}), .c ({new_AGEMA_signal_15075, new_AGEMA_signal_15074, new_AGEMA_signal_15073, MixColumnsOutput[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U31 ( .a ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_13725, new_AGEMA_signal_13724, new_AGEMA_signal_13723, MixColumnsIns_MixOneColumnInst_2_n24}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U30 ( .a ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .b ({new_AGEMA_signal_13728, new_AGEMA_signal_13727, new_AGEMA_signal_13726, MixColumnsIns_MixOneColumnInst_2_n60}), .c ({new_AGEMA_signal_14397, new_AGEMA_signal_14396, new_AGEMA_signal_14395, MixColumnsIns_MixOneColumnInst_2_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U29 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .c ({new_AGEMA_signal_13728, new_AGEMA_signal_13727, new_AGEMA_signal_13726, MixColumnsIns_MixOneColumnInst_2_n60}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U28 ( .a ({new_AGEMA_signal_14400, new_AGEMA_signal_14399, new_AGEMA_signal_14398, MixColumnsIns_MixOneColumnInst_2_n7}), .b ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, new_AGEMA_signal_13729, MixColumnsIns_MixOneColumnInst_2_n21}), .c ({new_AGEMA_signal_15078, new_AGEMA_signal_15077, new_AGEMA_signal_15076, MixColumnsOutput[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U27 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13335, new_AGEMA_signal_13334, new_AGEMA_signal_13333, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[15]}), .c ({new_AGEMA_signal_13731, new_AGEMA_signal_13730, new_AGEMA_signal_13729, MixColumnsIns_MixOneColumnInst_2_n21}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U26 ( .a ({new_AGEMA_signal_13734, new_AGEMA_signal_13733, new_AGEMA_signal_13732, MixColumnsIns_MixOneColumnInst_2_n56}), .b ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .c ({new_AGEMA_signal_14400, new_AGEMA_signal_14399, new_AGEMA_signal_14398, MixColumnsIns_MixOneColumnInst_2_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U25 ( .a ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_13734, new_AGEMA_signal_13733, new_AGEMA_signal_13732, MixColumnsIns_MixOneColumnInst_2_n56}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U24 ( .a ({new_AGEMA_signal_14403, new_AGEMA_signal_14402, new_AGEMA_signal_14401, MixColumnsIns_MixOneColumnInst_2_n6}), .b ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, new_AGEMA_signal_13735, MixColumnsIns_MixOneColumnInst_2_n19}), .c ({new_AGEMA_signal_15081, new_AGEMA_signal_15080, new_AGEMA_signal_15079, MixColumnsOutput[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U23 ( .a ({new_AGEMA_signal_13230, new_AGEMA_signal_13229, new_AGEMA_signal_13228, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[7]}), .b ({new_AGEMA_signal_13338, new_AGEMA_signal_13337, new_AGEMA_signal_13336, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[14]}), .c ({new_AGEMA_signal_13737, new_AGEMA_signal_13736, new_AGEMA_signal_13735, MixColumnsIns_MixOneColumnInst_2_n19}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U22 ( .a ({new_AGEMA_signal_13740, new_AGEMA_signal_13739, new_AGEMA_signal_13738, MixColumnsIns_MixOneColumnInst_2_n53}), .b ({new_AGEMA_signal_13104, new_AGEMA_signal_13103, new_AGEMA_signal_13102, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[23]}), .c ({new_AGEMA_signal_14403, new_AGEMA_signal_14402, new_AGEMA_signal_14401, MixColumnsIns_MixOneColumnInst_2_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U21 ( .a ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_13209, new_AGEMA_signal_13208, new_AGEMA_signal_13207, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[31]}), .c ({new_AGEMA_signal_13740, new_AGEMA_signal_13739, new_AGEMA_signal_13738, MixColumnsIns_MixOneColumnInst_2_n53}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U20 ( .a ({new_AGEMA_signal_14406, new_AGEMA_signal_14405, new_AGEMA_signal_14404, MixColumnsIns_MixOneColumnInst_2_n5}), .b ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, new_AGEMA_signal_13741, MixColumnsIns_MixOneColumnInst_2_n17}), .c ({new_AGEMA_signal_15084, new_AGEMA_signal_15083, new_AGEMA_signal_15082, MixColumnsOutput[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U19 ( .a ({new_AGEMA_signal_13233, new_AGEMA_signal_13232, new_AGEMA_signal_13231, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[6]}), .b ({new_AGEMA_signal_13341, new_AGEMA_signal_13340, new_AGEMA_signal_13339, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[13]}), .c ({new_AGEMA_signal_13743, new_AGEMA_signal_13742, new_AGEMA_signal_13741, MixColumnsIns_MixOneColumnInst_2_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U18 ( .a ({new_AGEMA_signal_13746, new_AGEMA_signal_13745, new_AGEMA_signal_13744, MixColumnsIns_MixOneColumnInst_2_n50}), .b ({new_AGEMA_signal_13107, new_AGEMA_signal_13106, new_AGEMA_signal_13105, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[22]}), .c ({new_AGEMA_signal_14406, new_AGEMA_signal_14405, new_AGEMA_signal_14404, MixColumnsIns_MixOneColumnInst_2_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U17 ( .a ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_13212, new_AGEMA_signal_13211, new_AGEMA_signal_13210, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[30]}), .c ({new_AGEMA_signal_13746, new_AGEMA_signal_13745, new_AGEMA_signal_13744, MixColumnsIns_MixOneColumnInst_2_n50}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U16 ( .a ({new_AGEMA_signal_15087, new_AGEMA_signal_15086, new_AGEMA_signal_15085, MixColumnsIns_MixOneColumnInst_2_n4}), .b ({new_AGEMA_signal_14409, new_AGEMA_signal_14408, new_AGEMA_signal_14407, MixColumnsIns_MixOneColumnInst_2_n15}), .c ({new_AGEMA_signal_15816, new_AGEMA_signal_15815, new_AGEMA_signal_15814, MixColumnsOutput[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U15 ( .a ({new_AGEMA_signal_13236, new_AGEMA_signal_13235, new_AGEMA_signal_13234, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[5]}), .b ({new_AGEMA_signal_13779, new_AGEMA_signal_13778, new_AGEMA_signal_13777, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}), .c ({new_AGEMA_signal_14409, new_AGEMA_signal_14408, new_AGEMA_signal_14407, MixColumnsIns_MixOneColumnInst_2_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U14 ( .a ({new_AGEMA_signal_14412, new_AGEMA_signal_14411, new_AGEMA_signal_14410, MixColumnsIns_MixOneColumnInst_2_n47}), .b ({new_AGEMA_signal_13110, new_AGEMA_signal_13109, new_AGEMA_signal_13108, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[21]}), .c ({new_AGEMA_signal_15087, new_AGEMA_signal_15086, new_AGEMA_signal_15085, MixColumnsIns_MixOneColumnInst_2_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U13 ( .a ({new_AGEMA_signal_13788, new_AGEMA_signal_13787, new_AGEMA_signal_13786, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}), .b ({new_AGEMA_signal_13215, new_AGEMA_signal_13214, new_AGEMA_signal_13213, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[29]}), .c ({new_AGEMA_signal_14412, new_AGEMA_signal_14411, new_AGEMA_signal_14410, MixColumnsIns_MixOneColumnInst_2_n47}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U12 ( .a ({new_AGEMA_signal_15090, new_AGEMA_signal_15089, new_AGEMA_signal_15088, MixColumnsIns_MixOneColumnInst_2_n3}), .b ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, new_AGEMA_signal_14413, MixColumnsIns_MixOneColumnInst_2_n12}), .c ({new_AGEMA_signal_15819, new_AGEMA_signal_15818, new_AGEMA_signal_15817, MixColumnsOutput[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U11 ( .a ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .b ({new_AGEMA_signal_13782, new_AGEMA_signal_13781, new_AGEMA_signal_13780, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}), .c ({new_AGEMA_signal_14415, new_AGEMA_signal_14414, new_AGEMA_signal_14413, MixColumnsIns_MixOneColumnInst_2_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U10 ( .a ({new_AGEMA_signal_14418, new_AGEMA_signal_14417, new_AGEMA_signal_14416, MixColumnsIns_MixOneColumnInst_2_n44}), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .c ({new_AGEMA_signal_15090, new_AGEMA_signal_15089, new_AGEMA_signal_15088, MixColumnsIns_MixOneColumnInst_2_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U9 ( .a ({new_AGEMA_signal_13791, new_AGEMA_signal_13790, new_AGEMA_signal_13789, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}), .b ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .c ({new_AGEMA_signal_14418, new_AGEMA_signal_14417, new_AGEMA_signal_14416, MixColumnsIns_MixOneColumnInst_2_n44}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U8 ( .a ({new_AGEMA_signal_14421, new_AGEMA_signal_14420, new_AGEMA_signal_14419, MixColumnsIns_MixOneColumnInst_2_n2}), .b ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, new_AGEMA_signal_13747, MixColumnsIns_MixOneColumnInst_2_n10}), .c ({new_AGEMA_signal_15093, new_AGEMA_signal_15092, new_AGEMA_signal_15091, MixColumnsOutput[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U7 ( .a ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .b ({new_AGEMA_signal_13350, new_AGEMA_signal_13349, new_AGEMA_signal_13348, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[10]}), .c ({new_AGEMA_signal_13749, new_AGEMA_signal_13748, new_AGEMA_signal_13747, MixColumnsIns_MixOneColumnInst_2_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U6 ( .a ({new_AGEMA_signal_13752, new_AGEMA_signal_13751, new_AGEMA_signal_13750, MixColumnsIns_MixOneColumnInst_2_n37}), .b ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .c ({new_AGEMA_signal_14421, new_AGEMA_signal_14420, new_AGEMA_signal_14419, MixColumnsIns_MixOneColumnInst_2_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U5 ( .a ({new_AGEMA_signal_13245, new_AGEMA_signal_13244, new_AGEMA_signal_13243, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[2]}), .b ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .c ({new_AGEMA_signal_13752, new_AGEMA_signal_13751, new_AGEMA_signal_13750, MixColumnsIns_MixOneColumnInst_2_n37}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U4 ( .a ({new_AGEMA_signal_14424, new_AGEMA_signal_14423, new_AGEMA_signal_14422, MixColumnsIns_MixOneColumnInst_2_n1}), .b ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .c ({new_AGEMA_signal_15096, new_AGEMA_signal_15095, new_AGEMA_signal_15094, MixColumnsOutput[32]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U3 ( .a ({new_AGEMA_signal_13758, new_AGEMA_signal_13757, new_AGEMA_signal_13756, MixColumnsIns_MixOneColumnInst_2_n59}), .b ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, new_AGEMA_signal_13753, MixColumnsIns_MixOneColumnInst_2_n23}), .c ({new_AGEMA_signal_14424, new_AGEMA_signal_14423, new_AGEMA_signal_14422, MixColumnsIns_MixOneColumnInst_2_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U2 ( .a ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .b ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .c ({new_AGEMA_signal_13755, new_AGEMA_signal_13754, new_AGEMA_signal_13753, MixColumnsIns_MixOneColumnInst_2_n23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_U1 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .c ({new_AGEMA_signal_13758, new_AGEMA_signal_13757, new_AGEMA_signal_13756, MixColumnsIns_MixOneColumnInst_2_n59}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_13218, new_AGEMA_signal_13217, new_AGEMA_signal_13216, MixColumnsInput[59]}), .c ({new_AGEMA_signal_13761, new_AGEMA_signal_13760, new_AGEMA_signal_13759, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_13221, new_AGEMA_signal_13220, new_AGEMA_signal_13219, MixColumnsInput[58]}), .c ({new_AGEMA_signal_13764, new_AGEMA_signal_13763, new_AGEMA_signal_13762, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13206, new_AGEMA_signal_13205, new_AGEMA_signal_13204, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[24]}), .b ({new_AGEMA_signal_12696, new_AGEMA_signal_12695, new_AGEMA_signal_12694, MixColumnsInput[56]}), .c ({new_AGEMA_signal_13767, new_AGEMA_signal_13766, new_AGEMA_signal_13765, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_13113, new_AGEMA_signal_13112, new_AGEMA_signal_13111, MixColumnsInput[51]}), .c ({new_AGEMA_signal_13770, new_AGEMA_signal_13769, new_AGEMA_signal_13768, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_13116, new_AGEMA_signal_13115, new_AGEMA_signal_13114, MixColumnsInput[50]}), .c ({new_AGEMA_signal_13773, new_AGEMA_signal_13772, new_AGEMA_signal_13771, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13101, new_AGEMA_signal_13100, new_AGEMA_signal_13099, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[16]}), .b ({new_AGEMA_signal_12531, new_AGEMA_signal_12530, new_AGEMA_signal_12529, MixColumnsInput[48]}), .c ({new_AGEMA_signal_13776, new_AGEMA_signal_13775, new_AGEMA_signal_13774, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_13344, new_AGEMA_signal_13343, new_AGEMA_signal_13342, MixColumnsInput[43]}), .c ({new_AGEMA_signal_13779, new_AGEMA_signal_13778, new_AGEMA_signal_13777, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_13347, new_AGEMA_signal_13346, new_AGEMA_signal_13345, MixColumnsInput[42]}), .c ({new_AGEMA_signal_13782, new_AGEMA_signal_13781, new_AGEMA_signal_13780, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13332, new_AGEMA_signal_13331, new_AGEMA_signal_13330, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[8]}), .b ({new_AGEMA_signal_12894, new_AGEMA_signal_12893, new_AGEMA_signal_12892, MixColumnsInput[40]}), .c ({new_AGEMA_signal_13785, new_AGEMA_signal_13784, new_AGEMA_signal_13783, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13239, new_AGEMA_signal_13238, new_AGEMA_signal_13237, MixColumnsInput[35]}), .c ({new_AGEMA_signal_13788, new_AGEMA_signal_13787, new_AGEMA_signal_13786, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_13242, new_AGEMA_signal_13241, new_AGEMA_signal_13240, MixColumnsInput[34]}), .c ({new_AGEMA_signal_13791, new_AGEMA_signal_13790, new_AGEMA_signal_13789, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_2_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13227, new_AGEMA_signal_13226, new_AGEMA_signal_13225, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[0]}), .b ({new_AGEMA_signal_12729, new_AGEMA_signal_12728, new_AGEMA_signal_12727, MixColumnsInput[32]}), .c ({new_AGEMA_signal_13794, new_AGEMA_signal_13793, new_AGEMA_signal_13792, MixColumnsIns_MixOneColumnInst_2_DoubleBytes[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U96 ( .a ({new_AGEMA_signal_15099, new_AGEMA_signal_15098, new_AGEMA_signal_15097, MixColumnsIns_MixOneColumnInst_3_n64}), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_15822, new_AGEMA_signal_15821, new_AGEMA_signal_15820, MixColumnsOutput[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U95 ( .a ({new_AGEMA_signal_14490, new_AGEMA_signal_14489, new_AGEMA_signal_14488, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_14478, new_AGEMA_signal_14477, new_AGEMA_signal_14476, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_15099, new_AGEMA_signal_15098, new_AGEMA_signal_15097, MixColumnsIns_MixOneColumnInst_3_n64}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U94 ( .a ({new_AGEMA_signal_14427, new_AGEMA_signal_14426, new_AGEMA_signal_14425, MixColumnsIns_MixOneColumnInst_3_n61}), .b ({new_AGEMA_signal_13824, new_AGEMA_signal_13823, new_AGEMA_signal_13822, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_15102, new_AGEMA_signal_15101, new_AGEMA_signal_15100, MixColumnsOutput[8]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U93 ( .a ({new_AGEMA_signal_13854, new_AGEMA_signal_13853, new_AGEMA_signal_13852, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .c ({new_AGEMA_signal_14427, new_AGEMA_signal_14426, new_AGEMA_signal_14425, MixColumnsIns_MixOneColumnInst_3_n61}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U92 ( .a ({new_AGEMA_signal_14430, new_AGEMA_signal_14429, new_AGEMA_signal_14428, MixColumnsIns_MixOneColumnInst_3_n58}), .b ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, new_AGEMA_signal_13795, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_15105, new_AGEMA_signal_15104, new_AGEMA_signal_15103, MixColumnsOutput[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U91 ( .a ({new_AGEMA_signal_13830, new_AGEMA_signal_13829, new_AGEMA_signal_13828, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .c ({new_AGEMA_signal_14430, new_AGEMA_signal_14429, new_AGEMA_signal_14428, MixColumnsIns_MixOneColumnInst_3_n58}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U90 ( .a ({new_AGEMA_signal_14433, new_AGEMA_signal_14432, new_AGEMA_signal_14431, MixColumnsIns_MixOneColumnInst_3_n55}), .b ({new_AGEMA_signal_13800, new_AGEMA_signal_13799, new_AGEMA_signal_13798, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_15108, new_AGEMA_signal_15107, new_AGEMA_signal_15106, MixColumnsOutput[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U89 ( .a ({new_AGEMA_signal_13836, new_AGEMA_signal_13835, new_AGEMA_signal_13834, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_14433, new_AGEMA_signal_14432, new_AGEMA_signal_14431, MixColumnsIns_MixOneColumnInst_3_n55}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U88 ( .a ({new_AGEMA_signal_14436, new_AGEMA_signal_14435, new_AGEMA_signal_14434, MixColumnsIns_MixOneColumnInst_3_n52}), .b ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, new_AGEMA_signal_13801, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_15111, new_AGEMA_signal_15110, new_AGEMA_signal_15109, MixColumnsOutput[5]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U87 ( .a ({new_AGEMA_signal_13842, new_AGEMA_signal_13841, new_AGEMA_signal_13840, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_14436, new_AGEMA_signal_14435, new_AGEMA_signal_14434, MixColumnsIns_MixOneColumnInst_3_n52}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U86 ( .a ({new_AGEMA_signal_15114, new_AGEMA_signal_15113, new_AGEMA_signal_15112, MixColumnsIns_MixOneColumnInst_3_n49}), .b ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, new_AGEMA_signal_14449, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_15825, new_AGEMA_signal_15824, new_AGEMA_signal_15823, MixColumnsOutput[4]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U85 ( .a ({new_AGEMA_signal_14508, new_AGEMA_signal_14507, new_AGEMA_signal_14506, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_15114, new_AGEMA_signal_15113, new_AGEMA_signal_15112, MixColumnsIns_MixOneColumnInst_3_n49}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U84 ( .a ({new_AGEMA_signal_15117, new_AGEMA_signal_15116, new_AGEMA_signal_15115, MixColumnsIns_MixOneColumnInst_3_n46}), .b ({new_AGEMA_signal_14454, new_AGEMA_signal_14453, new_AGEMA_signal_14452, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_15828, new_AGEMA_signal_15827, new_AGEMA_signal_15826, MixColumnsOutput[3]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U83 ( .a ({new_AGEMA_signal_14514, new_AGEMA_signal_14513, new_AGEMA_signal_14512, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .c ({new_AGEMA_signal_15117, new_AGEMA_signal_15116, new_AGEMA_signal_15115, MixColumnsIns_MixOneColumnInst_3_n46}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U82 ( .a ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, new_AGEMA_signal_14437, MixColumnsIns_MixOneColumnInst_3_n43}), .b ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, new_AGEMA_signal_13795, MixColumnsIns_MixOneColumnInst_3_n57}), .c ({new_AGEMA_signal_15120, new_AGEMA_signal_15119, new_AGEMA_signal_15118, MixColumnsOutput[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U81 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_13797, new_AGEMA_signal_13796, new_AGEMA_signal_13795, MixColumnsIns_MixOneColumnInst_3_n57}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U80 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, new_AGEMA_signal_13807, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_14439, new_AGEMA_signal_14438, new_AGEMA_signal_14437, MixColumnsIns_MixOneColumnInst_3_n43}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U79 ( .a ({new_AGEMA_signal_14442, new_AGEMA_signal_14441, new_AGEMA_signal_14440, MixColumnsIns_MixOneColumnInst_3_n41}), .b ({new_AGEMA_signal_13800, new_AGEMA_signal_13799, new_AGEMA_signal_13798, MixColumnsIns_MixOneColumnInst_3_n54}), .c ({new_AGEMA_signal_15123, new_AGEMA_signal_15122, new_AGEMA_signal_15121, MixColumnsOutput[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U78 ( .a ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .b ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_13800, new_AGEMA_signal_13799, new_AGEMA_signal_13798, MixColumnsIns_MixOneColumnInst_3_n54}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U77 ( .a ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_13812, new_AGEMA_signal_13811, new_AGEMA_signal_13810, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_14442, new_AGEMA_signal_14441, new_AGEMA_signal_14440, MixColumnsIns_MixOneColumnInst_3_n41}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U76 ( .a ({new_AGEMA_signal_14445, new_AGEMA_signal_14444, new_AGEMA_signal_14443, MixColumnsIns_MixOneColumnInst_3_n39}), .b ({new_AGEMA_signal_13806, new_AGEMA_signal_13805, new_AGEMA_signal_13804, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_15126, new_AGEMA_signal_15125, new_AGEMA_signal_15124, MixColumnsOutput[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U75 ( .a ({new_AGEMA_signal_13848, new_AGEMA_signal_13847, new_AGEMA_signal_13846, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .c ({new_AGEMA_signal_14445, new_AGEMA_signal_14444, new_AGEMA_signal_14443, MixColumnsIns_MixOneColumnInst_3_n39}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U74 ( .a ({new_AGEMA_signal_14448, new_AGEMA_signal_14447, new_AGEMA_signal_14446, MixColumnsIns_MixOneColumnInst_3_n36}), .b ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, new_AGEMA_signal_13801, MixColumnsIns_MixOneColumnInst_3_n51}), .c ({new_AGEMA_signal_15129, new_AGEMA_signal_15128, new_AGEMA_signal_15127, MixColumnsOutput[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U73 ( .a ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_13803, new_AGEMA_signal_13802, new_AGEMA_signal_13801, MixColumnsIns_MixOneColumnInst_3_n51}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U72 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, new_AGEMA_signal_13813, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_14448, new_AGEMA_signal_14447, new_AGEMA_signal_14446, MixColumnsIns_MixOneColumnInst_3_n36}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U71 ( .a ({new_AGEMA_signal_15132, new_AGEMA_signal_15131, new_AGEMA_signal_15130, MixColumnsIns_MixOneColumnInst_3_n34}), .b ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, new_AGEMA_signal_14449, MixColumnsIns_MixOneColumnInst_3_n48}), .c ({new_AGEMA_signal_15831, new_AGEMA_signal_15830, new_AGEMA_signal_15829, MixColumnsOutput[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U70 ( .a ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .b ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, new_AGEMA_signal_13855, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}), .c ({new_AGEMA_signal_14451, new_AGEMA_signal_14450, new_AGEMA_signal_14449, MixColumnsIns_MixOneColumnInst_3_n48}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U69 ( .a ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_14472, new_AGEMA_signal_14471, new_AGEMA_signal_14470, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_15132, new_AGEMA_signal_15131, new_AGEMA_signal_15130, MixColumnsIns_MixOneColumnInst_3_n34}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U68 ( .a ({new_AGEMA_signal_15135, new_AGEMA_signal_15134, new_AGEMA_signal_15133, MixColumnsIns_MixOneColumnInst_3_n32}), .b ({new_AGEMA_signal_14454, new_AGEMA_signal_14453, new_AGEMA_signal_14452, MixColumnsIns_MixOneColumnInst_3_n45}), .c ({new_AGEMA_signal_15834, new_AGEMA_signal_15833, new_AGEMA_signal_15832, MixColumnsOutput[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U67 ( .a ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .b ({new_AGEMA_signal_13860, new_AGEMA_signal_13859, new_AGEMA_signal_13858, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}), .c ({new_AGEMA_signal_14454, new_AGEMA_signal_14453, new_AGEMA_signal_14452, MixColumnsIns_MixOneColumnInst_3_n45}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U66 ( .a ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .b ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, new_AGEMA_signal_14479, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_15135, new_AGEMA_signal_15134, new_AGEMA_signal_15133, MixColumnsIns_MixOneColumnInst_3_n32}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U65 ( .a ({new_AGEMA_signal_14457, new_AGEMA_signal_14456, new_AGEMA_signal_14455, MixColumnsIns_MixOneColumnInst_3_n30}), .b ({new_AGEMA_signal_13806, new_AGEMA_signal_13805, new_AGEMA_signal_13804, MixColumnsIns_MixOneColumnInst_3_n38}), .c ({new_AGEMA_signal_15138, new_AGEMA_signal_15137, new_AGEMA_signal_15136, MixColumnsOutput[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U64 ( .a ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .b ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_13806, new_AGEMA_signal_13805, new_AGEMA_signal_13804, MixColumnsIns_MixOneColumnInst_3_n38}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U63 ( .a ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .b ({new_AGEMA_signal_13818, new_AGEMA_signal_13817, new_AGEMA_signal_13816, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_14457, new_AGEMA_signal_14456, new_AGEMA_signal_14455, MixColumnsIns_MixOneColumnInst_3_n30}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U62 ( .a ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, new_AGEMA_signal_15139, MixColumnsIns_MixOneColumnInst_3_n28}), .b ({new_AGEMA_signal_14475, new_AGEMA_signal_14474, new_AGEMA_signal_14473, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_15837, new_AGEMA_signal_15836, new_AGEMA_signal_15835, MixColumnsOutput[25]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U61 ( .a ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, new_AGEMA_signal_14485, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_15141, new_AGEMA_signal_15140, new_AGEMA_signal_15139, MixColumnsIns_MixOneColumnInst_3_n28}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U60 ( .a ({new_AGEMA_signal_14460, new_AGEMA_signal_14459, new_AGEMA_signal_14458, MixColumnsIns_MixOneColumnInst_3_n25}), .b ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, new_AGEMA_signal_13819, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_15144, new_AGEMA_signal_15143, new_AGEMA_signal_15142, MixColumnsOutput[24]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U59 ( .a ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, new_AGEMA_signal_13849, MixColumnsIns_MixOneColumnInst_3_n23}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .c ({new_AGEMA_signal_14460, new_AGEMA_signal_14459, new_AGEMA_signal_14458, MixColumnsIns_MixOneColumnInst_3_n25}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U58 ( .a ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, new_AGEMA_signal_14461, MixColumnsIns_MixOneColumnInst_3_n22}), .b ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, new_AGEMA_signal_13807, MixColumnsIns_MixOneColumnInst_3_n42}), .c ({new_AGEMA_signal_15147, new_AGEMA_signal_15146, new_AGEMA_signal_15145, MixColumnsOutput[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U57 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_13809, new_AGEMA_signal_13808, new_AGEMA_signal_13807, MixColumnsIns_MixOneColumnInst_3_n42}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U56 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, new_AGEMA_signal_13825, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_14463, new_AGEMA_signal_14462, new_AGEMA_signal_14461, MixColumnsIns_MixOneColumnInst_3_n22}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U55 ( .a ({new_AGEMA_signal_14466, new_AGEMA_signal_14465, new_AGEMA_signal_14464, MixColumnsIns_MixOneColumnInst_3_n20}), .b ({new_AGEMA_signal_13812, new_AGEMA_signal_13811, new_AGEMA_signal_13810, MixColumnsIns_MixOneColumnInst_3_n40}), .c ({new_AGEMA_signal_15150, new_AGEMA_signal_15149, new_AGEMA_signal_15148, MixColumnsOutput[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U54 ( .a ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_13812, new_AGEMA_signal_13811, new_AGEMA_signal_13810, MixColumnsIns_MixOneColumnInst_3_n40}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U53 ( .a ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .b ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, new_AGEMA_signal_13831, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_14466, new_AGEMA_signal_14465, new_AGEMA_signal_14464, MixColumnsIns_MixOneColumnInst_3_n20}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U52 ( .a ({new_AGEMA_signal_14469, new_AGEMA_signal_14468, new_AGEMA_signal_14467, MixColumnsIns_MixOneColumnInst_3_n18}), .b ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, new_AGEMA_signal_13813, MixColumnsIns_MixOneColumnInst_3_n35}), .c ({new_AGEMA_signal_15153, new_AGEMA_signal_15152, new_AGEMA_signal_15151, MixColumnsOutput[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U51 ( .a ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .b ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_13815, new_AGEMA_signal_13814, new_AGEMA_signal_13813, MixColumnsIns_MixOneColumnInst_3_n35}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U50 ( .a ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .b ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, new_AGEMA_signal_13837, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_14469, new_AGEMA_signal_14468, new_AGEMA_signal_14467, MixColumnsIns_MixOneColumnInst_3_n18}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U49 ( .a ({new_AGEMA_signal_15156, new_AGEMA_signal_15155, new_AGEMA_signal_15154, MixColumnsIns_MixOneColumnInst_3_n16}), .b ({new_AGEMA_signal_14472, new_AGEMA_signal_14471, new_AGEMA_signal_14470, MixColumnsIns_MixOneColumnInst_3_n33}), .c ({new_AGEMA_signal_15840, new_AGEMA_signal_15839, new_AGEMA_signal_15838, MixColumnsOutput[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U48 ( .a ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .b ({new_AGEMA_signal_13866, new_AGEMA_signal_13865, new_AGEMA_signal_13864, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}), .c ({new_AGEMA_signal_14472, new_AGEMA_signal_14471, new_AGEMA_signal_14470, MixColumnsIns_MixOneColumnInst_3_n33}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U47 ( .a ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .b ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, new_AGEMA_signal_14503, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_15156, new_AGEMA_signal_15155, new_AGEMA_signal_15154, MixColumnsIns_MixOneColumnInst_3_n16}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U46 ( .a ({new_AGEMA_signal_15159, new_AGEMA_signal_15158, new_AGEMA_signal_15157, MixColumnsIns_MixOneColumnInst_3_n14}), .b ({new_AGEMA_signal_14475, new_AGEMA_signal_14474, new_AGEMA_signal_14473, MixColumnsIns_MixOneColumnInst_3_n27}), .c ({new_AGEMA_signal_15843, new_AGEMA_signal_15842, new_AGEMA_signal_15841, MixColumnsOutput[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U45 ( .a ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .b ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, new_AGEMA_signal_13861, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}), .c ({new_AGEMA_signal_14475, new_AGEMA_signal_14474, new_AGEMA_signal_14473, MixColumnsIns_MixOneColumnInst_3_n27}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U44 ( .a ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .b ({new_AGEMA_signal_14478, new_AGEMA_signal_14477, new_AGEMA_signal_14476, MixColumnsIns_MixOneColumnInst_3_n62}), .c ({new_AGEMA_signal_15159, new_AGEMA_signal_15158, new_AGEMA_signal_15157, MixColumnsIns_MixOneColumnInst_3_n14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U43 ( .a ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .b ({new_AGEMA_signal_13890, new_AGEMA_signal_13889, new_AGEMA_signal_13888, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}), .c ({new_AGEMA_signal_14478, new_AGEMA_signal_14477, new_AGEMA_signal_14476, MixColumnsIns_MixOneColumnInst_3_n62}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U42 ( .a ({new_AGEMA_signal_15162, new_AGEMA_signal_15161, new_AGEMA_signal_15160, MixColumnsIns_MixOneColumnInst_3_n13}), .b ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, new_AGEMA_signal_14479, MixColumnsIns_MixOneColumnInst_3_n31}), .c ({new_AGEMA_signal_15846, new_AGEMA_signal_15845, new_AGEMA_signal_15844, MixColumnsOutput[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U41 ( .a ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .b ({new_AGEMA_signal_13869, new_AGEMA_signal_13868, new_AGEMA_signal_13867, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}), .c ({new_AGEMA_signal_14481, new_AGEMA_signal_14480, new_AGEMA_signal_14479, MixColumnsIns_MixOneColumnInst_3_n31}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U40 ( .a ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .b ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, new_AGEMA_signal_14509, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_15162, new_AGEMA_signal_15161, new_AGEMA_signal_15160, MixColumnsIns_MixOneColumnInst_3_n13}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U39 ( .a ({new_AGEMA_signal_14484, new_AGEMA_signal_14483, new_AGEMA_signal_14482, MixColumnsIns_MixOneColumnInst_3_n11}), .b ({new_AGEMA_signal_13818, new_AGEMA_signal_13817, new_AGEMA_signal_13816, MixColumnsIns_MixOneColumnInst_3_n29}), .c ({new_AGEMA_signal_15165, new_AGEMA_signal_15164, new_AGEMA_signal_15163, MixColumnsOutput[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U38 ( .a ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .b ({new_AGEMA_signal_13371, new_AGEMA_signal_13370, new_AGEMA_signal_13369, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[18]}), .c ({new_AGEMA_signal_13818, new_AGEMA_signal_13817, new_AGEMA_signal_13816, MixColumnsIns_MixOneColumnInst_3_n29}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U37 ( .a ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .b ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, new_AGEMA_signal_13843, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_14484, new_AGEMA_signal_14483, new_AGEMA_signal_14482, MixColumnsIns_MixOneColumnInst_3_n11}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U36 ( .a ({new_AGEMA_signal_15168, new_AGEMA_signal_15167, new_AGEMA_signal_15166, MixColumnsIns_MixOneColumnInst_3_n9}), .b ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, new_AGEMA_signal_14485, MixColumnsIns_MixOneColumnInst_3_n26}), .c ({new_AGEMA_signal_15849, new_AGEMA_signal_15848, new_AGEMA_signal_15847, MixColumnsOutput[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U35 ( .a ({new_AGEMA_signal_13872, new_AGEMA_signal_13871, new_AGEMA_signal_13870, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}), .b ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_14487, new_AGEMA_signal_14486, new_AGEMA_signal_14485, MixColumnsIns_MixOneColumnInst_3_n26}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U34 ( .a ({new_AGEMA_signal_14490, new_AGEMA_signal_14489, new_AGEMA_signal_14488, MixColumnsIns_MixOneColumnInst_3_n63}), .b ({new_AGEMA_signal_13140, new_AGEMA_signal_13139, new_AGEMA_signal_13138, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[26]}), .c ({new_AGEMA_signal_15168, new_AGEMA_signal_15167, new_AGEMA_signal_15166, MixColumnsIns_MixOneColumnInst_3_n9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U33 ( .a ({new_AGEMA_signal_13881, new_AGEMA_signal_13880, new_AGEMA_signal_13879, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}), .b ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .c ({new_AGEMA_signal_14490, new_AGEMA_signal_14489, new_AGEMA_signal_14488, MixColumnsIns_MixOneColumnInst_3_n63}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U32 ( .a ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, new_AGEMA_signal_14491, MixColumnsIns_MixOneColumnInst_3_n8}), .b ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, new_AGEMA_signal_13819, MixColumnsIns_MixOneColumnInst_3_n24}), .c ({new_AGEMA_signal_15171, new_AGEMA_signal_15170, new_AGEMA_signal_15169, MixColumnsOutput[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U31 ( .a ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_13821, new_AGEMA_signal_13820, new_AGEMA_signal_13819, MixColumnsIns_MixOneColumnInst_3_n24}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U30 ( .a ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .b ({new_AGEMA_signal_13824, new_AGEMA_signal_13823, new_AGEMA_signal_13822, MixColumnsIns_MixOneColumnInst_3_n60}), .c ({new_AGEMA_signal_14493, new_AGEMA_signal_14492, new_AGEMA_signal_14491, MixColumnsIns_MixOneColumnInst_3_n8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U29 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .c ({new_AGEMA_signal_13824, new_AGEMA_signal_13823, new_AGEMA_signal_13822, MixColumnsIns_MixOneColumnInst_3_n60}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U28 ( .a ({new_AGEMA_signal_14496, new_AGEMA_signal_14495, new_AGEMA_signal_14494, MixColumnsIns_MixOneColumnInst_3_n7}), .b ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, new_AGEMA_signal_13825, MixColumnsIns_MixOneColumnInst_3_n21}), .c ({new_AGEMA_signal_15174, new_AGEMA_signal_15173, new_AGEMA_signal_15172, MixColumnsOutput[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U27 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13251, new_AGEMA_signal_13250, new_AGEMA_signal_13249, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[15]}), .c ({new_AGEMA_signal_13827, new_AGEMA_signal_13826, new_AGEMA_signal_13825, MixColumnsIns_MixOneColumnInst_3_n21}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U26 ( .a ({new_AGEMA_signal_13830, new_AGEMA_signal_13829, new_AGEMA_signal_13828, MixColumnsIns_MixOneColumnInst_3_n56}), .b ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .c ({new_AGEMA_signal_14496, new_AGEMA_signal_14495, new_AGEMA_signal_14494, MixColumnsIns_MixOneColumnInst_3_n7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U25 ( .a ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_13830, new_AGEMA_signal_13829, new_AGEMA_signal_13828, MixColumnsIns_MixOneColumnInst_3_n56}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U24 ( .a ({new_AGEMA_signal_14499, new_AGEMA_signal_14498, new_AGEMA_signal_14497, MixColumnsIns_MixOneColumnInst_3_n6}), .b ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, new_AGEMA_signal_13831, MixColumnsIns_MixOneColumnInst_3_n19}), .c ({new_AGEMA_signal_15177, new_AGEMA_signal_15176, new_AGEMA_signal_15175, MixColumnsOutput[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U23 ( .a ({new_AGEMA_signal_13146, new_AGEMA_signal_13145, new_AGEMA_signal_13144, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[7]}), .b ({new_AGEMA_signal_13254, new_AGEMA_signal_13253, new_AGEMA_signal_13252, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[14]}), .c ({new_AGEMA_signal_13833, new_AGEMA_signal_13832, new_AGEMA_signal_13831, MixColumnsIns_MixOneColumnInst_3_n19}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U22 ( .a ({new_AGEMA_signal_13836, new_AGEMA_signal_13835, new_AGEMA_signal_13834, MixColumnsIns_MixOneColumnInst_3_n53}), .b ({new_AGEMA_signal_13356, new_AGEMA_signal_13355, new_AGEMA_signal_13354, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[23]}), .c ({new_AGEMA_signal_14499, new_AGEMA_signal_14498, new_AGEMA_signal_14497, MixColumnsIns_MixOneColumnInst_3_n6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U21 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_13125, new_AGEMA_signal_13124, new_AGEMA_signal_13123, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[31]}), .c ({new_AGEMA_signal_13836, new_AGEMA_signal_13835, new_AGEMA_signal_13834, MixColumnsIns_MixOneColumnInst_3_n53}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U20 ( .a ({new_AGEMA_signal_14502, new_AGEMA_signal_14501, new_AGEMA_signal_14500, MixColumnsIns_MixOneColumnInst_3_n5}), .b ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, new_AGEMA_signal_13837, MixColumnsIns_MixOneColumnInst_3_n17}), .c ({new_AGEMA_signal_15180, new_AGEMA_signal_15179, new_AGEMA_signal_15178, MixColumnsOutput[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U19 ( .a ({new_AGEMA_signal_13149, new_AGEMA_signal_13148, new_AGEMA_signal_13147, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[6]}), .b ({new_AGEMA_signal_13257, new_AGEMA_signal_13256, new_AGEMA_signal_13255, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[13]}), .c ({new_AGEMA_signal_13839, new_AGEMA_signal_13838, new_AGEMA_signal_13837, MixColumnsIns_MixOneColumnInst_3_n17}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U18 ( .a ({new_AGEMA_signal_13842, new_AGEMA_signal_13841, new_AGEMA_signal_13840, MixColumnsIns_MixOneColumnInst_3_n50}), .b ({new_AGEMA_signal_13359, new_AGEMA_signal_13358, new_AGEMA_signal_13357, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[22]}), .c ({new_AGEMA_signal_14502, new_AGEMA_signal_14501, new_AGEMA_signal_14500, MixColumnsIns_MixOneColumnInst_3_n5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U17 ( .a ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_13128, new_AGEMA_signal_13127, new_AGEMA_signal_13126, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[30]}), .c ({new_AGEMA_signal_13842, new_AGEMA_signal_13841, new_AGEMA_signal_13840, MixColumnsIns_MixOneColumnInst_3_n50}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U16 ( .a ({new_AGEMA_signal_15183, new_AGEMA_signal_15182, new_AGEMA_signal_15181, MixColumnsIns_MixOneColumnInst_3_n4}), .b ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, new_AGEMA_signal_14503, MixColumnsIns_MixOneColumnInst_3_n15}), .c ({new_AGEMA_signal_15852, new_AGEMA_signal_15851, new_AGEMA_signal_15850, MixColumnsOutput[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U15 ( .a ({new_AGEMA_signal_13152, new_AGEMA_signal_13151, new_AGEMA_signal_13150, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[5]}), .b ({new_AGEMA_signal_13875, new_AGEMA_signal_13874, new_AGEMA_signal_13873, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}), .c ({new_AGEMA_signal_14505, new_AGEMA_signal_14504, new_AGEMA_signal_14503, MixColumnsIns_MixOneColumnInst_3_n15}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U14 ( .a ({new_AGEMA_signal_14508, new_AGEMA_signal_14507, new_AGEMA_signal_14506, MixColumnsIns_MixOneColumnInst_3_n47}), .b ({new_AGEMA_signal_13362, new_AGEMA_signal_13361, new_AGEMA_signal_13360, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[21]}), .c ({new_AGEMA_signal_15183, new_AGEMA_signal_15182, new_AGEMA_signal_15181, MixColumnsIns_MixOneColumnInst_3_n4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U13 ( .a ({new_AGEMA_signal_13884, new_AGEMA_signal_13883, new_AGEMA_signal_13882, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}), .b ({new_AGEMA_signal_13131, new_AGEMA_signal_13130, new_AGEMA_signal_13129, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[29]}), .c ({new_AGEMA_signal_14508, new_AGEMA_signal_14507, new_AGEMA_signal_14506, MixColumnsIns_MixOneColumnInst_3_n47}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U12 ( .a ({new_AGEMA_signal_15186, new_AGEMA_signal_15185, new_AGEMA_signal_15184, MixColumnsIns_MixOneColumnInst_3_n3}), .b ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, new_AGEMA_signal_14509, MixColumnsIns_MixOneColumnInst_3_n12}), .c ({new_AGEMA_signal_15855, new_AGEMA_signal_15854, new_AGEMA_signal_15853, MixColumnsOutput[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U11 ( .a ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .b ({new_AGEMA_signal_13878, new_AGEMA_signal_13877, new_AGEMA_signal_13876, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}), .c ({new_AGEMA_signal_14511, new_AGEMA_signal_14510, new_AGEMA_signal_14509, MixColumnsIns_MixOneColumnInst_3_n12}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U10 ( .a ({new_AGEMA_signal_14514, new_AGEMA_signal_14513, new_AGEMA_signal_14512, MixColumnsIns_MixOneColumnInst_3_n44}), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .c ({new_AGEMA_signal_15186, new_AGEMA_signal_15185, new_AGEMA_signal_15184, MixColumnsIns_MixOneColumnInst_3_n3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U9 ( .a ({new_AGEMA_signal_13887, new_AGEMA_signal_13886, new_AGEMA_signal_13885, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}), .b ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .c ({new_AGEMA_signal_14514, new_AGEMA_signal_14513, new_AGEMA_signal_14512, MixColumnsIns_MixOneColumnInst_3_n44}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U8 ( .a ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, new_AGEMA_signal_14515, MixColumnsIns_MixOneColumnInst_3_n2}), .b ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, new_AGEMA_signal_13843, MixColumnsIns_MixOneColumnInst_3_n10}), .c ({new_AGEMA_signal_15189, new_AGEMA_signal_15188, new_AGEMA_signal_15187, MixColumnsOutput[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U7 ( .a ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .b ({new_AGEMA_signal_13266, new_AGEMA_signal_13265, new_AGEMA_signal_13264, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[10]}), .c ({new_AGEMA_signal_13845, new_AGEMA_signal_13844, new_AGEMA_signal_13843, MixColumnsIns_MixOneColumnInst_3_n10}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U6 ( .a ({new_AGEMA_signal_13848, new_AGEMA_signal_13847, new_AGEMA_signal_13846, MixColumnsIns_MixOneColumnInst_3_n37}), .b ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .c ({new_AGEMA_signal_14517, new_AGEMA_signal_14516, new_AGEMA_signal_14515, MixColumnsIns_MixOneColumnInst_3_n2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U5 ( .a ({new_AGEMA_signal_13161, new_AGEMA_signal_13160, new_AGEMA_signal_13159, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[2]}), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .c ({new_AGEMA_signal_13848, new_AGEMA_signal_13847, new_AGEMA_signal_13846, MixColumnsIns_MixOneColumnInst_3_n37}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U4 ( .a ({new_AGEMA_signal_14520, new_AGEMA_signal_14519, new_AGEMA_signal_14518, MixColumnsIns_MixOneColumnInst_3_n1}), .b ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .c ({new_AGEMA_signal_15192, new_AGEMA_signal_15191, new_AGEMA_signal_15190, MixColumnsOutput[0]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U3 ( .a ({new_AGEMA_signal_13854, new_AGEMA_signal_13853, new_AGEMA_signal_13852, MixColumnsIns_MixOneColumnInst_3_n59}), .b ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, new_AGEMA_signal_13849, MixColumnsIns_MixOneColumnInst_3_n23}), .c ({new_AGEMA_signal_14520, new_AGEMA_signal_14519, new_AGEMA_signal_14518, MixColumnsIns_MixOneColumnInst_3_n1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U2 ( .a ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .b ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .c ({new_AGEMA_signal_13851, new_AGEMA_signal_13850, new_AGEMA_signal_13849, MixColumnsIns_MixOneColumnInst_3_n23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_U1 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .c ({new_AGEMA_signal_13854, new_AGEMA_signal_13853, new_AGEMA_signal_13852, MixColumnsIns_MixOneColumnInst_3_n59}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U3 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_13134, new_AGEMA_signal_13133, new_AGEMA_signal_13132, MixColumnsInput[27]}), .c ({new_AGEMA_signal_13857, new_AGEMA_signal_13856, new_AGEMA_signal_13855, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U2 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_13137, new_AGEMA_signal_13136, new_AGEMA_signal_13135, MixColumnsInput[26]}), .c ({new_AGEMA_signal_13860, new_AGEMA_signal_13859, new_AGEMA_signal_13858, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_0_U1 ( .a ({new_AGEMA_signal_13122, new_AGEMA_signal_13121, new_AGEMA_signal_13120, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[24]}), .b ({new_AGEMA_signal_12564, new_AGEMA_signal_12563, new_AGEMA_signal_12562, MixColumnsInput[24]}), .c ({new_AGEMA_signal_13863, new_AGEMA_signal_13862, new_AGEMA_signal_13861, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U3 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_13365, new_AGEMA_signal_13364, new_AGEMA_signal_13363, MixColumnsInput[19]}), .c ({new_AGEMA_signal_13866, new_AGEMA_signal_13865, new_AGEMA_signal_13864, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U2 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_13368, new_AGEMA_signal_13367, new_AGEMA_signal_13366, MixColumnsInput[18]}), .c ({new_AGEMA_signal_13869, new_AGEMA_signal_13868, new_AGEMA_signal_13867, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_1_U1 ( .a ({new_AGEMA_signal_13353, new_AGEMA_signal_13352, new_AGEMA_signal_13351, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[16]}), .b ({new_AGEMA_signal_12927, new_AGEMA_signal_12926, new_AGEMA_signal_12925, MixColumnsInput[16]}), .c ({new_AGEMA_signal_13872, new_AGEMA_signal_13871, new_AGEMA_signal_13870, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U3 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_13260, new_AGEMA_signal_13259, new_AGEMA_signal_13258, MixColumnsInput[11]}), .c ({new_AGEMA_signal_13875, new_AGEMA_signal_13874, new_AGEMA_signal_13873, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U2 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_13263, new_AGEMA_signal_13262, new_AGEMA_signal_13261, MixColumnsInput[10]}), .c ({new_AGEMA_signal_13878, new_AGEMA_signal_13877, new_AGEMA_signal_13876, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_2_U1 ( .a ({new_AGEMA_signal_13248, new_AGEMA_signal_13247, new_AGEMA_signal_13246, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[8]}), .b ({new_AGEMA_signal_12762, new_AGEMA_signal_12761, new_AGEMA_signal_12760, MixColumnsInput[8]}), .c ({new_AGEMA_signal_13881, new_AGEMA_signal_13880, new_AGEMA_signal_13879, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U3 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13155, new_AGEMA_signal_13154, new_AGEMA_signal_13153, MixColumnsInput[3]}), .c ({new_AGEMA_signal_13884, new_AGEMA_signal_13883, new_AGEMA_signal_13882, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U2 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_13158, new_AGEMA_signal_13157, new_AGEMA_signal_13156, MixColumnsInput[2]}), .c ({new_AGEMA_signal_13887, new_AGEMA_signal_13886, new_AGEMA_signal_13885, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) MixColumnsIns_MixOneColumnInst_3_Mul2Inst_3_U1 ( .a ({new_AGEMA_signal_13143, new_AGEMA_signal_13142, new_AGEMA_signal_13141, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[0]}), .b ({new_AGEMA_signal_12597, new_AGEMA_signal_12596, new_AGEMA_signal_12595, MixColumnsInput[0]}), .c ({new_AGEMA_signal_13890, new_AGEMA_signal_13889, new_AGEMA_signal_13888, MixColumnsIns_MixOneColumnInst_3_DoubleBytes[1]}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_0_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14808, new_AGEMA_signal_14807, new_AGEMA_signal_14806, KeyExpansionOutput[0]}), .a ({key_s3[0], key_s2[0], key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_15198, new_AGEMA_signal_15197, new_AGEMA_signal_15196, KeyReg_Inst_ff_SDE_0_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_1_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15444, new_AGEMA_signal_15443, new_AGEMA_signal_15442, KeyExpansionOutput[1]}), .a ({key_s3[1], key_s2[1], key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_15861, new_AGEMA_signal_15860, new_AGEMA_signal_15859, KeyReg_Inst_ff_SDE_1_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_2_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15411, new_AGEMA_signal_15410, new_AGEMA_signal_15409, KeyExpansionOutput[2]}), .a ({key_s3[2], key_s2[2], key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_15867, new_AGEMA_signal_15866, new_AGEMA_signal_15865, KeyReg_Inst_ff_SDE_2_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_3_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15402, new_AGEMA_signal_15401, new_AGEMA_signal_15400, KeyExpansionOutput[3]}), .a ({key_s3[3], key_s2[3], key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_15873, new_AGEMA_signal_15872, new_AGEMA_signal_15871, KeyReg_Inst_ff_SDE_3_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_4_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15399, new_AGEMA_signal_15398, new_AGEMA_signal_15397, KeyExpansionOutput[4]}), .a ({key_s3[4], key_s2[4], key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_15879, new_AGEMA_signal_15878, new_AGEMA_signal_15877, KeyReg_Inst_ff_SDE_4_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_5_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15396, new_AGEMA_signal_15395, new_AGEMA_signal_15394, KeyExpansionOutput[5]}), .a ({key_s3[5], key_s2[5], key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_15885, new_AGEMA_signal_15884, new_AGEMA_signal_15883, KeyReg_Inst_ff_SDE_5_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_6_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15393, new_AGEMA_signal_15392, new_AGEMA_signal_15391, KeyExpansionOutput[6]}), .a ({key_s3[6], key_s2[6], key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_15891, new_AGEMA_signal_15890, new_AGEMA_signal_15889, KeyReg_Inst_ff_SDE_6_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_7_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15390, new_AGEMA_signal_15389, new_AGEMA_signal_15388, KeyExpansionOutput[7]}), .a ({key_s3[7], key_s2[7], key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_15897, new_AGEMA_signal_15896, new_AGEMA_signal_15895, KeyReg_Inst_ff_SDE_7_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_8_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, new_AGEMA_signal_14713, KeyExpansionOutput[8]}), .a ({key_s3[8], key_s2[8], key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_15204, new_AGEMA_signal_15203, new_AGEMA_signal_15202, KeyReg_Inst_ff_SDE_8_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_9_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15387, new_AGEMA_signal_15386, new_AGEMA_signal_15385, KeyExpansionOutput[9]}), .a ({key_s3[9], key_s2[9], key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_15903, new_AGEMA_signal_15902, new_AGEMA_signal_15901, KeyReg_Inst_ff_SDE_9_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_10_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15471, new_AGEMA_signal_15470, new_AGEMA_signal_15469, KeyExpansionOutput[10]}), .a ({key_s3[10], key_s2[10], key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_15909, new_AGEMA_signal_15908, new_AGEMA_signal_15907, KeyReg_Inst_ff_SDE_10_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_11_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15468, new_AGEMA_signal_15467, new_AGEMA_signal_15466, KeyExpansionOutput[11]}), .a ({key_s3[11], key_s2[11], key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_15915, new_AGEMA_signal_15914, new_AGEMA_signal_15913, KeyReg_Inst_ff_SDE_11_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_12_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15465, new_AGEMA_signal_15464, new_AGEMA_signal_15463, KeyExpansionOutput[12]}), .a ({key_s3[12], key_s2[12], key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_15921, new_AGEMA_signal_15920, new_AGEMA_signal_15919, KeyReg_Inst_ff_SDE_12_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_13_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15462, new_AGEMA_signal_15461, new_AGEMA_signal_15460, KeyExpansionOutput[13]}), .a ({key_s3[13], key_s2[13], key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_15927, new_AGEMA_signal_15926, new_AGEMA_signal_15925, KeyReg_Inst_ff_SDE_13_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_14_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15459, new_AGEMA_signal_15458, new_AGEMA_signal_15457, KeyExpansionOutput[14]}), .a ({key_s3[14], key_s2[14], key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_15933, new_AGEMA_signal_15932, new_AGEMA_signal_15931, KeyReg_Inst_ff_SDE_14_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_15_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15456, new_AGEMA_signal_15455, new_AGEMA_signal_15454, KeyExpansionOutput[15]}), .a ({key_s3[15], key_s2[15], key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_15939, new_AGEMA_signal_15938, new_AGEMA_signal_15937, KeyReg_Inst_ff_SDE_15_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_16_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14787, new_AGEMA_signal_14786, new_AGEMA_signal_14785, KeyExpansionOutput[16]}), .a ({key_s3[16], key_s2[16], key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_15210, new_AGEMA_signal_15209, new_AGEMA_signal_15208, KeyReg_Inst_ff_SDE_16_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_17_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15453, new_AGEMA_signal_15452, new_AGEMA_signal_15451, KeyExpansionOutput[17]}), .a ({key_s3[17], key_s2[17], key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_15945, new_AGEMA_signal_15944, new_AGEMA_signal_15943, KeyReg_Inst_ff_SDE_17_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_18_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15450, new_AGEMA_signal_15449, new_AGEMA_signal_15448, KeyExpansionOutput[18]}), .a ({key_s3[18], key_s2[18], key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_15951, new_AGEMA_signal_15950, new_AGEMA_signal_15949, KeyReg_Inst_ff_SDE_18_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_19_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15447, new_AGEMA_signal_15446, new_AGEMA_signal_15445, KeyExpansionOutput[19]}), .a ({key_s3[19], key_s2[19], key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_15957, new_AGEMA_signal_15956, new_AGEMA_signal_15955, KeyReg_Inst_ff_SDE_19_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_20_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15441, new_AGEMA_signal_15440, new_AGEMA_signal_15439, KeyExpansionOutput[20]}), .a ({key_s3[20], key_s2[20], key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_15963, new_AGEMA_signal_15962, new_AGEMA_signal_15961, KeyReg_Inst_ff_SDE_20_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_21_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15438, new_AGEMA_signal_15437, new_AGEMA_signal_15436, KeyExpansionOutput[21]}), .a ({key_s3[21], key_s2[21], key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_15969, new_AGEMA_signal_15968, new_AGEMA_signal_15967, KeyReg_Inst_ff_SDE_21_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_22_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15435, new_AGEMA_signal_15434, new_AGEMA_signal_15433, KeyExpansionOutput[22]}), .a ({key_s3[22], key_s2[22], key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_15975, new_AGEMA_signal_15974, new_AGEMA_signal_15973, KeyReg_Inst_ff_SDE_22_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_23_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15432, new_AGEMA_signal_15431, new_AGEMA_signal_15430, KeyExpansionOutput[23]}), .a ({key_s3[23], key_s2[23], key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_15981, new_AGEMA_signal_15980, new_AGEMA_signal_15979, KeyReg_Inst_ff_SDE_23_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_24_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15429, new_AGEMA_signal_15428, new_AGEMA_signal_15427, KeyExpansionOutput[24]}), .a ({key_s3[24], key_s2[24], key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_15987, new_AGEMA_signal_15986, new_AGEMA_signal_15985, KeyReg_Inst_ff_SDE_24_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_25_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16050, new_AGEMA_signal_16049, new_AGEMA_signal_16048, KeyExpansionOutput[25]}), .a ({key_s3[25], key_s2[25], key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_16680, new_AGEMA_signal_16679, new_AGEMA_signal_16678, KeyReg_Inst_ff_SDE_25_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_26_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, new_AGEMA_signal_16045, KeyExpansionOutput[26]}), .a ({key_s3[26], key_s2[26], key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_16686, new_AGEMA_signal_16685, new_AGEMA_signal_16684, KeyReg_Inst_ff_SDE_26_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_27_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16044, new_AGEMA_signal_16043, new_AGEMA_signal_16042, KeyExpansionOutput[27]}), .a ({key_s3[27], key_s2[27], key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_16692, new_AGEMA_signal_16691, new_AGEMA_signal_16690, KeyReg_Inst_ff_SDE_27_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_28_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, new_AGEMA_signal_16039, KeyExpansionOutput[28]}), .a ({key_s3[28], key_s2[28], key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_16698, new_AGEMA_signal_16697, new_AGEMA_signal_16696, KeyReg_Inst_ff_SDE_28_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_29_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16038, new_AGEMA_signal_16037, new_AGEMA_signal_16036, KeyExpansionOutput[29]}), .a ({key_s3[29], key_s2[29], key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_16704, new_AGEMA_signal_16703, new_AGEMA_signal_16702, KeyReg_Inst_ff_SDE_29_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_30_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16035, new_AGEMA_signal_16034, new_AGEMA_signal_16033, KeyExpansionOutput[30]}), .a ({key_s3[30], key_s2[30], key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_16710, new_AGEMA_signal_16709, new_AGEMA_signal_16708, KeyReg_Inst_ff_SDE_30_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_31_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_16032, new_AGEMA_signal_16031, new_AGEMA_signal_16030, KeyExpansionOutput[31]}), .a ({key_s3[31], key_s2[31], key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_16716, new_AGEMA_signal_16715, new_AGEMA_signal_16714, KeyReg_Inst_ff_SDE_31_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_32_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14136, new_AGEMA_signal_14135, new_AGEMA_signal_14134, KeyExpansionOutput[32]}), .a ({key_s3[32], key_s2[32], key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_14526, new_AGEMA_signal_14525, new_AGEMA_signal_14524, KeyReg_Inst_ff_SDE_32_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_33_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, new_AGEMA_signal_14773, KeyExpansionOutput[33]}), .a ({key_s3[33], key_s2[33], key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_15216, new_AGEMA_signal_15215, new_AGEMA_signal_15214, KeyReg_Inst_ff_SDE_33_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_34_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14742, new_AGEMA_signal_14741, new_AGEMA_signal_14740, KeyExpansionOutput[34]}), .a ({key_s3[34], key_s2[34], key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_15222, new_AGEMA_signal_15221, new_AGEMA_signal_15220, KeyReg_Inst_ff_SDE_34_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_35_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, new_AGEMA_signal_14731, KeyExpansionOutput[35]}), .a ({key_s3[35], key_s2[35], key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_15228, new_AGEMA_signal_15227, new_AGEMA_signal_15226, KeyReg_Inst_ff_SDE_35_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_36_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14730, new_AGEMA_signal_14729, new_AGEMA_signal_14728, KeyExpansionOutput[36]}), .a ({key_s3[36], key_s2[36], key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_15234, new_AGEMA_signal_15233, new_AGEMA_signal_15232, KeyReg_Inst_ff_SDE_36_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_37_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, new_AGEMA_signal_14725, KeyExpansionOutput[37]}), .a ({key_s3[37], key_s2[37], key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_15240, new_AGEMA_signal_15239, new_AGEMA_signal_15238, KeyReg_Inst_ff_SDE_37_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_38_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14724, new_AGEMA_signal_14723, new_AGEMA_signal_14722, KeyExpansionOutput[38]}), .a ({key_s3[38], key_s2[38], key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_15246, new_AGEMA_signal_15245, new_AGEMA_signal_15244, KeyReg_Inst_ff_SDE_38_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_39_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, new_AGEMA_signal_14719, KeyExpansionOutput[39]}), .a ({key_s3[39], key_s2[39], key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_15252, new_AGEMA_signal_15251, new_AGEMA_signal_15250, KeyReg_Inst_ff_SDE_39_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_40_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14046, new_AGEMA_signal_14045, new_AGEMA_signal_14044, KeyExpansionOutput[40]}), .a ({key_s3[40], key_s2[40], key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_14532, new_AGEMA_signal_14531, new_AGEMA_signal_14530, KeyReg_Inst_ff_SDE_40_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_41_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14718, new_AGEMA_signal_14717, new_AGEMA_signal_14716, KeyExpansionOutput[41]}), .a ({key_s3[41], key_s2[41], key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_15258, new_AGEMA_signal_15257, new_AGEMA_signal_15256, KeyReg_Inst_ff_SDE_41_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_42_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14805, new_AGEMA_signal_14804, new_AGEMA_signal_14803, KeyExpansionOutput[42]}), .a ({key_s3[42], key_s2[42], key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_15264, new_AGEMA_signal_15263, new_AGEMA_signal_15262, KeyReg_Inst_ff_SDE_42_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_43_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14802, new_AGEMA_signal_14801, new_AGEMA_signal_14800, KeyExpansionOutput[43]}), .a ({key_s3[43], key_s2[43], key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_15270, new_AGEMA_signal_15269, new_AGEMA_signal_15268, KeyReg_Inst_ff_SDE_43_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_44_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, new_AGEMA_signal_14797, KeyExpansionOutput[44]}), .a ({key_s3[44], key_s2[44], key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_15276, new_AGEMA_signal_15275, new_AGEMA_signal_15274, KeyReg_Inst_ff_SDE_44_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_45_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14796, new_AGEMA_signal_14795, new_AGEMA_signal_14794, KeyExpansionOutput[45]}), .a ({key_s3[45], key_s2[45], key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_15282, new_AGEMA_signal_15281, new_AGEMA_signal_15280, KeyReg_Inst_ff_SDE_45_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_46_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, new_AGEMA_signal_14791, KeyExpansionOutput[46]}), .a ({key_s3[46], key_s2[46], key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_15288, new_AGEMA_signal_15287, new_AGEMA_signal_15286, KeyReg_Inst_ff_SDE_46_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_47_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14790, new_AGEMA_signal_14789, new_AGEMA_signal_14788, KeyExpansionOutput[47]}), .a ({key_s3[47], key_s2[47], key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_15294, new_AGEMA_signal_15293, new_AGEMA_signal_15292, KeyReg_Inst_ff_SDE_47_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_48_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14094, new_AGEMA_signal_14093, new_AGEMA_signal_14092, KeyExpansionOutput[48]}), .a ({key_s3[48], key_s2[48], key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_14538, new_AGEMA_signal_14537, new_AGEMA_signal_14536, KeyReg_Inst_ff_SDE_48_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_49_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14784, new_AGEMA_signal_14783, new_AGEMA_signal_14782, KeyExpansionOutput[49]}), .a ({key_s3[49], key_s2[49], key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_15300, new_AGEMA_signal_15299, new_AGEMA_signal_15298, KeyReg_Inst_ff_SDE_49_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_50_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, new_AGEMA_signal_14779, KeyExpansionOutput[50]}), .a ({key_s3[50], key_s2[50], key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_15306, new_AGEMA_signal_15305, new_AGEMA_signal_15304, KeyReg_Inst_ff_SDE_50_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_51_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14778, new_AGEMA_signal_14777, new_AGEMA_signal_14776, KeyExpansionOutput[51]}), .a ({key_s3[51], key_s2[51], key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_15312, new_AGEMA_signal_15311, new_AGEMA_signal_15310, KeyReg_Inst_ff_SDE_51_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_52_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14772, new_AGEMA_signal_14771, new_AGEMA_signal_14770, KeyExpansionOutput[52]}), .a ({key_s3[52], key_s2[52], key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_15318, new_AGEMA_signal_15317, new_AGEMA_signal_15316, KeyReg_Inst_ff_SDE_52_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_53_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, new_AGEMA_signal_14767, KeyExpansionOutput[53]}), .a ({key_s3[53], key_s2[53], key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_15324, new_AGEMA_signal_15323, new_AGEMA_signal_15322, KeyReg_Inst_ff_SDE_53_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_54_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14766, new_AGEMA_signal_14765, new_AGEMA_signal_14764, KeyExpansionOutput[54]}), .a ({key_s3[54], key_s2[54], key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_15330, new_AGEMA_signal_15329, new_AGEMA_signal_15328, KeyReg_Inst_ff_SDE_54_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_55_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, new_AGEMA_signal_14761, KeyExpansionOutput[55]}), .a ({key_s3[55], key_s2[55], key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_15336, new_AGEMA_signal_15335, new_AGEMA_signal_15334, KeyReg_Inst_ff_SDE_55_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_56_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14760, new_AGEMA_signal_14759, new_AGEMA_signal_14758, KeyExpansionOutput[56]}), .a ({key_s3[56], key_s2[56], key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_15342, new_AGEMA_signal_15341, new_AGEMA_signal_15340, KeyReg_Inst_ff_SDE_56_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_57_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15426, new_AGEMA_signal_15425, new_AGEMA_signal_15424, KeyExpansionOutput[57]}), .a ({key_s3[57], key_s2[57], key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_15993, new_AGEMA_signal_15992, new_AGEMA_signal_15991, KeyReg_Inst_ff_SDE_57_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_58_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15423, new_AGEMA_signal_15422, new_AGEMA_signal_15421, KeyExpansionOutput[58]}), .a ({key_s3[58], key_s2[58], key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_15999, new_AGEMA_signal_15998, new_AGEMA_signal_15997, KeyReg_Inst_ff_SDE_58_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_59_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15420, new_AGEMA_signal_15419, new_AGEMA_signal_15418, KeyExpansionOutput[59]}), .a ({key_s3[59], key_s2[59], key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, new_AGEMA_signal_16003, KeyReg_Inst_ff_SDE_59_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_60_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15417, new_AGEMA_signal_15416, new_AGEMA_signal_15415, KeyExpansionOutput[60]}), .a ({key_s3[60], key_s2[60], key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, new_AGEMA_signal_16009, KeyReg_Inst_ff_SDE_60_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_61_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15414, new_AGEMA_signal_15413, new_AGEMA_signal_15412, KeyExpansionOutput[61]}), .a ({key_s3[61], key_s2[61], key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_16017, new_AGEMA_signal_16016, new_AGEMA_signal_16015, KeyReg_Inst_ff_SDE_61_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_62_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15408, new_AGEMA_signal_15407, new_AGEMA_signal_15406, KeyExpansionOutput[62]}), .a ({key_s3[62], key_s2[62], key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_16023, new_AGEMA_signal_16022, new_AGEMA_signal_16021, KeyReg_Inst_ff_SDE_62_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_63_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_15405, new_AGEMA_signal_15404, new_AGEMA_signal_15403, KeyExpansionOutput[63]}), .a ({key_s3[63], key_s2[63], key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, new_AGEMA_signal_16027, KeyReg_Inst_ff_SDE_63_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_64_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, new_AGEMA_signal_13483, KeyExpansionOutput[64]}), .a ({key_s3[64], key_s2[64], key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_13896, new_AGEMA_signal_13895, new_AGEMA_signal_13894, KeyReg_Inst_ff_SDE_64_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_65_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14082, new_AGEMA_signal_14081, new_AGEMA_signal_14080, KeyExpansionOutput[65]}), .a ({key_s3[65], key_s2[65], key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_14544, new_AGEMA_signal_14543, new_AGEMA_signal_14542, KeyReg_Inst_ff_SDE_65_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_66_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14064, new_AGEMA_signal_14063, new_AGEMA_signal_14062, KeyExpansionOutput[66]}), .a ({key_s3[66], key_s2[66], key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_14550, new_AGEMA_signal_14549, new_AGEMA_signal_14548, KeyReg_Inst_ff_SDE_66_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_67_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, new_AGEMA_signal_14059, KeyExpansionOutput[67]}), .a ({key_s3[67], key_s2[67], key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_14556, new_AGEMA_signal_14555, new_AGEMA_signal_14554, KeyReg_Inst_ff_SDE_67_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_68_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14058, new_AGEMA_signal_14057, new_AGEMA_signal_14056, KeyExpansionOutput[68]}), .a ({key_s3[68], key_s2[68], key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_14562, new_AGEMA_signal_14561, new_AGEMA_signal_14560, KeyReg_Inst_ff_SDE_68_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_69_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, new_AGEMA_signal_14053, KeyExpansionOutput[69]}), .a ({key_s3[69], key_s2[69], key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_14568, new_AGEMA_signal_14567, new_AGEMA_signal_14566, KeyReg_Inst_ff_SDE_69_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_70_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14052, new_AGEMA_signal_14051, new_AGEMA_signal_14050, KeyExpansionOutput[70]}), .a ({key_s3[70], key_s2[70], key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_14574, new_AGEMA_signal_14573, new_AGEMA_signal_14572, KeyReg_Inst_ff_SDE_70_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_71_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, new_AGEMA_signal_14047, KeyExpansionOutput[71]}), .a ({key_s3[71], key_s2[71], key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_14580, new_AGEMA_signal_14579, new_AGEMA_signal_14578, KeyReg_Inst_ff_SDE_71_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_72_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, new_AGEMA_signal_13411, KeyExpansionOutput[72]}), .a ({key_s3[72], key_s2[72], key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_13902, new_AGEMA_signal_13901, new_AGEMA_signal_13900, KeyReg_Inst_ff_SDE_72_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_73_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, new_AGEMA_signal_14041, KeyExpansionOutput[73]}), .a ({key_s3[73], key_s2[73], key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_14586, new_AGEMA_signal_14585, new_AGEMA_signal_14584, KeyReg_Inst_ff_SDE_73_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_74_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, new_AGEMA_signal_14131, KeyExpansionOutput[74]}), .a ({key_s3[74], key_s2[74], key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_14592, new_AGEMA_signal_14591, new_AGEMA_signal_14590, KeyReg_Inst_ff_SDE_74_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_75_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14130, new_AGEMA_signal_14129, new_AGEMA_signal_14128, KeyExpansionOutput[75]}), .a ({key_s3[75], key_s2[75], key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_14598, new_AGEMA_signal_14597, new_AGEMA_signal_14596, KeyReg_Inst_ff_SDE_75_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_76_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14106, new_AGEMA_signal_14105, new_AGEMA_signal_14104, KeyExpansionOutput[76]}), .a ({key_s3[76], key_s2[76], key_s1[76], key_s0[76]}), .c ({new_AGEMA_signal_14604, new_AGEMA_signal_14603, new_AGEMA_signal_14602, KeyReg_Inst_ff_SDE_76_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_77_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, new_AGEMA_signal_14101, KeyExpansionOutput[77]}), .a ({key_s3[77], key_s2[77], key_s1[77], key_s0[77]}), .c ({new_AGEMA_signal_14610, new_AGEMA_signal_14609, new_AGEMA_signal_14608, KeyReg_Inst_ff_SDE_77_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_78_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14100, new_AGEMA_signal_14099, new_AGEMA_signal_14098, KeyExpansionOutput[78]}), .a ({key_s3[78], key_s2[78], key_s1[78], key_s0[78]}), .c ({new_AGEMA_signal_14616, new_AGEMA_signal_14615, new_AGEMA_signal_14614, KeyReg_Inst_ff_SDE_78_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_79_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, new_AGEMA_signal_14095, KeyExpansionOutput[79]}), .a ({key_s3[79], key_s2[79], key_s1[79], key_s0[79]}), .c ({new_AGEMA_signal_14622, new_AGEMA_signal_14621, new_AGEMA_signal_14620, KeyReg_Inst_ff_SDE_79_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_80_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, new_AGEMA_signal_13423, KeyExpansionOutput[80]}), .a ({key_s3[80], key_s2[80], key_s1[80], key_s0[80]}), .c ({new_AGEMA_signal_13908, new_AGEMA_signal_13907, new_AGEMA_signal_13906, KeyReg_Inst_ff_SDE_80_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_81_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, new_AGEMA_signal_14089, KeyExpansionOutput[81]}), .a ({key_s3[81], key_s2[81], key_s1[81], key_s0[81]}), .c ({new_AGEMA_signal_14628, new_AGEMA_signal_14627, new_AGEMA_signal_14626, KeyReg_Inst_ff_SDE_81_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_82_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14088, new_AGEMA_signal_14087, new_AGEMA_signal_14086, KeyExpansionOutput[82]}), .a ({key_s3[82], key_s2[82], key_s1[82], key_s0[82]}), .c ({new_AGEMA_signal_14634, new_AGEMA_signal_14633, new_AGEMA_signal_14632, KeyReg_Inst_ff_SDE_82_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_83_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, new_AGEMA_signal_14083, KeyExpansionOutput[83]}), .a ({key_s3[83], key_s2[83], key_s1[83], key_s0[83]}), .c ({new_AGEMA_signal_14640, new_AGEMA_signal_14639, new_AGEMA_signal_14638, KeyReg_Inst_ff_SDE_83_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_84_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, new_AGEMA_signal_14077, KeyExpansionOutput[84]}), .a ({key_s3[84], key_s2[84], key_s1[84], key_s0[84]}), .c ({new_AGEMA_signal_14646, new_AGEMA_signal_14645, new_AGEMA_signal_14644, KeyReg_Inst_ff_SDE_84_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_85_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14076, new_AGEMA_signal_14075, new_AGEMA_signal_14074, KeyExpansionOutput[85]}), .a ({key_s3[85], key_s2[85], key_s1[85], key_s0[85]}), .c ({new_AGEMA_signal_14652, new_AGEMA_signal_14651, new_AGEMA_signal_14650, KeyReg_Inst_ff_SDE_85_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_86_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, new_AGEMA_signal_14071, KeyExpansionOutput[86]}), .a ({key_s3[86], key_s2[86], key_s1[86], key_s0[86]}), .c ({new_AGEMA_signal_14658, new_AGEMA_signal_14657, new_AGEMA_signal_14656, KeyReg_Inst_ff_SDE_86_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_87_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14070, new_AGEMA_signal_14069, new_AGEMA_signal_14068, KeyExpansionOutput[87]}), .a ({key_s3[87], key_s2[87], key_s1[87], key_s0[87]}), .c ({new_AGEMA_signal_14664, new_AGEMA_signal_14663, new_AGEMA_signal_14662, KeyReg_Inst_ff_SDE_87_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_88_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, new_AGEMA_signal_14065, KeyExpansionOutput[88]}), .a ({key_s3[88], key_s2[88], key_s1[88], key_s0[88]}), .c ({new_AGEMA_signal_14670, new_AGEMA_signal_14669, new_AGEMA_signal_14668, KeyReg_Inst_ff_SDE_88_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_89_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, new_AGEMA_signal_14755, KeyExpansionOutput[89]}), .a ({key_s3[89], key_s2[89], key_s1[89], key_s0[89]}), .c ({new_AGEMA_signal_15348, new_AGEMA_signal_15347, new_AGEMA_signal_15346, KeyReg_Inst_ff_SDE_89_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_90_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14754, new_AGEMA_signal_14753, new_AGEMA_signal_14752, KeyExpansionOutput[90]}), .a ({key_s3[90], key_s2[90], key_s1[90], key_s0[90]}), .c ({new_AGEMA_signal_15354, new_AGEMA_signal_15353, new_AGEMA_signal_15352, KeyReg_Inst_ff_SDE_90_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_91_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, new_AGEMA_signal_14749, KeyExpansionOutput[91]}), .a ({key_s3[91], key_s2[91], key_s1[91], key_s0[91]}), .c ({new_AGEMA_signal_15360, new_AGEMA_signal_15359, new_AGEMA_signal_15358, KeyReg_Inst_ff_SDE_91_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_92_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14748, new_AGEMA_signal_14747, new_AGEMA_signal_14746, KeyExpansionOutput[92]}), .a ({key_s3[92], key_s2[92], key_s1[92], key_s0[92]}), .c ({new_AGEMA_signal_15366, new_AGEMA_signal_15365, new_AGEMA_signal_15364, KeyReg_Inst_ff_SDE_92_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_93_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, new_AGEMA_signal_14743, KeyExpansionOutput[93]}), .a ({key_s3[93], key_s2[93], key_s1[93], key_s0[93]}), .c ({new_AGEMA_signal_15372, new_AGEMA_signal_15371, new_AGEMA_signal_15370, KeyReg_Inst_ff_SDE_93_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_94_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, new_AGEMA_signal_14737, KeyExpansionOutput[94]}), .a ({key_s3[94], key_s2[94], key_s1[94], key_s0[94]}), .c ({new_AGEMA_signal_15378, new_AGEMA_signal_15377, new_AGEMA_signal_15376, KeyReg_Inst_ff_SDE_94_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_95_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14736, new_AGEMA_signal_14735, new_AGEMA_signal_14734, KeyExpansionOutput[95]}), .a ({key_s3[95], key_s2[95], key_s1[95], key_s0[95]}), .c ({new_AGEMA_signal_15384, new_AGEMA_signal_15383, new_AGEMA_signal_15382, KeyReg_Inst_ff_SDE_95_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_96_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, new_AGEMA_signal_12967, KeyExpansionOutput[96]}), .a ({key_s3[96], key_s2[96], key_s1[96], key_s0[96]}), .c ({new_AGEMA_signal_13398, new_AGEMA_signal_13397, new_AGEMA_signal_13396, KeyReg_Inst_ff_SDE_96_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_97_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13422, new_AGEMA_signal_13421, new_AGEMA_signal_13420, KeyExpansionOutput[97]}), .a ({key_s3[97], key_s2[97], key_s1[97], key_s0[97]}), .c ({new_AGEMA_signal_13914, new_AGEMA_signal_13913, new_AGEMA_signal_13912, KeyReg_Inst_ff_SDE_97_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_98_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, new_AGEMA_signal_13417, KeyExpansionOutput[98]}), .a ({key_s3[98], key_s2[98], key_s1[98], key_s0[98]}), .c ({new_AGEMA_signal_13920, new_AGEMA_signal_13919, new_AGEMA_signal_13918, KeyReg_Inst_ff_SDE_98_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_99_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13416, new_AGEMA_signal_13415, new_AGEMA_signal_13414, KeyExpansionOutput[99]}), .a ({key_s3[99], key_s2[99], key_s1[99], key_s0[99]}), .c ({new_AGEMA_signal_13926, new_AGEMA_signal_13925, new_AGEMA_signal_13924, KeyReg_Inst_ff_SDE_99_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_100_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13482, new_AGEMA_signal_13481, new_AGEMA_signal_13480, KeyExpansionOutput[100]}), .a ({key_s3[100], key_s2[100], key_s1[100], key_s0[100]}), .c ({new_AGEMA_signal_13932, new_AGEMA_signal_13931, new_AGEMA_signal_13930, KeyReg_Inst_ff_SDE_100_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_101_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, new_AGEMA_signal_13477, KeyExpansionOutput[101]}), .a ({key_s3[101], key_s2[101], key_s1[101], key_s0[101]}), .c ({new_AGEMA_signal_13938, new_AGEMA_signal_13937, new_AGEMA_signal_13936, KeyReg_Inst_ff_SDE_101_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_102_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13476, new_AGEMA_signal_13475, new_AGEMA_signal_13474, KeyExpansionOutput[102]}), .a ({key_s3[102], key_s2[102], key_s1[102], key_s0[102]}), .c ({new_AGEMA_signal_13944, new_AGEMA_signal_13943, new_AGEMA_signal_13942, KeyReg_Inst_ff_SDE_102_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_103_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, new_AGEMA_signal_13471, KeyExpansionOutput[103]}), .a ({key_s3[103], key_s2[103], key_s1[103], key_s0[103]}), .c ({new_AGEMA_signal_13950, new_AGEMA_signal_13949, new_AGEMA_signal_13948, KeyReg_Inst_ff_SDE_103_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_104_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12966, new_AGEMA_signal_12965, new_AGEMA_signal_12964, KeyExpansionOutput[104]}), .a ({key_s3[104], key_s2[104], key_s1[104], key_s0[104]}), .c ({new_AGEMA_signal_13404, new_AGEMA_signal_13403, new_AGEMA_signal_13402, KeyReg_Inst_ff_SDE_104_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_105_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13470, new_AGEMA_signal_13469, new_AGEMA_signal_13468, KeyExpansionOutput[105]}), .a ({key_s3[105], key_s2[105], key_s1[105], key_s0[105]}), .c ({new_AGEMA_signal_13956, new_AGEMA_signal_13955, new_AGEMA_signal_13954, KeyReg_Inst_ff_SDE_105_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_106_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, new_AGEMA_signal_13465, KeyExpansionOutput[106]}), .a ({key_s3[106], key_s2[106], key_s1[106], key_s0[106]}), .c ({new_AGEMA_signal_13962, new_AGEMA_signal_13961, new_AGEMA_signal_13960, KeyReg_Inst_ff_SDE_106_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_107_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13464, new_AGEMA_signal_13463, new_AGEMA_signal_13462, KeyExpansionOutput[107]}), .a ({key_s3[107], key_s2[107], key_s1[107], key_s0[107]}), .c ({new_AGEMA_signal_13968, new_AGEMA_signal_13967, new_AGEMA_signal_13966, KeyReg_Inst_ff_SDE_107_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_108_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, new_AGEMA_signal_13459, KeyExpansionOutput[108]}), .a ({key_s3[108], key_s2[108], key_s1[108], key_s0[108]}), .c ({new_AGEMA_signal_13974, new_AGEMA_signal_13973, new_AGEMA_signal_13972, KeyReg_Inst_ff_SDE_108_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_109_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13458, new_AGEMA_signal_13457, new_AGEMA_signal_13456, KeyExpansionOutput[109]}), .a ({key_s3[109], key_s2[109], key_s1[109], key_s0[109]}), .c ({new_AGEMA_signal_13980, new_AGEMA_signal_13979, new_AGEMA_signal_13978, KeyReg_Inst_ff_SDE_109_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_110_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, new_AGEMA_signal_13453, KeyExpansionOutput[110]}), .a ({key_s3[110], key_s2[110], key_s1[110], key_s0[110]}), .c ({new_AGEMA_signal_13986, new_AGEMA_signal_13985, new_AGEMA_signal_13984, KeyReg_Inst_ff_SDE_110_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_111_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13452, new_AGEMA_signal_13451, new_AGEMA_signal_13450, KeyExpansionOutput[111]}), .a ({key_s3[111], key_s2[111], key_s1[111], key_s0[111]}), .c ({new_AGEMA_signal_13992, new_AGEMA_signal_13991, new_AGEMA_signal_13990, KeyReg_Inst_ff_SDE_111_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_112_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, new_AGEMA_signal_12961, KeyExpansionOutput[112]}), .a ({key_s3[112], key_s2[112], key_s1[112], key_s0[112]}), .c ({new_AGEMA_signal_13410, new_AGEMA_signal_13409, new_AGEMA_signal_13408, KeyReg_Inst_ff_SDE_112_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_113_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, new_AGEMA_signal_13447, KeyExpansionOutput[113]}), .a ({key_s3[113], key_s2[113], key_s1[113], key_s0[113]}), .c ({new_AGEMA_signal_13998, new_AGEMA_signal_13997, new_AGEMA_signal_13996, KeyReg_Inst_ff_SDE_113_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_114_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13446, new_AGEMA_signal_13445, new_AGEMA_signal_13444, KeyExpansionOutput[114]}), .a ({key_s3[114], key_s2[114], key_s1[114], key_s0[114]}), .c ({new_AGEMA_signal_14004, new_AGEMA_signal_14003, new_AGEMA_signal_14002, KeyReg_Inst_ff_SDE_114_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_115_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, new_AGEMA_signal_13441, KeyExpansionOutput[115]}), .a ({key_s3[115], key_s2[115], key_s1[115], key_s0[115]}), .c ({new_AGEMA_signal_14010, new_AGEMA_signal_14009, new_AGEMA_signal_14008, KeyReg_Inst_ff_SDE_115_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_116_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13440, new_AGEMA_signal_13439, new_AGEMA_signal_13438, KeyExpansionOutput[116]}), .a ({key_s3[116], key_s2[116], key_s1[116], key_s0[116]}), .c ({new_AGEMA_signal_14016, new_AGEMA_signal_14015, new_AGEMA_signal_14014, KeyReg_Inst_ff_SDE_116_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_117_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, new_AGEMA_signal_13435, KeyExpansionOutput[117]}), .a ({key_s3[117], key_s2[117], key_s1[117], key_s0[117]}), .c ({new_AGEMA_signal_14022, new_AGEMA_signal_14021, new_AGEMA_signal_14020, KeyReg_Inst_ff_SDE_117_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_118_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13434, new_AGEMA_signal_13433, new_AGEMA_signal_13432, KeyExpansionOutput[118]}), .a ({key_s3[118], key_s2[118], key_s1[118], key_s0[118]}), .c ({new_AGEMA_signal_14028, new_AGEMA_signal_14027, new_AGEMA_signal_14026, KeyReg_Inst_ff_SDE_118_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_119_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, new_AGEMA_signal_13429, KeyExpansionOutput[119]}), .a ({key_s3[119], key_s2[119], key_s1[119], key_s0[119]}), .c ({new_AGEMA_signal_14034, new_AGEMA_signal_14033, new_AGEMA_signal_14032, KeyReg_Inst_ff_SDE_119_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_120_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_13428, new_AGEMA_signal_13427, new_AGEMA_signal_13426, KeyExpansionOutput[120]}), .a ({key_s3[120], key_s2[120], key_s1[120], key_s0[120]}), .c ({new_AGEMA_signal_14040, new_AGEMA_signal_14039, new_AGEMA_signal_14038, KeyReg_Inst_ff_SDE_120_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_121_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, new_AGEMA_signal_14125, KeyExpansionOutput[121]}), .a ({key_s3[121], key_s2[121], key_s1[121], key_s0[121]}), .c ({new_AGEMA_signal_14676, new_AGEMA_signal_14675, new_AGEMA_signal_14674, KeyReg_Inst_ff_SDE_121_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_122_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14124, new_AGEMA_signal_14123, new_AGEMA_signal_14122, KeyExpansionOutput[122]}), .a ({key_s3[122], key_s2[122], key_s1[122], key_s0[122]}), .c ({new_AGEMA_signal_14682, new_AGEMA_signal_14681, new_AGEMA_signal_14680, KeyReg_Inst_ff_SDE_122_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_123_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, new_AGEMA_signal_14119, KeyExpansionOutput[123]}), .a ({key_s3[123], key_s2[123], key_s1[123], key_s0[123]}), .c ({new_AGEMA_signal_14688, new_AGEMA_signal_14687, new_AGEMA_signal_14686, KeyReg_Inst_ff_SDE_123_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_124_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14118, new_AGEMA_signal_14117, new_AGEMA_signal_14116, KeyExpansionOutput[124]}), .a ({key_s3[124], key_s2[124], key_s1[124], key_s0[124]}), .c ({new_AGEMA_signal_14694, new_AGEMA_signal_14693, new_AGEMA_signal_14692, KeyReg_Inst_ff_SDE_124_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_125_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, new_AGEMA_signal_14113, KeyExpansionOutput[125]}), .a ({key_s3[125], key_s2[125], key_s1[125], key_s0[125]}), .c ({new_AGEMA_signal_14700, new_AGEMA_signal_14699, new_AGEMA_signal_14698, KeyReg_Inst_ff_SDE_125_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_126_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14112, new_AGEMA_signal_14111, new_AGEMA_signal_14110, KeyExpansionOutput[126]}), .a ({key_s3[126], key_s2[126], key_s1[126], key_s0[126]}), .c ({new_AGEMA_signal_14706, new_AGEMA_signal_14705, new_AGEMA_signal_14704, KeyReg_Inst_ff_SDE_126_next_state}) ) ;
    mux2_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_127_MUX_inst_U1 ( .s (reset), .b ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, new_AGEMA_signal_14107, KeyExpansionOutput[127]}), .a ({key_s3[127], key_s2[127], key_s1[127], key_s0[127]}), .c ({new_AGEMA_signal_14712, new_AGEMA_signal_14711, new_AGEMA_signal_14710, KeyReg_Inst_ff_SDE_127_next_state}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U128 ( .a ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}), .b ({new_AGEMA_signal_14718, new_AGEMA_signal_14717, new_AGEMA_signal_14716, KeyExpansionOutput[41]}), .c ({new_AGEMA_signal_15387, new_AGEMA_signal_15386, new_AGEMA_signal_15385, KeyExpansionOutput[9]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U127 ( .a ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .b ({new_AGEMA_signal_14046, new_AGEMA_signal_14045, new_AGEMA_signal_14044, KeyExpansionOutput[40]}), .c ({new_AGEMA_signal_14715, new_AGEMA_signal_14714, new_AGEMA_signal_14713, KeyExpansionOutput[8]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U126 ( .a ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}), .b ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, new_AGEMA_signal_14719, KeyExpansionOutput[39]}), .c ({new_AGEMA_signal_15390, new_AGEMA_signal_15389, new_AGEMA_signal_15388, KeyExpansionOutput[7]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U125 ( .a ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}), .b ({new_AGEMA_signal_14724, new_AGEMA_signal_14723, new_AGEMA_signal_14722, KeyExpansionOutput[38]}), .c ({new_AGEMA_signal_15393, new_AGEMA_signal_15392, new_AGEMA_signal_15391, KeyExpansionOutput[6]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U124 ( .a ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}), .b ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, new_AGEMA_signal_14725, KeyExpansionOutput[37]}), .c ({new_AGEMA_signal_15396, new_AGEMA_signal_15395, new_AGEMA_signal_15394, KeyExpansionOutput[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U123 ( .a ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}), .b ({new_AGEMA_signal_14730, new_AGEMA_signal_14729, new_AGEMA_signal_14728, KeyExpansionOutput[36]}), .c ({new_AGEMA_signal_15399, new_AGEMA_signal_15398, new_AGEMA_signal_15397, KeyExpansionOutput[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U122 ( .a ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundKey[41]}), .b ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, new_AGEMA_signal_14041, KeyExpansionOutput[73]}), .c ({new_AGEMA_signal_14718, new_AGEMA_signal_14717, new_AGEMA_signal_14716, KeyExpansionOutput[41]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U121 ( .a ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, RoundKey[73]}), .b ({new_AGEMA_signal_13470, new_AGEMA_signal_13469, new_AGEMA_signal_13468, KeyExpansionOutput[105]}), .c ({new_AGEMA_signal_14043, new_AGEMA_signal_14042, new_AGEMA_signal_14041, KeyExpansionOutput[73]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U120 ( .a ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, RoundKey[40]}), .b ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, new_AGEMA_signal_13411, KeyExpansionOutput[72]}), .c ({new_AGEMA_signal_14046, new_AGEMA_signal_14045, new_AGEMA_signal_14044, KeyExpansionOutput[40]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U119 ( .a ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, RoundKey[72]}), .b ({new_AGEMA_signal_12966, new_AGEMA_signal_12965, new_AGEMA_signal_12964, KeyExpansionOutput[104]}), .c ({new_AGEMA_signal_13413, new_AGEMA_signal_13412, new_AGEMA_signal_13411, KeyExpansionOutput[72]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U118 ( .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}), .b ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, new_AGEMA_signal_14731, KeyExpansionOutput[35]}), .c ({new_AGEMA_signal_15402, new_AGEMA_signal_15401, new_AGEMA_signal_15400, KeyExpansionOutput[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U117 ( .a ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKey[39]}), .b ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, new_AGEMA_signal_14047, KeyExpansionOutput[71]}), .c ({new_AGEMA_signal_14721, new_AGEMA_signal_14720, new_AGEMA_signal_14719, KeyExpansionOutput[39]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U116 ( .a ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, RoundKey[71]}), .b ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, new_AGEMA_signal_13471, KeyExpansionOutput[103]}), .c ({new_AGEMA_signal_14049, new_AGEMA_signal_14048, new_AGEMA_signal_14047, KeyExpansionOutput[71]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U115 ( .a ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundKey[38]}), .b ({new_AGEMA_signal_14052, new_AGEMA_signal_14051, new_AGEMA_signal_14050, KeyExpansionOutput[70]}), .c ({new_AGEMA_signal_14724, new_AGEMA_signal_14723, new_AGEMA_signal_14722, KeyExpansionOutput[38]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U114 ( .a ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, RoundKey[70]}), .b ({new_AGEMA_signal_13476, new_AGEMA_signal_13475, new_AGEMA_signal_13474, KeyExpansionOutput[102]}), .c ({new_AGEMA_signal_14052, new_AGEMA_signal_14051, new_AGEMA_signal_14050, KeyExpansionOutput[70]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U113 ( .a ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKey[37]}), .b ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, new_AGEMA_signal_14053, KeyExpansionOutput[69]}), .c ({new_AGEMA_signal_14727, new_AGEMA_signal_14726, new_AGEMA_signal_14725, KeyExpansionOutput[37]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U112 ( .a ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, RoundKey[69]}), .b ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, new_AGEMA_signal_13477, KeyExpansionOutput[101]}), .c ({new_AGEMA_signal_14055, new_AGEMA_signal_14054, new_AGEMA_signal_14053, KeyExpansionOutput[69]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U111 ( .a ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundKey[36]}), .b ({new_AGEMA_signal_14058, new_AGEMA_signal_14057, new_AGEMA_signal_14056, KeyExpansionOutput[68]}), .c ({new_AGEMA_signal_14730, new_AGEMA_signal_14729, new_AGEMA_signal_14728, KeyExpansionOutput[36]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U110 ( .a ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKey[68]}), .b ({new_AGEMA_signal_13482, new_AGEMA_signal_13481, new_AGEMA_signal_13480, KeyExpansionOutput[100]}), .c ({new_AGEMA_signal_14058, new_AGEMA_signal_14057, new_AGEMA_signal_14056, KeyExpansionOutput[68]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U109 ( .a ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKey[35]}), .b ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, new_AGEMA_signal_14059, KeyExpansionOutput[67]}), .c ({new_AGEMA_signal_14733, new_AGEMA_signal_14732, new_AGEMA_signal_14731, KeyExpansionOutput[35]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U108 ( .a ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, RoundKey[67]}), .b ({new_AGEMA_signal_13416, new_AGEMA_signal_13415, new_AGEMA_signal_13414, KeyExpansionOutput[99]}), .c ({new_AGEMA_signal_14061, new_AGEMA_signal_14060, new_AGEMA_signal_14059, KeyExpansionOutput[67]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U107 ( .a ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKey[99]}), .b ({new_AGEMA_signal_13050, new_AGEMA_signal_13049, new_AGEMA_signal_13048, KeyExpansionIns_tmp[3]}), .c ({new_AGEMA_signal_13416, new_AGEMA_signal_13415, new_AGEMA_signal_13414, KeyExpansionOutput[99]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U106 ( .a ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}), .b ({new_AGEMA_signal_15405, new_AGEMA_signal_15404, new_AGEMA_signal_15403, KeyExpansionOutput[63]}), .c ({new_AGEMA_signal_16032, new_AGEMA_signal_16031, new_AGEMA_signal_16030, KeyExpansionOutput[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U105 ( .a ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, RoundKey[63]}), .b ({new_AGEMA_signal_14736, new_AGEMA_signal_14735, new_AGEMA_signal_14734, KeyExpansionOutput[95]}), .c ({new_AGEMA_signal_15405, new_AGEMA_signal_15404, new_AGEMA_signal_15403, KeyExpansionOutput[63]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U104 ( .a ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKey[95]}), .b ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, new_AGEMA_signal_14107, KeyExpansionOutput[127]}), .c ({new_AGEMA_signal_14736, new_AGEMA_signal_14735, new_AGEMA_signal_14734, KeyExpansionOutput[95]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U103 ( .a ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}), .b ({new_AGEMA_signal_15408, new_AGEMA_signal_15407, new_AGEMA_signal_15406, KeyExpansionOutput[62]}), .c ({new_AGEMA_signal_16035, new_AGEMA_signal_16034, new_AGEMA_signal_16033, KeyExpansionOutput[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U102 ( .a ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, RoundKey[62]}), .b ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, new_AGEMA_signal_14737, KeyExpansionOutput[94]}), .c ({new_AGEMA_signal_15408, new_AGEMA_signal_15407, new_AGEMA_signal_15406, KeyExpansionOutput[62]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U101 ( .a ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, RoundKey[94]}), .b ({new_AGEMA_signal_14112, new_AGEMA_signal_14111, new_AGEMA_signal_14110, KeyExpansionOutput[126]}), .c ({new_AGEMA_signal_14739, new_AGEMA_signal_14738, new_AGEMA_signal_14737, KeyExpansionOutput[94]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U100 ( .a ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}), .b ({new_AGEMA_signal_14742, new_AGEMA_signal_14741, new_AGEMA_signal_14740, KeyExpansionOutput[34]}), .c ({new_AGEMA_signal_15411, new_AGEMA_signal_15410, new_AGEMA_signal_15409, KeyExpansionOutput[2]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U99 ( .a ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundKey[34]}), .b ({new_AGEMA_signal_14064, new_AGEMA_signal_14063, new_AGEMA_signal_14062, KeyExpansionOutput[66]}), .c ({new_AGEMA_signal_14742, new_AGEMA_signal_14741, new_AGEMA_signal_14740, KeyExpansionOutput[34]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U98 ( .a ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKey[66]}), .b ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, new_AGEMA_signal_13417, KeyExpansionOutput[98]}), .c ({new_AGEMA_signal_14064, new_AGEMA_signal_14063, new_AGEMA_signal_14062, KeyExpansionOutput[66]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U97 ( .a ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, RoundKey[98]}), .b ({new_AGEMA_signal_13053, new_AGEMA_signal_13052, new_AGEMA_signal_13051, KeyExpansionIns_tmp[2]}), .c ({new_AGEMA_signal_13419, new_AGEMA_signal_13418, new_AGEMA_signal_13417, KeyExpansionOutput[98]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U96 ( .a ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}), .b ({new_AGEMA_signal_15414, new_AGEMA_signal_15413, new_AGEMA_signal_15412, KeyExpansionOutput[61]}), .c ({new_AGEMA_signal_16038, new_AGEMA_signal_16037, new_AGEMA_signal_16036, KeyExpansionOutput[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U95 ( .a ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, RoundKey[61]}), .b ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, new_AGEMA_signal_14743, KeyExpansionOutput[93]}), .c ({new_AGEMA_signal_15414, new_AGEMA_signal_15413, new_AGEMA_signal_15412, KeyExpansionOutput[61]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U94 ( .a ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, RoundKey[93]}), .b ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, new_AGEMA_signal_14113, KeyExpansionOutput[125]}), .c ({new_AGEMA_signal_14745, new_AGEMA_signal_14744, new_AGEMA_signal_14743, KeyExpansionOutput[93]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U93 ( .a ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}), .b ({new_AGEMA_signal_15417, new_AGEMA_signal_15416, new_AGEMA_signal_15415, KeyExpansionOutput[60]}), .c ({new_AGEMA_signal_16041, new_AGEMA_signal_16040, new_AGEMA_signal_16039, KeyExpansionOutput[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U92 ( .a ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, RoundKey[60]}), .b ({new_AGEMA_signal_14748, new_AGEMA_signal_14747, new_AGEMA_signal_14746, KeyExpansionOutput[92]}), .c ({new_AGEMA_signal_15417, new_AGEMA_signal_15416, new_AGEMA_signal_15415, KeyExpansionOutput[60]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U91 ( .a ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, RoundKey[92]}), .b ({new_AGEMA_signal_14118, new_AGEMA_signal_14117, new_AGEMA_signal_14116, KeyExpansionOutput[124]}), .c ({new_AGEMA_signal_14748, new_AGEMA_signal_14747, new_AGEMA_signal_14746, KeyExpansionOutput[92]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U90 ( .a ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}), .b ({new_AGEMA_signal_15420, new_AGEMA_signal_15419, new_AGEMA_signal_15418, KeyExpansionOutput[59]}), .c ({new_AGEMA_signal_16044, new_AGEMA_signal_16043, new_AGEMA_signal_16042, KeyExpansionOutput[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U89 ( .a ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, RoundKey[59]}), .b ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, new_AGEMA_signal_14749, KeyExpansionOutput[91]}), .c ({new_AGEMA_signal_15420, new_AGEMA_signal_15419, new_AGEMA_signal_15418, KeyExpansionOutput[59]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U88 ( .a ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, RoundKey[91]}), .b ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, new_AGEMA_signal_14119, KeyExpansionOutput[123]}), .c ({new_AGEMA_signal_14751, new_AGEMA_signal_14750, new_AGEMA_signal_14749, KeyExpansionOutput[91]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U87 ( .a ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}), .b ({new_AGEMA_signal_15423, new_AGEMA_signal_15422, new_AGEMA_signal_15421, KeyExpansionOutput[58]}), .c ({new_AGEMA_signal_16047, new_AGEMA_signal_16046, new_AGEMA_signal_16045, KeyExpansionOutput[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U86 ( .a ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundKey[58]}), .b ({new_AGEMA_signal_14754, new_AGEMA_signal_14753, new_AGEMA_signal_14752, KeyExpansionOutput[90]}), .c ({new_AGEMA_signal_15423, new_AGEMA_signal_15422, new_AGEMA_signal_15421, KeyExpansionOutput[58]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U85 ( .a ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, RoundKey[90]}), .b ({new_AGEMA_signal_14124, new_AGEMA_signal_14123, new_AGEMA_signal_14122, KeyExpansionOutput[122]}), .c ({new_AGEMA_signal_14754, new_AGEMA_signal_14753, new_AGEMA_signal_14752, KeyExpansionOutput[90]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U84 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}), .b ({new_AGEMA_signal_15426, new_AGEMA_signal_15425, new_AGEMA_signal_15424, KeyExpansionOutput[57]}), .c ({new_AGEMA_signal_16050, new_AGEMA_signal_16049, new_AGEMA_signal_16048, KeyExpansionOutput[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U83 ( .a ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, RoundKey[57]}), .b ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, new_AGEMA_signal_14755, KeyExpansionOutput[89]}), .c ({new_AGEMA_signal_15426, new_AGEMA_signal_15425, new_AGEMA_signal_15424, KeyExpansionOutput[57]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U82 ( .a ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, RoundKey[89]}), .b ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, new_AGEMA_signal_14125, KeyExpansionOutput[121]}), .c ({new_AGEMA_signal_14757, new_AGEMA_signal_14756, new_AGEMA_signal_14755, KeyExpansionOutput[89]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U81 ( .a ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .b ({new_AGEMA_signal_14760, new_AGEMA_signal_14759, new_AGEMA_signal_14758, KeyExpansionOutput[56]}), .c ({new_AGEMA_signal_15429, new_AGEMA_signal_15428, new_AGEMA_signal_15427, KeyExpansionOutput[24]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U80 ( .a ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundKey[56]}), .b ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, new_AGEMA_signal_14065, KeyExpansionOutput[88]}), .c ({new_AGEMA_signal_14760, new_AGEMA_signal_14759, new_AGEMA_signal_14758, KeyExpansionOutput[56]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U79 ( .a ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, RoundKey[88]}), .b ({new_AGEMA_signal_13428, new_AGEMA_signal_13427, new_AGEMA_signal_13426, KeyExpansionOutput[120]}), .c ({new_AGEMA_signal_14067, new_AGEMA_signal_14066, new_AGEMA_signal_14065, KeyExpansionOutput[88]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U78 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}), .b ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, new_AGEMA_signal_14761, KeyExpansionOutput[55]}), .c ({new_AGEMA_signal_15432, new_AGEMA_signal_15431, new_AGEMA_signal_15430, KeyExpansionOutput[23]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U77 ( .a ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, RoundKey[55]}), .b ({new_AGEMA_signal_14070, new_AGEMA_signal_14069, new_AGEMA_signal_14068, KeyExpansionOutput[87]}), .c ({new_AGEMA_signal_14763, new_AGEMA_signal_14762, new_AGEMA_signal_14761, KeyExpansionOutput[55]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U76 ( .a ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, RoundKey[87]}), .b ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, new_AGEMA_signal_13429, KeyExpansionOutput[119]}), .c ({new_AGEMA_signal_14070, new_AGEMA_signal_14069, new_AGEMA_signal_14068, KeyExpansionOutput[87]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U75 ( .a ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}), .b ({new_AGEMA_signal_14766, new_AGEMA_signal_14765, new_AGEMA_signal_14764, KeyExpansionOutput[54]}), .c ({new_AGEMA_signal_15435, new_AGEMA_signal_15434, new_AGEMA_signal_15433, KeyExpansionOutput[22]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U74 ( .a ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundKey[54]}), .b ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, new_AGEMA_signal_14071, KeyExpansionOutput[86]}), .c ({new_AGEMA_signal_14766, new_AGEMA_signal_14765, new_AGEMA_signal_14764, KeyExpansionOutput[54]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U73 ( .a ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, RoundKey[86]}), .b ({new_AGEMA_signal_13434, new_AGEMA_signal_13433, new_AGEMA_signal_13432, KeyExpansionOutput[118]}), .c ({new_AGEMA_signal_14073, new_AGEMA_signal_14072, new_AGEMA_signal_14071, KeyExpansionOutput[86]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U72 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}), .b ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, new_AGEMA_signal_14767, KeyExpansionOutput[53]}), .c ({new_AGEMA_signal_15438, new_AGEMA_signal_15437, new_AGEMA_signal_15436, KeyExpansionOutput[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U71 ( .a ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, RoundKey[53]}), .b ({new_AGEMA_signal_14076, new_AGEMA_signal_14075, new_AGEMA_signal_14074, KeyExpansionOutput[85]}), .c ({new_AGEMA_signal_14769, new_AGEMA_signal_14768, new_AGEMA_signal_14767, KeyExpansionOutput[53]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U70 ( .a ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, RoundKey[85]}), .b ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, new_AGEMA_signal_13435, KeyExpansionOutput[117]}), .c ({new_AGEMA_signal_14076, new_AGEMA_signal_14075, new_AGEMA_signal_14074, KeyExpansionOutput[85]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U69 ( .a ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}), .b ({new_AGEMA_signal_14772, new_AGEMA_signal_14771, new_AGEMA_signal_14770, KeyExpansionOutput[52]}), .c ({new_AGEMA_signal_15441, new_AGEMA_signal_15440, new_AGEMA_signal_15439, KeyExpansionOutput[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U68 ( .a ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundKey[52]}), .b ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, new_AGEMA_signal_14077, KeyExpansionOutput[84]}), .c ({new_AGEMA_signal_14772, new_AGEMA_signal_14771, new_AGEMA_signal_14770, KeyExpansionOutput[52]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U67 ( .a ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, RoundKey[84]}), .b ({new_AGEMA_signal_13440, new_AGEMA_signal_13439, new_AGEMA_signal_13438, KeyExpansionOutput[116]}), .c ({new_AGEMA_signal_14079, new_AGEMA_signal_14078, new_AGEMA_signal_14077, KeyExpansionOutput[84]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U66 ( .a ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}), .b ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, new_AGEMA_signal_14773, KeyExpansionOutput[33]}), .c ({new_AGEMA_signal_15444, new_AGEMA_signal_15443, new_AGEMA_signal_15442, KeyExpansionOutput[1]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U65 ( .a ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, RoundKey[33]}), .b ({new_AGEMA_signal_14082, new_AGEMA_signal_14081, new_AGEMA_signal_14080, KeyExpansionOutput[65]}), .c ({new_AGEMA_signal_14775, new_AGEMA_signal_14774, new_AGEMA_signal_14773, KeyExpansionOutput[33]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U64 ( .a ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, RoundKey[65]}), .b ({new_AGEMA_signal_13422, new_AGEMA_signal_13421, new_AGEMA_signal_13420, KeyExpansionOutput[97]}), .c ({new_AGEMA_signal_14082, new_AGEMA_signal_14081, new_AGEMA_signal_14080, KeyExpansionOutput[65]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U63 ( .a ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKey[97]}), .b ({new_AGEMA_signal_13056, new_AGEMA_signal_13055, new_AGEMA_signal_13054, KeyExpansionIns_tmp[1]}), .c ({new_AGEMA_signal_13422, new_AGEMA_signal_13421, new_AGEMA_signal_13420, KeyExpansionOutput[97]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U62 ( .a ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}), .b ({new_AGEMA_signal_14778, new_AGEMA_signal_14777, new_AGEMA_signal_14776, KeyExpansionOutput[51]}), .c ({new_AGEMA_signal_15447, new_AGEMA_signal_15446, new_AGEMA_signal_15445, KeyExpansionOutput[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U61 ( .a ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, RoundKey[51]}), .b ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, new_AGEMA_signal_14083, KeyExpansionOutput[83]}), .c ({new_AGEMA_signal_14778, new_AGEMA_signal_14777, new_AGEMA_signal_14776, KeyExpansionOutput[51]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U60 ( .a ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, RoundKey[83]}), .b ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, new_AGEMA_signal_13441, KeyExpansionOutput[115]}), .c ({new_AGEMA_signal_14085, new_AGEMA_signal_14084, new_AGEMA_signal_14083, KeyExpansionOutput[83]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U59 ( .a ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}), .b ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, new_AGEMA_signal_14779, KeyExpansionOutput[50]}), .c ({new_AGEMA_signal_15450, new_AGEMA_signal_15449, new_AGEMA_signal_15448, KeyExpansionOutput[18]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U58 ( .a ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundKey[50]}), .b ({new_AGEMA_signal_14088, new_AGEMA_signal_14087, new_AGEMA_signal_14086, KeyExpansionOutput[82]}), .c ({new_AGEMA_signal_14781, new_AGEMA_signal_14780, new_AGEMA_signal_14779, KeyExpansionOutput[50]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U57 ( .a ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, RoundKey[82]}), .b ({new_AGEMA_signal_13446, new_AGEMA_signal_13445, new_AGEMA_signal_13444, KeyExpansionOutput[114]}), .c ({new_AGEMA_signal_14088, new_AGEMA_signal_14087, new_AGEMA_signal_14086, KeyExpansionOutput[82]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U56 ( .a ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}), .b ({new_AGEMA_signal_14784, new_AGEMA_signal_14783, new_AGEMA_signal_14782, KeyExpansionOutput[49]}), .c ({new_AGEMA_signal_15453, new_AGEMA_signal_15452, new_AGEMA_signal_15451, KeyExpansionOutput[17]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U55 ( .a ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundKey[49]}), .b ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, new_AGEMA_signal_14089, KeyExpansionOutput[81]}), .c ({new_AGEMA_signal_14784, new_AGEMA_signal_14783, new_AGEMA_signal_14782, KeyExpansionOutput[49]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U54 ( .a ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, RoundKey[81]}), .b ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, new_AGEMA_signal_13447, KeyExpansionOutput[113]}), .c ({new_AGEMA_signal_14091, new_AGEMA_signal_14090, new_AGEMA_signal_14089, KeyExpansionOutput[81]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U53 ( .a ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .b ({new_AGEMA_signal_14094, new_AGEMA_signal_14093, new_AGEMA_signal_14092, KeyExpansionOutput[48]}), .c ({new_AGEMA_signal_14787, new_AGEMA_signal_14786, new_AGEMA_signal_14785, KeyExpansionOutput[16]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U52 ( .a ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, RoundKey[48]}), .b ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, new_AGEMA_signal_13423, KeyExpansionOutput[80]}), .c ({new_AGEMA_signal_14094, new_AGEMA_signal_14093, new_AGEMA_signal_14092, KeyExpansionOutput[48]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U51 ( .a ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, RoundKey[80]}), .b ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, new_AGEMA_signal_12961, KeyExpansionOutput[112]}), .c ({new_AGEMA_signal_13425, new_AGEMA_signal_13424, new_AGEMA_signal_13423, KeyExpansionOutput[80]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U50 ( .a ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}), .b ({new_AGEMA_signal_14790, new_AGEMA_signal_14789, new_AGEMA_signal_14788, KeyExpansionOutput[47]}), .c ({new_AGEMA_signal_15456, new_AGEMA_signal_15455, new_AGEMA_signal_15454, KeyExpansionOutput[15]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U49 ( .a ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundKey[47]}), .b ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, new_AGEMA_signal_14095, KeyExpansionOutput[79]}), .c ({new_AGEMA_signal_14790, new_AGEMA_signal_14789, new_AGEMA_signal_14788, KeyExpansionOutput[47]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U48 ( .a ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, RoundKey[79]}), .b ({new_AGEMA_signal_13452, new_AGEMA_signal_13451, new_AGEMA_signal_13450, KeyExpansionOutput[111]}), .c ({new_AGEMA_signal_14097, new_AGEMA_signal_14096, new_AGEMA_signal_14095, KeyExpansionOutput[79]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U47 ( .a ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}), .b ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, new_AGEMA_signal_14791, KeyExpansionOutput[46]}), .c ({new_AGEMA_signal_15459, new_AGEMA_signal_15458, new_AGEMA_signal_15457, KeyExpansionOutput[14]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U46 ( .a ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, RoundKey[46]}), .b ({new_AGEMA_signal_14100, new_AGEMA_signal_14099, new_AGEMA_signal_14098, KeyExpansionOutput[78]}), .c ({new_AGEMA_signal_14793, new_AGEMA_signal_14792, new_AGEMA_signal_14791, KeyExpansionOutput[46]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U45 ( .a ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, RoundKey[78]}), .b ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, new_AGEMA_signal_13453, KeyExpansionOutput[110]}), .c ({new_AGEMA_signal_14100, new_AGEMA_signal_14099, new_AGEMA_signal_14098, KeyExpansionOutput[78]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U44 ( .a ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}), .b ({new_AGEMA_signal_14796, new_AGEMA_signal_14795, new_AGEMA_signal_14794, KeyExpansionOutput[45]}), .c ({new_AGEMA_signal_15462, new_AGEMA_signal_15461, new_AGEMA_signal_15460, KeyExpansionOutput[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U43 ( .a ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundKey[45]}), .b ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, new_AGEMA_signal_14101, KeyExpansionOutput[77]}), .c ({new_AGEMA_signal_14796, new_AGEMA_signal_14795, new_AGEMA_signal_14794, KeyExpansionOutput[45]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U42 ( .a ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, RoundKey[77]}), .b ({new_AGEMA_signal_13458, new_AGEMA_signal_13457, new_AGEMA_signal_13456, KeyExpansionOutput[109]}), .c ({new_AGEMA_signal_14103, new_AGEMA_signal_14102, new_AGEMA_signal_14101, KeyExpansionOutput[77]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U41 ( .a ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}), .b ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, new_AGEMA_signal_14797, KeyExpansionOutput[44]}), .c ({new_AGEMA_signal_15465, new_AGEMA_signal_15464, new_AGEMA_signal_15463, KeyExpansionOutput[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U40 ( .a ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, RoundKey[44]}), .b ({new_AGEMA_signal_14106, new_AGEMA_signal_14105, new_AGEMA_signal_14104, KeyExpansionOutput[76]}), .c ({new_AGEMA_signal_14799, new_AGEMA_signal_14798, new_AGEMA_signal_14797, KeyExpansionOutput[44]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U39 ( .a ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, RoundKey[76]}), .b ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, new_AGEMA_signal_13459, KeyExpansionOutput[108]}), .c ({new_AGEMA_signal_14106, new_AGEMA_signal_14105, new_AGEMA_signal_14104, KeyExpansionOutput[76]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U38 ( .a ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, RoundKey[127]}), .b ({new_AGEMA_signal_13488, new_AGEMA_signal_13487, new_AGEMA_signal_13486, KeyExpansionIns_tmp[31]}), .c ({new_AGEMA_signal_14109, new_AGEMA_signal_14108, new_AGEMA_signal_14107, KeyExpansionOutput[127]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U37 ( .a ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundKey[126]}), .b ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, new_AGEMA_signal_13489, KeyExpansionIns_tmp[30]}), .c ({new_AGEMA_signal_14112, new_AGEMA_signal_14111, new_AGEMA_signal_14110, KeyExpansionOutput[126]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U36 ( .a ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, RoundKey[125]}), .b ({new_AGEMA_signal_13494, new_AGEMA_signal_13493, new_AGEMA_signal_13492, KeyExpansionIns_tmp[29]}), .c ({new_AGEMA_signal_14115, new_AGEMA_signal_14114, new_AGEMA_signal_14113, KeyExpansionOutput[125]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U35 ( .a ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundKey[124]}), .b ({new_AGEMA_signal_13497, new_AGEMA_signal_13496, new_AGEMA_signal_13495, KeyExpansionIns_tmp[28]}), .c ({new_AGEMA_signal_14118, new_AGEMA_signal_14117, new_AGEMA_signal_14116, KeyExpansionOutput[124]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U34 ( .a ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, RoundKey[123]}), .b ({new_AGEMA_signal_13500, new_AGEMA_signal_13499, new_AGEMA_signal_13498, KeyExpansionIns_tmp[27]}), .c ({new_AGEMA_signal_14121, new_AGEMA_signal_14120, new_AGEMA_signal_14119, KeyExpansionOutput[123]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U33 ( .a ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundKey[122]}), .b ({new_AGEMA_signal_13503, new_AGEMA_signal_13502, new_AGEMA_signal_13501, KeyExpansionIns_tmp[26]}), .c ({new_AGEMA_signal_14124, new_AGEMA_signal_14123, new_AGEMA_signal_14122, KeyExpansionOutput[122]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U32 ( .a ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, RoundKey[121]}), .b ({new_AGEMA_signal_13506, new_AGEMA_signal_13505, new_AGEMA_signal_13504, KeyExpansionIns_tmp[25]}), .c ({new_AGEMA_signal_14127, new_AGEMA_signal_14126, new_AGEMA_signal_14125, KeyExpansionOutput[121]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U31 ( .a ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundKey[120]}), .b ({new_AGEMA_signal_12972, new_AGEMA_signal_12971, new_AGEMA_signal_12970, KeyExpansionIns_tmp[24]}), .c ({new_AGEMA_signal_13428, new_AGEMA_signal_13427, new_AGEMA_signal_13426, KeyExpansionOutput[120]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U30 ( .a ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}), .b ({new_AGEMA_signal_14802, new_AGEMA_signal_14801, new_AGEMA_signal_14800, KeyExpansionOutput[43]}), .c ({new_AGEMA_signal_15468, new_AGEMA_signal_15467, new_AGEMA_signal_15466, KeyExpansionOutput[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U29 ( .a ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundKey[43]}), .b ({new_AGEMA_signal_14130, new_AGEMA_signal_14129, new_AGEMA_signal_14128, KeyExpansionOutput[75]}), .c ({new_AGEMA_signal_14802, new_AGEMA_signal_14801, new_AGEMA_signal_14800, KeyExpansionOutput[43]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U28 ( .a ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, RoundKey[75]}), .b ({new_AGEMA_signal_13464, new_AGEMA_signal_13463, new_AGEMA_signal_13462, KeyExpansionOutput[107]}), .c ({new_AGEMA_signal_14130, new_AGEMA_signal_14129, new_AGEMA_signal_14128, KeyExpansionOutput[75]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U27 ( .a ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundKey[119]}), .b ({new_AGEMA_signal_12996, new_AGEMA_signal_12995, new_AGEMA_signal_12994, KeyExpansionIns_tmp[23]}), .c ({new_AGEMA_signal_13431, new_AGEMA_signal_13430, new_AGEMA_signal_13429, KeyExpansionOutput[119]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U26 ( .a ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, RoundKey[118]}), .b ({new_AGEMA_signal_12999, new_AGEMA_signal_12998, new_AGEMA_signal_12997, KeyExpansionIns_tmp[22]}), .c ({new_AGEMA_signal_13434, new_AGEMA_signal_13433, new_AGEMA_signal_13432, KeyExpansionOutput[118]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U25 ( .a ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundKey[117]}), .b ({new_AGEMA_signal_13002, new_AGEMA_signal_13001, new_AGEMA_signal_13000, KeyExpansionIns_tmp[21]}), .c ({new_AGEMA_signal_13437, new_AGEMA_signal_13436, new_AGEMA_signal_13435, KeyExpansionOutput[117]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U24 ( .a ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, RoundKey[116]}), .b ({new_AGEMA_signal_13005, new_AGEMA_signal_13004, new_AGEMA_signal_13003, KeyExpansionIns_tmp[20]}), .c ({new_AGEMA_signal_13440, new_AGEMA_signal_13439, new_AGEMA_signal_13438, KeyExpansionOutput[116]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U23 ( .a ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundKey[115]}), .b ({new_AGEMA_signal_13008, new_AGEMA_signal_13007, new_AGEMA_signal_13006, KeyExpansionIns_tmp[19]}), .c ({new_AGEMA_signal_13443, new_AGEMA_signal_13442, new_AGEMA_signal_13441, KeyExpansionOutput[115]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U22 ( .a ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, RoundKey[114]}), .b ({new_AGEMA_signal_13011, new_AGEMA_signal_13010, new_AGEMA_signal_13009, KeyExpansionIns_tmp[18]}), .c ({new_AGEMA_signal_13446, new_AGEMA_signal_13445, new_AGEMA_signal_13444, KeyExpansionOutput[114]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U21 ( .a ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundKey[113]}), .b ({new_AGEMA_signal_13014, new_AGEMA_signal_13013, new_AGEMA_signal_13012, KeyExpansionIns_tmp[17]}), .c ({new_AGEMA_signal_13449, new_AGEMA_signal_13448, new_AGEMA_signal_13447, KeyExpansionOutput[113]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U20 ( .a ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, RoundKey[112]}), .b ({new_AGEMA_signal_12366, new_AGEMA_signal_12365, new_AGEMA_signal_12364, KeyExpansionIns_tmp[16]}), .c ({new_AGEMA_signal_12963, new_AGEMA_signal_12962, new_AGEMA_signal_12961, KeyExpansionOutput[112]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U19 ( .a ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundKey[111]}), .b ({new_AGEMA_signal_13017, new_AGEMA_signal_13016, new_AGEMA_signal_13015, KeyExpansionIns_tmp[15]}), .c ({new_AGEMA_signal_13452, new_AGEMA_signal_13451, new_AGEMA_signal_13450, KeyExpansionOutput[111]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U18 ( .a ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, RoundKey[110]}), .b ({new_AGEMA_signal_13020, new_AGEMA_signal_13019, new_AGEMA_signal_13018, KeyExpansionIns_tmp[14]}), .c ({new_AGEMA_signal_13455, new_AGEMA_signal_13454, new_AGEMA_signal_13453, KeyExpansionOutput[110]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U17 ( .a ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}), .b ({new_AGEMA_signal_14805, new_AGEMA_signal_14804, new_AGEMA_signal_14803, KeyExpansionOutput[42]}), .c ({new_AGEMA_signal_15471, new_AGEMA_signal_15470, new_AGEMA_signal_15469, KeyExpansionOutput[10]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U16 ( .a ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, RoundKey[42]}), .b ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, new_AGEMA_signal_14131, KeyExpansionOutput[74]}), .c ({new_AGEMA_signal_14805, new_AGEMA_signal_14804, new_AGEMA_signal_14803, KeyExpansionOutput[42]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U15 ( .a ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, RoundKey[74]}), .b ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, new_AGEMA_signal_13465, KeyExpansionOutput[106]}), .c ({new_AGEMA_signal_14133, new_AGEMA_signal_14132, new_AGEMA_signal_14131, KeyExpansionOutput[74]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U14 ( .a ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, RoundKey[109]}), .b ({new_AGEMA_signal_13023, new_AGEMA_signal_13022, new_AGEMA_signal_13021, KeyExpansionIns_tmp[13]}), .c ({new_AGEMA_signal_13458, new_AGEMA_signal_13457, new_AGEMA_signal_13456, KeyExpansionOutput[109]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U13 ( .a ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundKey[108]}), .b ({new_AGEMA_signal_13026, new_AGEMA_signal_13025, new_AGEMA_signal_13024, KeyExpansionIns_tmp[12]}), .c ({new_AGEMA_signal_13461, new_AGEMA_signal_13460, new_AGEMA_signal_13459, KeyExpansionOutput[108]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U12 ( .a ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, RoundKey[107]}), .b ({new_AGEMA_signal_13029, new_AGEMA_signal_13028, new_AGEMA_signal_13027, KeyExpansionIns_tmp[11]}), .c ({new_AGEMA_signal_13464, new_AGEMA_signal_13463, new_AGEMA_signal_13462, KeyExpansionOutput[107]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U11 ( .a ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundKey[106]}), .b ({new_AGEMA_signal_13032, new_AGEMA_signal_13031, new_AGEMA_signal_13030, KeyExpansionIns_tmp[10]}), .c ({new_AGEMA_signal_13467, new_AGEMA_signal_13466, new_AGEMA_signal_13465, KeyExpansionOutput[106]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U10 ( .a ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, RoundKey[105]}), .b ({new_AGEMA_signal_13035, new_AGEMA_signal_13034, new_AGEMA_signal_13033, KeyExpansionIns_tmp[9]}), .c ({new_AGEMA_signal_13470, new_AGEMA_signal_13469, new_AGEMA_signal_13468, KeyExpansionOutput[105]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U9 ( .a ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundKey[104]}), .b ({new_AGEMA_signal_12399, new_AGEMA_signal_12398, new_AGEMA_signal_12397, KeyExpansionIns_tmp[8]}), .c ({new_AGEMA_signal_12966, new_AGEMA_signal_12965, new_AGEMA_signal_12964, KeyExpansionOutput[104]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U8 ( .a ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, RoundKey[103]}), .b ({new_AGEMA_signal_13038, new_AGEMA_signal_13037, new_AGEMA_signal_13036, KeyExpansionIns_tmp[7]}), .c ({new_AGEMA_signal_13473, new_AGEMA_signal_13472, new_AGEMA_signal_13471, KeyExpansionOutput[103]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U7 ( .a ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundKey[102]}), .b ({new_AGEMA_signal_13041, new_AGEMA_signal_13040, new_AGEMA_signal_13039, KeyExpansionIns_tmp[6]}), .c ({new_AGEMA_signal_13476, new_AGEMA_signal_13475, new_AGEMA_signal_13474, KeyExpansionOutput[102]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U6 ( .a ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, RoundKey[101]}), .b ({new_AGEMA_signal_13044, new_AGEMA_signal_13043, new_AGEMA_signal_13042, KeyExpansionIns_tmp[5]}), .c ({new_AGEMA_signal_13479, new_AGEMA_signal_13478, new_AGEMA_signal_13477, KeyExpansionOutput[101]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U5 ( .a ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundKey[100]}), .b ({new_AGEMA_signal_13047, new_AGEMA_signal_13046, new_AGEMA_signal_13045, KeyExpansionIns_tmp[4]}), .c ({new_AGEMA_signal_13482, new_AGEMA_signal_13481, new_AGEMA_signal_13480, KeyExpansionOutput[100]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U4 ( .a ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .b ({new_AGEMA_signal_14136, new_AGEMA_signal_14135, new_AGEMA_signal_14134, KeyExpansionOutput[32]}), .c ({new_AGEMA_signal_14808, new_AGEMA_signal_14807, new_AGEMA_signal_14806, KeyExpansionOutput[0]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U3 ( .a ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundKey[32]}), .b ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, new_AGEMA_signal_13483, KeyExpansionOutput[64]}), .c ({new_AGEMA_signal_14136, new_AGEMA_signal_14135, new_AGEMA_signal_14134, KeyExpansionOutput[32]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U2 ( .a ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKey[64]}), .b ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, new_AGEMA_signal_12967, KeyExpansionOutput[96]}), .c ({new_AGEMA_signal_13485, new_AGEMA_signal_13484, new_AGEMA_signal_13483, KeyExpansionOutput[64]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_U1 ( .a ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, RoundKey[96]}), .b ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, new_AGEMA_signal_12430, KeyExpansionIns_tmp[0]}), .c ({new_AGEMA_signal_12969, new_AGEMA_signal_12968, new_AGEMA_signal_12967, KeyExpansionOutput[96]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U8 ( .a ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, new_AGEMA_signal_12973, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}), .b ({1'b0, 1'b0, 1'b0, n283}), .c ({new_AGEMA_signal_13488, new_AGEMA_signal_13487, new_AGEMA_signal_13486, KeyExpansionIns_tmp[31]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U7 ( .a ({new_AGEMA_signal_12978, new_AGEMA_signal_12977, new_AGEMA_signal_12976, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}), .b ({1'b0, 1'b0, 1'b0, n285}), .c ({new_AGEMA_signal_13491, new_AGEMA_signal_13490, new_AGEMA_signal_13489, KeyExpansionIns_tmp[30]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U6 ( .a ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, new_AGEMA_signal_12979, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}), .b ({1'b0, 1'b0, 1'b0, Rcon[5]}), .c ({new_AGEMA_signal_13494, new_AGEMA_signal_13493, new_AGEMA_signal_13492, KeyExpansionIns_tmp[29]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U5 ( .a ({new_AGEMA_signal_12984, new_AGEMA_signal_12983, new_AGEMA_signal_12982, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}), .b ({1'b0, 1'b0, 1'b0, Rcon[4]}), .c ({new_AGEMA_signal_13497, new_AGEMA_signal_13496, new_AGEMA_signal_13495, KeyExpansionIns_tmp[28]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U4 ( .a ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, new_AGEMA_signal_12985, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}), .b ({1'b0, 1'b0, 1'b0, Rcon[3]}), .c ({new_AGEMA_signal_13500, new_AGEMA_signal_13499, new_AGEMA_signal_13498, KeyExpansionIns_tmp[27]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U3 ( .a ({new_AGEMA_signal_12990, new_AGEMA_signal_12989, new_AGEMA_signal_12988, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}), .b ({1'b0, 1'b0, 1'b0, Rcon[2]}), .c ({new_AGEMA_signal_13503, new_AGEMA_signal_13502, new_AGEMA_signal_13501, KeyExpansionIns_tmp[26]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U2 ( .a ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, new_AGEMA_signal_12991, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}), .b ({1'b0, 1'b0, 1'b0, Rcon[1]}), .c ({new_AGEMA_signal_13506, new_AGEMA_signal_13505, new_AGEMA_signal_13504, KeyExpansionIns_tmp[25]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_U1 ( .a ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, new_AGEMA_signal_12331, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}), .b ({1'b0, 1'b0, 1'b0, Rcon[0]}), .c ({new_AGEMA_signal_12972, new_AGEMA_signal_12971, new_AGEMA_signal_12970, KeyExpansionIns_tmp[24]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M46_U1 ( .a ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, new_AGEMA_signal_9730, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_6303, new_AGEMA_signal_6302, new_AGEMA_signal_6301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T6}), .clk (clk), .r ({Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648]}), .c ({new_AGEMA_signal_10446, new_AGEMA_signal_10445, new_AGEMA_signal_10444, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M47_U1 ( .a ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6783, new_AGEMA_signal_6782, new_AGEMA_signal_6781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T8}), .clk (clk), .r ({Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654]}), .c ({new_AGEMA_signal_9735, new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M48_U1 ( .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}), .clk (clk), .r ({Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660]}), .c ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, new_AGEMA_signal_9736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M49_U1 ( .a ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_6315, new_AGEMA_signal_6314, new_AGEMA_signal_6313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T16}), .clk (clk), .r ({Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666]}), .c ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M50_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6306, new_AGEMA_signal_6305, new_AGEMA_signal_6304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T9}), .clk (clk), .r ({Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672]}), .c ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M51_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6792, new_AGEMA_signal_6791, new_AGEMA_signal_6790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T17}), .clk (clk), .r ({Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678]}), .c ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, new_AGEMA_signal_9742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M52_U1 ( .a ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_6312, new_AGEMA_signal_6311, new_AGEMA_signal_6310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T15}), .clk (clk), .r ({Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684]}), .c ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, new_AGEMA_signal_10450, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M53_U1 ( .a ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, new_AGEMA_signal_10441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_6324, new_AGEMA_signal_6323, new_AGEMA_signal_6322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T27}), .clk (clk), .r ({Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690]}), .c ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, new_AGEMA_signal_11161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M54_U1 ( .a ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_6786, new_AGEMA_signal_6785, new_AGEMA_signal_6784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T10}), .clk (clk), .r ({Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696]}), .c ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, new_AGEMA_signal_10453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M55_U1 ( .a ({new_AGEMA_signal_9732, new_AGEMA_signal_9731, new_AGEMA_signal_9730, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M44}), .b ({new_AGEMA_signal_6309, new_AGEMA_signal_6308, new_AGEMA_signal_6307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T13}), .clk (clk), .r ({Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702]}), .c ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, new_AGEMA_signal_10456, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M56_U1 ( .a ({new_AGEMA_signal_9492, new_AGEMA_signal_9491, new_AGEMA_signal_9490, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M40}), .b ({new_AGEMA_signal_6798, new_AGEMA_signal_6797, new_AGEMA_signal_6796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T23}), .clk (clk), .r ({Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708]}), .c ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M57_U1 ( .a ({new_AGEMA_signal_9489, new_AGEMA_signal_9488, new_AGEMA_signal_9487, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M39}), .b ({new_AGEMA_signal_6318, new_AGEMA_signal_6317, new_AGEMA_signal_6316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T19}), .clk (clk), .r ({Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714]}), .c ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, new_AGEMA_signal_9748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M58_U1 ( .a ({new_AGEMA_signal_9729, new_AGEMA_signal_9728, new_AGEMA_signal_9727, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M43}), .b ({new_AGEMA_signal_5709, new_AGEMA_signal_5708, new_AGEMA_signal_5707, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T3}), .clk (clk), .r ({Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720]}), .c ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M59_U1 ( .a ({new_AGEMA_signal_9486, new_AGEMA_signal_9485, new_AGEMA_signal_9484, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M38}), .b ({new_AGEMA_signal_6321, new_AGEMA_signal_6320, new_AGEMA_signal_6319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T22}), .clk (clk), .r ({Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726]}), .c ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M60_U1 ( .a ({new_AGEMA_signal_9483, new_AGEMA_signal_9482, new_AGEMA_signal_9481, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M37}), .b ({new_AGEMA_signal_6795, new_AGEMA_signal_6794, new_AGEMA_signal_6793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T20}), .clk (clk), .r ({Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732]}), .c ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, new_AGEMA_signal_9754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M61_U1 ( .a ({new_AGEMA_signal_9726, new_AGEMA_signal_9725, new_AGEMA_signal_9724, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M42}), .b ({new_AGEMA_signal_5703, new_AGEMA_signal_5702, new_AGEMA_signal_5701, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T1}), .clk (clk), .r ({Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738]}), .c ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M62_U1 ( .a ({new_AGEMA_signal_10443, new_AGEMA_signal_10442, new_AGEMA_signal_10441, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M45}), .b ({new_AGEMA_signal_5712, new_AGEMA_signal_5711, new_AGEMA_signal_5710, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T4}), .clk (clk), .r ({Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744]}), .c ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, new_AGEMA_signal_11164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_AND_M63_U1 ( .a ({new_AGEMA_signal_9723, new_AGEMA_signal_9722, new_AGEMA_signal_9721, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M41}), .b ({new_AGEMA_signal_5706, new_AGEMA_signal_5705, new_AGEMA_signal_5704, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_T2}), .clk (clk), .r ({Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750]}), .c ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L0_U1 ( .a ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .b ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, new_AGEMA_signal_11164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .c ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L1_U1 ( .a ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .c ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L2_U1 ( .a ({new_AGEMA_signal_10446, new_AGEMA_signal_10445, new_AGEMA_signal_10444, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, new_AGEMA_signal_9736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .c ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, new_AGEMA_signal_11167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L3_U1 ( .a ({new_AGEMA_signal_9735, new_AGEMA_signal_9734, new_AGEMA_signal_9733, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M47}), .b ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, new_AGEMA_signal_10456, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .c ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, new_AGEMA_signal_11170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L4_U1 ( .a ({new_AGEMA_signal_10455, new_AGEMA_signal_10454, new_AGEMA_signal_10453, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M54}), .b ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .c ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, new_AGEMA_signal_11173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L5_U1 ( .a ({new_AGEMA_signal_10449, new_AGEMA_signal_10448, new_AGEMA_signal_10447, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M49}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, new_AGEMA_signal_11176, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L6_U1 ( .a ({new_AGEMA_signal_11166, new_AGEMA_signal_11165, new_AGEMA_signal_11164, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M62}), .b ({new_AGEMA_signal_11178, new_AGEMA_signal_11177, new_AGEMA_signal_11176, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L5}), .c ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L7_U1 ( .a ({new_AGEMA_signal_10446, new_AGEMA_signal_10445, new_AGEMA_signal_10444, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M46}), .b ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, new_AGEMA_signal_11170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .c ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L8_U1 ( .a ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, new_AGEMA_signal_9742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .b ({new_AGEMA_signal_9753, new_AGEMA_signal_9752, new_AGEMA_signal_9751, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M59}), .c ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L9_U1 ( .a ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, new_AGEMA_signal_10450, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, new_AGEMA_signal_11161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .c ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, new_AGEMA_signal_11770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L10_U1 ( .a ({new_AGEMA_signal_11163, new_AGEMA_signal_11162, new_AGEMA_signal_11161, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M53}), .b ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, new_AGEMA_signal_11173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L11_U1 ( .a ({new_AGEMA_signal_9756, new_AGEMA_signal_9755, new_AGEMA_signal_9754, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M60}), .b ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, new_AGEMA_signal_11167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, new_AGEMA_signal_11776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L12_U1 ( .a ({new_AGEMA_signal_9738, new_AGEMA_signal_9737, new_AGEMA_signal_9736, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M48}), .b ({new_AGEMA_signal_9744, new_AGEMA_signal_9743, new_AGEMA_signal_9742, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M51}), .c ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, new_AGEMA_signal_10474, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L13_U1 ( .a ({new_AGEMA_signal_9741, new_AGEMA_signal_9740, new_AGEMA_signal_9739, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M50}), .b ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, new_AGEMA_signal_12301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L14_U1 ( .a ({new_AGEMA_signal_10452, new_AGEMA_signal_10451, new_AGEMA_signal_10450, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M52}), .b ({new_AGEMA_signal_10464, new_AGEMA_signal_10463, new_AGEMA_signal_10462, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M61}), .c ({new_AGEMA_signal_11181, new_AGEMA_signal_11180, new_AGEMA_signal_11179, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L15_U1 ( .a ({new_AGEMA_signal_10458, new_AGEMA_signal_10457, new_AGEMA_signal_10456, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M55}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, new_AGEMA_signal_11182, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L16_U1 ( .a ({new_AGEMA_signal_9747, new_AGEMA_signal_9746, new_AGEMA_signal_9745, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M56}), .b ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .c ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, new_AGEMA_signal_12304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L17_U1 ( .a ({new_AGEMA_signal_9750, new_AGEMA_signal_9749, new_AGEMA_signal_9748, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M57}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_11187, new_AGEMA_signal_11186, new_AGEMA_signal_11185, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L18_U1 ( .a ({new_AGEMA_signal_10461, new_AGEMA_signal_10460, new_AGEMA_signal_10459, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M58}), .b ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .c ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, new_AGEMA_signal_11188, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L19_U1 ( .a ({new_AGEMA_signal_10467, new_AGEMA_signal_10466, new_AGEMA_signal_10465, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_M63}), .b ({new_AGEMA_signal_11175, new_AGEMA_signal_11174, new_AGEMA_signal_11173, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L4}), .c ({new_AGEMA_signal_11781, new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L20_U1 ( .a ({new_AGEMA_signal_11763, new_AGEMA_signal_11762, new_AGEMA_signal_11761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L0}), .b ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .c ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, new_AGEMA_signal_12307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L21_U1 ( .a ({new_AGEMA_signal_10470, new_AGEMA_signal_10469, new_AGEMA_signal_10468, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L1}), .b ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .c ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, new_AGEMA_signal_12310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L22_U1 ( .a ({new_AGEMA_signal_11172, new_AGEMA_signal_11171, new_AGEMA_signal_11170, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L3}), .b ({new_AGEMA_signal_10476, new_AGEMA_signal_10475, new_AGEMA_signal_10474, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L12}), .c ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, new_AGEMA_signal_11782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L23_U1 ( .a ({new_AGEMA_signal_11190, new_AGEMA_signal_11189, new_AGEMA_signal_11188, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L18}), .b ({new_AGEMA_signal_11169, new_AGEMA_signal_11168, new_AGEMA_signal_11167, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L2}), .c ({new_AGEMA_signal_11787, new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L24_U1 ( .a ({new_AGEMA_signal_11184, new_AGEMA_signal_11183, new_AGEMA_signal_11182, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L15}), .b ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, new_AGEMA_signal_11770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12315, new_AGEMA_signal_12314, new_AGEMA_signal_12313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L25_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12318, new_AGEMA_signal_12317, new_AGEMA_signal_12316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L26_U1 ( .a ({new_AGEMA_signal_11769, new_AGEMA_signal_11768, new_AGEMA_signal_11767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L7}), .b ({new_AGEMA_signal_11772, new_AGEMA_signal_11771, new_AGEMA_signal_11770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L9}), .c ({new_AGEMA_signal_12321, new_AGEMA_signal_12320, new_AGEMA_signal_12319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L27_U1 ( .a ({new_AGEMA_signal_10473, new_AGEMA_signal_10472, new_AGEMA_signal_10471, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L8}), .b ({new_AGEMA_signal_11775, new_AGEMA_signal_11774, new_AGEMA_signal_11773, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L10}), .c ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, new_AGEMA_signal_12322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L28_U1 ( .a ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, new_AGEMA_signal_11776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11181, new_AGEMA_signal_11180, new_AGEMA_signal_11179, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L14}), .c ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, new_AGEMA_signal_12325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_L29_U1 ( .a ({new_AGEMA_signal_11778, new_AGEMA_signal_11777, new_AGEMA_signal_11776, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L11}), .b ({new_AGEMA_signal_11187, new_AGEMA_signal_11186, new_AGEMA_signal_11185, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L17}), .c ({new_AGEMA_signal_12330, new_AGEMA_signal_12329, new_AGEMA_signal_12328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S0_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12315, new_AGEMA_signal_12314, new_AGEMA_signal_12313, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L24}), .c ({new_AGEMA_signal_12975, new_AGEMA_signal_12974, new_AGEMA_signal_12973, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__7_}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S1_U1 ( .a ({new_AGEMA_signal_12306, new_AGEMA_signal_12305, new_AGEMA_signal_12304, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L16}), .b ({new_AGEMA_signal_12321, new_AGEMA_signal_12320, new_AGEMA_signal_12319, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L26}), .c ({new_AGEMA_signal_12978, new_AGEMA_signal_12977, new_AGEMA_signal_12976, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__6_}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S2_U1 ( .a ({new_AGEMA_signal_11781, new_AGEMA_signal_11780, new_AGEMA_signal_11779, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L19}), .b ({new_AGEMA_signal_12327, new_AGEMA_signal_12326, new_AGEMA_signal_12325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L28}), .c ({new_AGEMA_signal_12981, new_AGEMA_signal_12980, new_AGEMA_signal_12979, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__5_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S3_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_12312, new_AGEMA_signal_12311, new_AGEMA_signal_12310, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L21}), .c ({new_AGEMA_signal_12984, new_AGEMA_signal_12983, new_AGEMA_signal_12982, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__4_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S4_U1 ( .a ({new_AGEMA_signal_12309, new_AGEMA_signal_12308, new_AGEMA_signal_12307, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L20}), .b ({new_AGEMA_signal_11784, new_AGEMA_signal_11783, new_AGEMA_signal_11782, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L22}), .c ({new_AGEMA_signal_12987, new_AGEMA_signal_12986, new_AGEMA_signal_12985, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__3_}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S5_U1 ( .a ({new_AGEMA_signal_12318, new_AGEMA_signal_12317, new_AGEMA_signal_12316, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L25}), .b ({new_AGEMA_signal_12330, new_AGEMA_signal_12329, new_AGEMA_signal_12328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L29}), .c ({new_AGEMA_signal_12990, new_AGEMA_signal_12989, new_AGEMA_signal_12988, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__2_}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S6_U1 ( .a ({new_AGEMA_signal_12303, new_AGEMA_signal_12302, new_AGEMA_signal_12301, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L13}), .b ({new_AGEMA_signal_12324, new_AGEMA_signal_12323, new_AGEMA_signal_12322, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L27}), .c ({new_AGEMA_signal_12993, new_AGEMA_signal_12992, new_AGEMA_signal_12991, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__1_}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_XOR_S7_U1 ( .a ({new_AGEMA_signal_11766, new_AGEMA_signal_11765, new_AGEMA_signal_11764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L6}), .b ({new_AGEMA_signal_11787, new_AGEMA_signal_11786, new_AGEMA_signal_11785, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_0_L23}), .c ({new_AGEMA_signal_12333, new_AGEMA_signal_12332, new_AGEMA_signal_12331, KeyExpansionIns_KeySchedCoreInst_OutBytes_0__0_}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M46_U1 ( .a ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, new_AGEMA_signal_9766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_6327, new_AGEMA_signal_6326, new_AGEMA_signal_6325, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T6}), .clk (clk), .r ({Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756]}), .c ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, new_AGEMA_signal_10480, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M47_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6822, new_AGEMA_signal_6821, new_AGEMA_signal_6820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T8}), .clk (clk), .r ({Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762]}), .c ({new_AGEMA_signal_9771, new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M48_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}), .clk (clk), .r ({Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768]}), .c ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, new_AGEMA_signal_9772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M49_U1 ( .a ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_6339, new_AGEMA_signal_6338, new_AGEMA_signal_6337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T16}), .clk (clk), .r ({Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774]}), .c ({new_AGEMA_signal_10485, new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M50_U1 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6330, new_AGEMA_signal_6329, new_AGEMA_signal_6328, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T9}), .clk (clk), .r ({Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780]}), .c ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M51_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6831, new_AGEMA_signal_6830, new_AGEMA_signal_6829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T17}), .clk (clk), .r ({Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786]}), .c ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, new_AGEMA_signal_9778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M52_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_6336, new_AGEMA_signal_6335, new_AGEMA_signal_6334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T15}), .clk (clk), .r ({Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792]}), .c ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, new_AGEMA_signal_10486, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M53_U1 ( .a ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_6348, new_AGEMA_signal_6347, new_AGEMA_signal_6346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T27}), .clk (clk), .r ({Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798]}), .c ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, new_AGEMA_signal_11191, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M54_U1 ( .a ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_6825, new_AGEMA_signal_6824, new_AGEMA_signal_6823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T10}), .clk (clk), .r ({Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804]}), .c ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M55_U1 ( .a ({new_AGEMA_signal_9768, new_AGEMA_signal_9767, new_AGEMA_signal_9766, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M44}), .b ({new_AGEMA_signal_6333, new_AGEMA_signal_6332, new_AGEMA_signal_6331, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T13}), .clk (clk), .r ({Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810]}), .c ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, new_AGEMA_signal_10492, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M56_U1 ( .a ({new_AGEMA_signal_9504, new_AGEMA_signal_9503, new_AGEMA_signal_9502, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M40}), .b ({new_AGEMA_signal_6837, new_AGEMA_signal_6836, new_AGEMA_signal_6835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T23}), .clk (clk), .r ({Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816]}), .c ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M57_U1 ( .a ({new_AGEMA_signal_9501, new_AGEMA_signal_9500, new_AGEMA_signal_9499, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M39}), .b ({new_AGEMA_signal_6342, new_AGEMA_signal_6341, new_AGEMA_signal_6340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T19}), .clk (clk), .r ({Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822]}), .c ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, new_AGEMA_signal_9784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M58_U1 ( .a ({new_AGEMA_signal_9765, new_AGEMA_signal_9764, new_AGEMA_signal_9763, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M43}), .b ({new_AGEMA_signal_5739, new_AGEMA_signal_5738, new_AGEMA_signal_5737, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T3}), .clk (clk), .r ({Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828]}), .c ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M59_U1 ( .a ({new_AGEMA_signal_9498, new_AGEMA_signal_9497, new_AGEMA_signal_9496, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M38}), .b ({new_AGEMA_signal_6345, new_AGEMA_signal_6344, new_AGEMA_signal_6343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T22}), .clk (clk), .r ({Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834]}), .c ({new_AGEMA_signal_9789, new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M60_U1 ( .a ({new_AGEMA_signal_9495, new_AGEMA_signal_9494, new_AGEMA_signal_9493, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M37}), .b ({new_AGEMA_signal_6834, new_AGEMA_signal_6833, new_AGEMA_signal_6832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T20}), .clk (clk), .r ({Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840]}), .c ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, new_AGEMA_signal_9790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M61_U1 ( .a ({new_AGEMA_signal_9762, new_AGEMA_signal_9761, new_AGEMA_signal_9760, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M42}), .b ({new_AGEMA_signal_5733, new_AGEMA_signal_5732, new_AGEMA_signal_5731, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T1}), .clk (clk), .r ({Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846]}), .c ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M62_U1 ( .a ({new_AGEMA_signal_10479, new_AGEMA_signal_10478, new_AGEMA_signal_10477, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M45}), .b ({new_AGEMA_signal_5742, new_AGEMA_signal_5741, new_AGEMA_signal_5740, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T4}), .clk (clk), .r ({Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852]}), .c ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, new_AGEMA_signal_11194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_AND_M63_U1 ( .a ({new_AGEMA_signal_9759, new_AGEMA_signal_9758, new_AGEMA_signal_9757, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M41}), .b ({new_AGEMA_signal_5736, new_AGEMA_signal_5735, new_AGEMA_signal_5734, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_T2}), .clk (clk), .r ({Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858]}), .c ({new_AGEMA_signal_10503, new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L0_U1 ( .a ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .b ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, new_AGEMA_signal_11194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .c ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L1_U1 ( .a ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .c ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L2_U1 ( .a ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, new_AGEMA_signal_10480, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, new_AGEMA_signal_9772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .c ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, new_AGEMA_signal_11197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L3_U1 ( .a ({new_AGEMA_signal_9771, new_AGEMA_signal_9770, new_AGEMA_signal_9769, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M47}), .b ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, new_AGEMA_signal_10492, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .c ({new_AGEMA_signal_11202, new_AGEMA_signal_11201, new_AGEMA_signal_11200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L4_U1 ( .a ({new_AGEMA_signal_10491, new_AGEMA_signal_10490, new_AGEMA_signal_10489, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M54}), .b ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .c ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L5_U1 ( .a ({new_AGEMA_signal_10485, new_AGEMA_signal_10484, new_AGEMA_signal_10483, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M49}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, new_AGEMA_signal_11206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L6_U1 ( .a ({new_AGEMA_signal_11196, new_AGEMA_signal_11195, new_AGEMA_signal_11194, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M62}), .b ({new_AGEMA_signal_11208, new_AGEMA_signal_11207, new_AGEMA_signal_11206, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L5}), .c ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L7_U1 ( .a ({new_AGEMA_signal_10482, new_AGEMA_signal_10481, new_AGEMA_signal_10480, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M46}), .b ({new_AGEMA_signal_11202, new_AGEMA_signal_11201, new_AGEMA_signal_11200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .c ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, new_AGEMA_signal_11794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L8_U1 ( .a ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, new_AGEMA_signal_9778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .b ({new_AGEMA_signal_9789, new_AGEMA_signal_9788, new_AGEMA_signal_9787, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M59}), .c ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L9_U1 ( .a ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, new_AGEMA_signal_10486, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, new_AGEMA_signal_11191, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .c ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L10_U1 ( .a ({new_AGEMA_signal_11193, new_AGEMA_signal_11192, new_AGEMA_signal_11191, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M53}), .b ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, new_AGEMA_signal_11800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L11_U1 ( .a ({new_AGEMA_signal_9792, new_AGEMA_signal_9791, new_AGEMA_signal_9790, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M60}), .b ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, new_AGEMA_signal_11197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L12_U1 ( .a ({new_AGEMA_signal_9774, new_AGEMA_signal_9773, new_AGEMA_signal_9772, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M48}), .b ({new_AGEMA_signal_9780, new_AGEMA_signal_9779, new_AGEMA_signal_9778, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M51}), .c ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, new_AGEMA_signal_10510, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L13_U1 ( .a ({new_AGEMA_signal_9777, new_AGEMA_signal_9776, new_AGEMA_signal_9775, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M50}), .b ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, new_AGEMA_signal_12334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L14_U1 ( .a ({new_AGEMA_signal_10488, new_AGEMA_signal_10487, new_AGEMA_signal_10486, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M52}), .b ({new_AGEMA_signal_10500, new_AGEMA_signal_10499, new_AGEMA_signal_10498, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M61}), .c ({new_AGEMA_signal_11211, new_AGEMA_signal_11210, new_AGEMA_signal_11209, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L15_U1 ( .a ({new_AGEMA_signal_10494, new_AGEMA_signal_10493, new_AGEMA_signal_10492, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M55}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11214, new_AGEMA_signal_11213, new_AGEMA_signal_11212, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L16_U1 ( .a ({new_AGEMA_signal_9783, new_AGEMA_signal_9782, new_AGEMA_signal_9781, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M56}), .b ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .c ({new_AGEMA_signal_12339, new_AGEMA_signal_12338, new_AGEMA_signal_12337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L17_U1 ( .a ({new_AGEMA_signal_9786, new_AGEMA_signal_9785, new_AGEMA_signal_9784, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M57}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_11217, new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L18_U1 ( .a ({new_AGEMA_signal_10497, new_AGEMA_signal_10496, new_AGEMA_signal_10495, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M58}), .b ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .c ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, new_AGEMA_signal_11218, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L19_U1 ( .a ({new_AGEMA_signal_10503, new_AGEMA_signal_10502, new_AGEMA_signal_10501, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_M63}), .b ({new_AGEMA_signal_11205, new_AGEMA_signal_11204, new_AGEMA_signal_11203, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L4}), .c ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, new_AGEMA_signal_11806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L20_U1 ( .a ({new_AGEMA_signal_11790, new_AGEMA_signal_11789, new_AGEMA_signal_11788, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L0}), .b ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .c ({new_AGEMA_signal_12342, new_AGEMA_signal_12341, new_AGEMA_signal_12340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L21_U1 ( .a ({new_AGEMA_signal_10506, new_AGEMA_signal_10505, new_AGEMA_signal_10504, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L1}), .b ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, new_AGEMA_signal_11794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .c ({new_AGEMA_signal_12345, new_AGEMA_signal_12344, new_AGEMA_signal_12343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L22_U1 ( .a ({new_AGEMA_signal_11202, new_AGEMA_signal_11201, new_AGEMA_signal_11200, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L3}), .b ({new_AGEMA_signal_10512, new_AGEMA_signal_10511, new_AGEMA_signal_10510, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L12}), .c ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L23_U1 ( .a ({new_AGEMA_signal_11220, new_AGEMA_signal_11219, new_AGEMA_signal_11218, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L18}), .b ({new_AGEMA_signal_11199, new_AGEMA_signal_11198, new_AGEMA_signal_11197, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L2}), .c ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, new_AGEMA_signal_11812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L24_U1 ( .a ({new_AGEMA_signal_11214, new_AGEMA_signal_11213, new_AGEMA_signal_11212, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L15}), .b ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, new_AGEMA_signal_12346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L25_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, new_AGEMA_signal_11800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12351, new_AGEMA_signal_12350, new_AGEMA_signal_12349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L26_U1 ( .a ({new_AGEMA_signal_11796, new_AGEMA_signal_11795, new_AGEMA_signal_11794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L7}), .b ({new_AGEMA_signal_11799, new_AGEMA_signal_11798, new_AGEMA_signal_11797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L9}), .c ({new_AGEMA_signal_12354, new_AGEMA_signal_12353, new_AGEMA_signal_12352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L27_U1 ( .a ({new_AGEMA_signal_10509, new_AGEMA_signal_10508, new_AGEMA_signal_10507, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L8}), .b ({new_AGEMA_signal_11802, new_AGEMA_signal_11801, new_AGEMA_signal_11800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L10}), .c ({new_AGEMA_signal_12357, new_AGEMA_signal_12356, new_AGEMA_signal_12355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L28_U1 ( .a ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11211, new_AGEMA_signal_11210, new_AGEMA_signal_11209, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L14}), .c ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, new_AGEMA_signal_12358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_L29_U1 ( .a ({new_AGEMA_signal_11805, new_AGEMA_signal_11804, new_AGEMA_signal_11803, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L11}), .b ({new_AGEMA_signal_11217, new_AGEMA_signal_11216, new_AGEMA_signal_11215, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L17}), .c ({new_AGEMA_signal_12363, new_AGEMA_signal_12362, new_AGEMA_signal_12361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S0_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12348, new_AGEMA_signal_12347, new_AGEMA_signal_12346, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L24}), .c ({new_AGEMA_signal_12996, new_AGEMA_signal_12995, new_AGEMA_signal_12994, KeyExpansionIns_tmp[23]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S1_U1 ( .a ({new_AGEMA_signal_12339, new_AGEMA_signal_12338, new_AGEMA_signal_12337, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L16}), .b ({new_AGEMA_signal_12354, new_AGEMA_signal_12353, new_AGEMA_signal_12352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L26}), .c ({new_AGEMA_signal_12999, new_AGEMA_signal_12998, new_AGEMA_signal_12997, KeyExpansionIns_tmp[22]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S2_U1 ( .a ({new_AGEMA_signal_11808, new_AGEMA_signal_11807, new_AGEMA_signal_11806, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L19}), .b ({new_AGEMA_signal_12360, new_AGEMA_signal_12359, new_AGEMA_signal_12358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L28}), .c ({new_AGEMA_signal_13002, new_AGEMA_signal_13001, new_AGEMA_signal_13000, KeyExpansionIns_tmp[21]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S3_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_12345, new_AGEMA_signal_12344, new_AGEMA_signal_12343, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L21}), .c ({new_AGEMA_signal_13005, new_AGEMA_signal_13004, new_AGEMA_signal_13003, KeyExpansionIns_tmp[20]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S4_U1 ( .a ({new_AGEMA_signal_12342, new_AGEMA_signal_12341, new_AGEMA_signal_12340, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L20}), .b ({new_AGEMA_signal_11811, new_AGEMA_signal_11810, new_AGEMA_signal_11809, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L22}), .c ({new_AGEMA_signal_13008, new_AGEMA_signal_13007, new_AGEMA_signal_13006, KeyExpansionIns_tmp[19]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S5_U1 ( .a ({new_AGEMA_signal_12351, new_AGEMA_signal_12350, new_AGEMA_signal_12349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L25}), .b ({new_AGEMA_signal_12363, new_AGEMA_signal_12362, new_AGEMA_signal_12361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L29}), .c ({new_AGEMA_signal_13011, new_AGEMA_signal_13010, new_AGEMA_signal_13009, KeyExpansionIns_tmp[18]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S6_U1 ( .a ({new_AGEMA_signal_12336, new_AGEMA_signal_12335, new_AGEMA_signal_12334, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L13}), .b ({new_AGEMA_signal_12357, new_AGEMA_signal_12356, new_AGEMA_signal_12355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L27}), .c ({new_AGEMA_signal_13014, new_AGEMA_signal_13013, new_AGEMA_signal_13012, KeyExpansionIns_tmp[17]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_XOR_S7_U1 ( .a ({new_AGEMA_signal_11793, new_AGEMA_signal_11792, new_AGEMA_signal_11791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L6}), .b ({new_AGEMA_signal_11814, new_AGEMA_signal_11813, new_AGEMA_signal_11812, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_1_L23}), .c ({new_AGEMA_signal_12366, new_AGEMA_signal_12365, new_AGEMA_signal_12364, KeyExpansionIns_tmp[16]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M46_U1 ( .a ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, new_AGEMA_signal_9802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_6351, new_AGEMA_signal_6350, new_AGEMA_signal_6349, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T6}), .clk (clk), .r ({Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864]}), .c ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, new_AGEMA_signal_10516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M47_U1 ( .a ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_6861, new_AGEMA_signal_6860, new_AGEMA_signal_6859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T8}), .clk (clk), .r ({Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870]}), .c ({new_AGEMA_signal_9807, new_AGEMA_signal_9806, new_AGEMA_signal_9805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M48_U1 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}), .clk (clk), .r ({Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876]}), .c ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, new_AGEMA_signal_9808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M49_U1 ( .a ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_6363, new_AGEMA_signal_6362, new_AGEMA_signal_6361, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T16}), .clk (clk), .r ({Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882]}), .c ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M50_U1 ( .a ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6354, new_AGEMA_signal_6353, new_AGEMA_signal_6352, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T9}), .clk (clk), .r ({Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888]}), .c ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, new_AGEMA_signal_9811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M51_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6870, new_AGEMA_signal_6869, new_AGEMA_signal_6868, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T17}), .clk (clk), .r ({Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894]}), .c ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, new_AGEMA_signal_9814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M52_U1 ( .a ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_6360, new_AGEMA_signal_6359, new_AGEMA_signal_6358, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T15}), .clk (clk), .r ({Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900]}), .c ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, new_AGEMA_signal_10522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M53_U1 ( .a ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_6372, new_AGEMA_signal_6371, new_AGEMA_signal_6370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T27}), .clk (clk), .r ({Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906]}), .c ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, new_AGEMA_signal_11221, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M54_U1 ( .a ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_6864, new_AGEMA_signal_6863, new_AGEMA_signal_6862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T10}), .clk (clk), .r ({Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912]}), .c ({new_AGEMA_signal_10527, new_AGEMA_signal_10526, new_AGEMA_signal_10525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M55_U1 ( .a ({new_AGEMA_signal_9804, new_AGEMA_signal_9803, new_AGEMA_signal_9802, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M44}), .b ({new_AGEMA_signal_6357, new_AGEMA_signal_6356, new_AGEMA_signal_6355, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T13}), .clk (clk), .r ({Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918]}), .c ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, new_AGEMA_signal_10528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M56_U1 ( .a ({new_AGEMA_signal_9516, new_AGEMA_signal_9515, new_AGEMA_signal_9514, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M40}), .b ({new_AGEMA_signal_6876, new_AGEMA_signal_6875, new_AGEMA_signal_6874, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T23}), .clk (clk), .r ({Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924]}), .c ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, new_AGEMA_signal_9817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M57_U1 ( .a ({new_AGEMA_signal_9513, new_AGEMA_signal_9512, new_AGEMA_signal_9511, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M39}), .b ({new_AGEMA_signal_6366, new_AGEMA_signal_6365, new_AGEMA_signal_6364, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T19}), .clk (clk), .r ({Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930]}), .c ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, new_AGEMA_signal_9820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M58_U1 ( .a ({new_AGEMA_signal_9801, new_AGEMA_signal_9800, new_AGEMA_signal_9799, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M43}), .b ({new_AGEMA_signal_5769, new_AGEMA_signal_5768, new_AGEMA_signal_5767, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T3}), .clk (clk), .r ({Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936]}), .c ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, new_AGEMA_signal_10531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M59_U1 ( .a ({new_AGEMA_signal_9510, new_AGEMA_signal_9509, new_AGEMA_signal_9508, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M38}), .b ({new_AGEMA_signal_6369, new_AGEMA_signal_6368, new_AGEMA_signal_6367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T22}), .clk (clk), .r ({Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942]}), .c ({new_AGEMA_signal_9825, new_AGEMA_signal_9824, new_AGEMA_signal_9823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M60_U1 ( .a ({new_AGEMA_signal_9507, new_AGEMA_signal_9506, new_AGEMA_signal_9505, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M37}), .b ({new_AGEMA_signal_6873, new_AGEMA_signal_6872, new_AGEMA_signal_6871, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T20}), .clk (clk), .r ({Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948]}), .c ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, new_AGEMA_signal_9826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M61_U1 ( .a ({new_AGEMA_signal_9798, new_AGEMA_signal_9797, new_AGEMA_signal_9796, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M42}), .b ({new_AGEMA_signal_5763, new_AGEMA_signal_5762, new_AGEMA_signal_5761, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T1}), .clk (clk), .r ({Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954]}), .c ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M62_U1 ( .a ({new_AGEMA_signal_10515, new_AGEMA_signal_10514, new_AGEMA_signal_10513, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M45}), .b ({new_AGEMA_signal_5772, new_AGEMA_signal_5771, new_AGEMA_signal_5770, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T4}), .clk (clk), .r ({Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960]}), .c ({new_AGEMA_signal_11226, new_AGEMA_signal_11225, new_AGEMA_signal_11224, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_AND_M63_U1 ( .a ({new_AGEMA_signal_9795, new_AGEMA_signal_9794, new_AGEMA_signal_9793, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M41}), .b ({new_AGEMA_signal_5766, new_AGEMA_signal_5765, new_AGEMA_signal_5764, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_T2}), .clk (clk), .r ({Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966]}), .c ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, new_AGEMA_signal_10537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L0_U1 ( .a ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .b ({new_AGEMA_signal_11226, new_AGEMA_signal_11225, new_AGEMA_signal_11224, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .c ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L1_U1 ( .a ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, new_AGEMA_signal_9811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, new_AGEMA_signal_9817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .c ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L2_U1 ( .a ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, new_AGEMA_signal_10516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, new_AGEMA_signal_9808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .c ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L3_U1 ( .a ({new_AGEMA_signal_9807, new_AGEMA_signal_9806, new_AGEMA_signal_9805, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M47}), .b ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, new_AGEMA_signal_10528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .c ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, new_AGEMA_signal_11230, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L4_U1 ( .a ({new_AGEMA_signal_10527, new_AGEMA_signal_10526, new_AGEMA_signal_10525, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M54}), .b ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, new_AGEMA_signal_10531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .c ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, new_AGEMA_signal_11233, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L5_U1 ( .a ({new_AGEMA_signal_10521, new_AGEMA_signal_10520, new_AGEMA_signal_10519, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M49}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11238, new_AGEMA_signal_11237, new_AGEMA_signal_11236, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L6_U1 ( .a ({new_AGEMA_signal_11226, new_AGEMA_signal_11225, new_AGEMA_signal_11224, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M62}), .b ({new_AGEMA_signal_11238, new_AGEMA_signal_11237, new_AGEMA_signal_11236, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L5}), .c ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L7_U1 ( .a ({new_AGEMA_signal_10518, new_AGEMA_signal_10517, new_AGEMA_signal_10516, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M46}), .b ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, new_AGEMA_signal_11230, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .c ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L8_U1 ( .a ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, new_AGEMA_signal_9814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .b ({new_AGEMA_signal_9825, new_AGEMA_signal_9824, new_AGEMA_signal_9823, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M59}), .c ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, new_AGEMA_signal_10543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L9_U1 ( .a ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, new_AGEMA_signal_10522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, new_AGEMA_signal_11221, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .c ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, new_AGEMA_signal_11824, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L10_U1 ( .a ({new_AGEMA_signal_11223, new_AGEMA_signal_11222, new_AGEMA_signal_11221, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M53}), .b ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, new_AGEMA_signal_11233, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L11_U1 ( .a ({new_AGEMA_signal_9828, new_AGEMA_signal_9827, new_AGEMA_signal_9826, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M60}), .b ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, new_AGEMA_signal_11830, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L12_U1 ( .a ({new_AGEMA_signal_9810, new_AGEMA_signal_9809, new_AGEMA_signal_9808, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M48}), .b ({new_AGEMA_signal_9816, new_AGEMA_signal_9815, new_AGEMA_signal_9814, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M51}), .c ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, new_AGEMA_signal_10546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L13_U1 ( .a ({new_AGEMA_signal_9813, new_AGEMA_signal_9812, new_AGEMA_signal_9811, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M50}), .b ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, new_AGEMA_signal_12367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L14_U1 ( .a ({new_AGEMA_signal_10524, new_AGEMA_signal_10523, new_AGEMA_signal_10522, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M52}), .b ({new_AGEMA_signal_10536, new_AGEMA_signal_10535, new_AGEMA_signal_10534, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M61}), .c ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L15_U1 ( .a ({new_AGEMA_signal_10530, new_AGEMA_signal_10529, new_AGEMA_signal_10528, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M55}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, new_AGEMA_signal_11242, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L16_U1 ( .a ({new_AGEMA_signal_9819, new_AGEMA_signal_9818, new_AGEMA_signal_9817, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M56}), .b ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .c ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, new_AGEMA_signal_12370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L17_U1 ( .a ({new_AGEMA_signal_9822, new_AGEMA_signal_9821, new_AGEMA_signal_9820, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M57}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_11247, new_AGEMA_signal_11246, new_AGEMA_signal_11245, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L18_U1 ( .a ({new_AGEMA_signal_10533, new_AGEMA_signal_10532, new_AGEMA_signal_10531, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M58}), .b ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, new_AGEMA_signal_10543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .c ({new_AGEMA_signal_11250, new_AGEMA_signal_11249, new_AGEMA_signal_11248, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L19_U1 ( .a ({new_AGEMA_signal_10539, new_AGEMA_signal_10538, new_AGEMA_signal_10537, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_M63}), .b ({new_AGEMA_signal_11235, new_AGEMA_signal_11234, new_AGEMA_signal_11233, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L4}), .c ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, new_AGEMA_signal_11833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L20_U1 ( .a ({new_AGEMA_signal_11817, new_AGEMA_signal_11816, new_AGEMA_signal_11815, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L0}), .b ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .c ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, new_AGEMA_signal_12373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L21_U1 ( .a ({new_AGEMA_signal_10542, new_AGEMA_signal_10541, new_AGEMA_signal_10540, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L1}), .b ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .c ({new_AGEMA_signal_12378, new_AGEMA_signal_12377, new_AGEMA_signal_12376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L22_U1 ( .a ({new_AGEMA_signal_11232, new_AGEMA_signal_11231, new_AGEMA_signal_11230, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L3}), .b ({new_AGEMA_signal_10548, new_AGEMA_signal_10547, new_AGEMA_signal_10546, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L12}), .c ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, new_AGEMA_signal_11836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L23_U1 ( .a ({new_AGEMA_signal_11250, new_AGEMA_signal_11249, new_AGEMA_signal_11248, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L18}), .b ({new_AGEMA_signal_11229, new_AGEMA_signal_11228, new_AGEMA_signal_11227, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L2}), .c ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, new_AGEMA_signal_11839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L24_U1 ( .a ({new_AGEMA_signal_11244, new_AGEMA_signal_11243, new_AGEMA_signal_11242, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L15}), .b ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, new_AGEMA_signal_11824, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, new_AGEMA_signal_12379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L25_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, new_AGEMA_signal_12382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L26_U1 ( .a ({new_AGEMA_signal_11823, new_AGEMA_signal_11822, new_AGEMA_signal_11821, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L7}), .b ({new_AGEMA_signal_11826, new_AGEMA_signal_11825, new_AGEMA_signal_11824, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L9}), .c ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, new_AGEMA_signal_12385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L27_U1 ( .a ({new_AGEMA_signal_10545, new_AGEMA_signal_10544, new_AGEMA_signal_10543, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L8}), .b ({new_AGEMA_signal_11829, new_AGEMA_signal_11828, new_AGEMA_signal_11827, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L10}), .c ({new_AGEMA_signal_12390, new_AGEMA_signal_12389, new_AGEMA_signal_12388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L28_U1 ( .a ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, new_AGEMA_signal_11830, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11241, new_AGEMA_signal_11240, new_AGEMA_signal_11239, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L14}), .c ({new_AGEMA_signal_12393, new_AGEMA_signal_12392, new_AGEMA_signal_12391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_L29_U1 ( .a ({new_AGEMA_signal_11832, new_AGEMA_signal_11831, new_AGEMA_signal_11830, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L11}), .b ({new_AGEMA_signal_11247, new_AGEMA_signal_11246, new_AGEMA_signal_11245, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L17}), .c ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, new_AGEMA_signal_12394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S0_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12381, new_AGEMA_signal_12380, new_AGEMA_signal_12379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L24}), .c ({new_AGEMA_signal_13017, new_AGEMA_signal_13016, new_AGEMA_signal_13015, KeyExpansionIns_tmp[15]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S1_U1 ( .a ({new_AGEMA_signal_12372, new_AGEMA_signal_12371, new_AGEMA_signal_12370, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L16}), .b ({new_AGEMA_signal_12387, new_AGEMA_signal_12386, new_AGEMA_signal_12385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L26}), .c ({new_AGEMA_signal_13020, new_AGEMA_signal_13019, new_AGEMA_signal_13018, KeyExpansionIns_tmp[14]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S2_U1 ( .a ({new_AGEMA_signal_11835, new_AGEMA_signal_11834, new_AGEMA_signal_11833, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L19}), .b ({new_AGEMA_signal_12393, new_AGEMA_signal_12392, new_AGEMA_signal_12391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L28}), .c ({new_AGEMA_signal_13023, new_AGEMA_signal_13022, new_AGEMA_signal_13021, KeyExpansionIns_tmp[13]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S3_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_12378, new_AGEMA_signal_12377, new_AGEMA_signal_12376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L21}), .c ({new_AGEMA_signal_13026, new_AGEMA_signal_13025, new_AGEMA_signal_13024, KeyExpansionIns_tmp[12]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S4_U1 ( .a ({new_AGEMA_signal_12375, new_AGEMA_signal_12374, new_AGEMA_signal_12373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L20}), .b ({new_AGEMA_signal_11838, new_AGEMA_signal_11837, new_AGEMA_signal_11836, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L22}), .c ({new_AGEMA_signal_13029, new_AGEMA_signal_13028, new_AGEMA_signal_13027, KeyExpansionIns_tmp[11]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S5_U1 ( .a ({new_AGEMA_signal_12384, new_AGEMA_signal_12383, new_AGEMA_signal_12382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L25}), .b ({new_AGEMA_signal_12396, new_AGEMA_signal_12395, new_AGEMA_signal_12394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L29}), .c ({new_AGEMA_signal_13032, new_AGEMA_signal_13031, new_AGEMA_signal_13030, KeyExpansionIns_tmp[10]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S6_U1 ( .a ({new_AGEMA_signal_12369, new_AGEMA_signal_12368, new_AGEMA_signal_12367, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L13}), .b ({new_AGEMA_signal_12390, new_AGEMA_signal_12389, new_AGEMA_signal_12388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L27}), .c ({new_AGEMA_signal_13035, new_AGEMA_signal_13034, new_AGEMA_signal_13033, KeyExpansionIns_tmp[9]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_XOR_S7_U1 ( .a ({new_AGEMA_signal_11820, new_AGEMA_signal_11819, new_AGEMA_signal_11818, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L6}), .b ({new_AGEMA_signal_11841, new_AGEMA_signal_11840, new_AGEMA_signal_11839, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_2_L23}), .c ({new_AGEMA_signal_12399, new_AGEMA_signal_12398, new_AGEMA_signal_12397, KeyExpansionIns_tmp[8]}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M46_U1 ( .a ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, new_AGEMA_signal_9838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_6375, new_AGEMA_signal_6374, new_AGEMA_signal_6373, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T6}), .clk (clk), .r ({Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972]}), .c ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, new_AGEMA_signal_10552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M47_U1 ( .a ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_6900, new_AGEMA_signal_6899, new_AGEMA_signal_6898, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T8}), .clk (clk), .r ({Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978]}), .c ({new_AGEMA_signal_9843, new_AGEMA_signal_9842, new_AGEMA_signal_9841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M48_U1 ( .a ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}), .clk (clk), .r ({Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984]}), .c ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, new_AGEMA_signal_9844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M49_U1 ( .a ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, new_AGEMA_signal_9835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_6387, new_AGEMA_signal_6386, new_AGEMA_signal_6385, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T16}), .clk (clk), .r ({Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990]}), .c ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, new_AGEMA_signal_10555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M50_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6378, new_AGEMA_signal_6377, new_AGEMA_signal_6376, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T9}), .clk (clk), .r ({Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996]}), .c ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, new_AGEMA_signal_9847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M51_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6909, new_AGEMA_signal_6908, new_AGEMA_signal_6907, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T17}), .clk (clk), .r ({Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002]}), .c ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, new_AGEMA_signal_9850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M52_U1 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_6384, new_AGEMA_signal_6383, new_AGEMA_signal_6382, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T15}), .clk (clk), .r ({Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008]}), .c ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, new_AGEMA_signal_10558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M53_U1 ( .a ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, new_AGEMA_signal_10549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_6396, new_AGEMA_signal_6395, new_AGEMA_signal_6394, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T27}), .clk (clk), .r ({Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014]}), .c ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M54_U1 ( .a ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_6903, new_AGEMA_signal_6902, new_AGEMA_signal_6901, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T10}), .clk (clk), .r ({Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020]}), .c ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, new_AGEMA_signal_10561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M55_U1 ( .a ({new_AGEMA_signal_9840, new_AGEMA_signal_9839, new_AGEMA_signal_9838, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M44}), .b ({new_AGEMA_signal_6381, new_AGEMA_signal_6380, new_AGEMA_signal_6379, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T13}), .clk (clk), .r ({Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026]}), .c ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, new_AGEMA_signal_10564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M56_U1 ( .a ({new_AGEMA_signal_9528, new_AGEMA_signal_9527, new_AGEMA_signal_9526, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M40}), .b ({new_AGEMA_signal_6915, new_AGEMA_signal_6914, new_AGEMA_signal_6913, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T23}), .clk (clk), .r ({Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032]}), .c ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, new_AGEMA_signal_9853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M57_U1 ( .a ({new_AGEMA_signal_9525, new_AGEMA_signal_9524, new_AGEMA_signal_9523, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M39}), .b ({new_AGEMA_signal_6390, new_AGEMA_signal_6389, new_AGEMA_signal_6388, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T19}), .clk (clk), .r ({Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038]}), .c ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, new_AGEMA_signal_9856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M58_U1 ( .a ({new_AGEMA_signal_9837, new_AGEMA_signal_9836, new_AGEMA_signal_9835, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M43}), .b ({new_AGEMA_signal_5799, new_AGEMA_signal_5798, new_AGEMA_signal_5797, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T3}), .clk (clk), .r ({Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044]}), .c ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, new_AGEMA_signal_10567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M59_U1 ( .a ({new_AGEMA_signal_9522, new_AGEMA_signal_9521, new_AGEMA_signal_9520, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M38}), .b ({new_AGEMA_signal_6393, new_AGEMA_signal_6392, new_AGEMA_signal_6391, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T22}), .clk (clk), .r ({Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050]}), .c ({new_AGEMA_signal_9861, new_AGEMA_signal_9860, new_AGEMA_signal_9859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M60_U1 ( .a ({new_AGEMA_signal_9519, new_AGEMA_signal_9518, new_AGEMA_signal_9517, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M37}), .b ({new_AGEMA_signal_6912, new_AGEMA_signal_6911, new_AGEMA_signal_6910, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T20}), .clk (clk), .r ({Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056]}), .c ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, new_AGEMA_signal_9862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M61_U1 ( .a ({new_AGEMA_signal_9834, new_AGEMA_signal_9833, new_AGEMA_signal_9832, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M42}), .b ({new_AGEMA_signal_5793, new_AGEMA_signal_5792, new_AGEMA_signal_5791, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T1}), .clk (clk), .r ({Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062]}), .c ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M62_U1 ( .a ({new_AGEMA_signal_10551, new_AGEMA_signal_10550, new_AGEMA_signal_10549, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M45}), .b ({new_AGEMA_signal_5802, new_AGEMA_signal_5801, new_AGEMA_signal_5800, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T4}), .clk (clk), .r ({Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068]}), .c ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, new_AGEMA_signal_11254, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}) ) ;
    and_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_AND_M63_U1 ( .a ({new_AGEMA_signal_9831, new_AGEMA_signal_9830, new_AGEMA_signal_9829, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M41}), .b ({new_AGEMA_signal_5796, new_AGEMA_signal_5795, new_AGEMA_signal_5794, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_T2}), .clk (clk), .r ({Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074]}), .c ({new_AGEMA_signal_10575, new_AGEMA_signal_10574, new_AGEMA_signal_10573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L0_U1 ( .a ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .b ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, new_AGEMA_signal_11254, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .c ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L1_U1 ( .a ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, new_AGEMA_signal_9847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, new_AGEMA_signal_9853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .c ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L2_U1 ( .a ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, new_AGEMA_signal_10552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, new_AGEMA_signal_9844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .c ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, new_AGEMA_signal_11257, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L3_U1 ( .a ({new_AGEMA_signal_9843, new_AGEMA_signal_9842, new_AGEMA_signal_9841, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M47}), .b ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, new_AGEMA_signal_10564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .c ({new_AGEMA_signal_11262, new_AGEMA_signal_11261, new_AGEMA_signal_11260, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L4_U1 ( .a ({new_AGEMA_signal_10563, new_AGEMA_signal_10562, new_AGEMA_signal_10561, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M54}), .b ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, new_AGEMA_signal_10567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .c ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L5_U1 ( .a ({new_AGEMA_signal_10557, new_AGEMA_signal_10556, new_AGEMA_signal_10555, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M49}), .b ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, new_AGEMA_signal_11266, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L6_U1 ( .a ({new_AGEMA_signal_11256, new_AGEMA_signal_11255, new_AGEMA_signal_11254, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M62}), .b ({new_AGEMA_signal_11268, new_AGEMA_signal_11267, new_AGEMA_signal_11266, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L5}), .c ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L7_U1 ( .a ({new_AGEMA_signal_10554, new_AGEMA_signal_10553, new_AGEMA_signal_10552, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M46}), .b ({new_AGEMA_signal_11262, new_AGEMA_signal_11261, new_AGEMA_signal_11260, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .c ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, new_AGEMA_signal_11848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L8_U1 ( .a ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, new_AGEMA_signal_9850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .b ({new_AGEMA_signal_9861, new_AGEMA_signal_9860, new_AGEMA_signal_9859, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M59}), .c ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, new_AGEMA_signal_10579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L9_U1 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, new_AGEMA_signal_10558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .c ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, new_AGEMA_signal_11851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L10_U1 ( .a ({new_AGEMA_signal_11253, new_AGEMA_signal_11252, new_AGEMA_signal_11251, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M53}), .b ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, new_AGEMA_signal_11854, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L11_U1 ( .a ({new_AGEMA_signal_9864, new_AGEMA_signal_9863, new_AGEMA_signal_9862, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M60}), .b ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, new_AGEMA_signal_11257, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, new_AGEMA_signal_11857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L12_U1 ( .a ({new_AGEMA_signal_9846, new_AGEMA_signal_9845, new_AGEMA_signal_9844, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M48}), .b ({new_AGEMA_signal_9852, new_AGEMA_signal_9851, new_AGEMA_signal_9850, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M51}), .c ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, new_AGEMA_signal_10582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L13_U1 ( .a ({new_AGEMA_signal_9849, new_AGEMA_signal_9848, new_AGEMA_signal_9847, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M50}), .b ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12402, new_AGEMA_signal_12401, new_AGEMA_signal_12400, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L14_U1 ( .a ({new_AGEMA_signal_10560, new_AGEMA_signal_10559, new_AGEMA_signal_10558, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M52}), .b ({new_AGEMA_signal_10572, new_AGEMA_signal_10571, new_AGEMA_signal_10570, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M61}), .c ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, new_AGEMA_signal_11269, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L15_U1 ( .a ({new_AGEMA_signal_10566, new_AGEMA_signal_10565, new_AGEMA_signal_10564, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M55}), .b ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11274, new_AGEMA_signal_11273, new_AGEMA_signal_11272, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L16_U1 ( .a ({new_AGEMA_signal_9855, new_AGEMA_signal_9854, new_AGEMA_signal_9853, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M56}), .b ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .c ({new_AGEMA_signal_12405, new_AGEMA_signal_12404, new_AGEMA_signal_12403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L17_U1 ( .a ({new_AGEMA_signal_9858, new_AGEMA_signal_9857, new_AGEMA_signal_9856, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M57}), .b ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L18_U1 ( .a ({new_AGEMA_signal_10569, new_AGEMA_signal_10568, new_AGEMA_signal_10567, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M58}), .b ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, new_AGEMA_signal_10579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .c ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, new_AGEMA_signal_11278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L19_U1 ( .a ({new_AGEMA_signal_10575, new_AGEMA_signal_10574, new_AGEMA_signal_10573, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_M63}), .b ({new_AGEMA_signal_11265, new_AGEMA_signal_11264, new_AGEMA_signal_11263, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L4}), .c ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, new_AGEMA_signal_11860, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L20_U1 ( .a ({new_AGEMA_signal_11844, new_AGEMA_signal_11843, new_AGEMA_signal_11842, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L0}), .b ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .c ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, new_AGEMA_signal_12406, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L21_U1 ( .a ({new_AGEMA_signal_10578, new_AGEMA_signal_10577, new_AGEMA_signal_10576, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L1}), .b ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, new_AGEMA_signal_11848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .c ({new_AGEMA_signal_12411, new_AGEMA_signal_12410, new_AGEMA_signal_12409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L22_U1 ( .a ({new_AGEMA_signal_11262, new_AGEMA_signal_11261, new_AGEMA_signal_11260, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L3}), .b ({new_AGEMA_signal_10584, new_AGEMA_signal_10583, new_AGEMA_signal_10582, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L12}), .c ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, new_AGEMA_signal_11863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L23_U1 ( .a ({new_AGEMA_signal_11280, new_AGEMA_signal_11279, new_AGEMA_signal_11278, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L18}), .b ({new_AGEMA_signal_11259, new_AGEMA_signal_11258, new_AGEMA_signal_11257, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L2}), .c ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, new_AGEMA_signal_11866, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L24_U1 ( .a ({new_AGEMA_signal_11274, new_AGEMA_signal_11273, new_AGEMA_signal_11272, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L15}), .b ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, new_AGEMA_signal_11851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12414, new_AGEMA_signal_12413, new_AGEMA_signal_12412, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L25_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, new_AGEMA_signal_11854, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, new_AGEMA_signal_12415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L26_U1 ( .a ({new_AGEMA_signal_11850, new_AGEMA_signal_11849, new_AGEMA_signal_11848, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L7}), .b ({new_AGEMA_signal_11853, new_AGEMA_signal_11852, new_AGEMA_signal_11851, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L9}), .c ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, new_AGEMA_signal_12418, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L27_U1 ( .a ({new_AGEMA_signal_10581, new_AGEMA_signal_10580, new_AGEMA_signal_10579, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L8}), .b ({new_AGEMA_signal_11856, new_AGEMA_signal_11855, new_AGEMA_signal_11854, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L10}), .c ({new_AGEMA_signal_12423, new_AGEMA_signal_12422, new_AGEMA_signal_12421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L28_U1 ( .a ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, new_AGEMA_signal_11857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11271, new_AGEMA_signal_11270, new_AGEMA_signal_11269, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L14}), .c ({new_AGEMA_signal_12426, new_AGEMA_signal_12425, new_AGEMA_signal_12424, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_L29_U1 ( .a ({new_AGEMA_signal_11859, new_AGEMA_signal_11858, new_AGEMA_signal_11857, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L11}), .b ({new_AGEMA_signal_11277, new_AGEMA_signal_11276, new_AGEMA_signal_11275, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L17}), .c ({new_AGEMA_signal_12429, new_AGEMA_signal_12428, new_AGEMA_signal_12427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S0_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12414, new_AGEMA_signal_12413, new_AGEMA_signal_12412, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L24}), .c ({new_AGEMA_signal_13038, new_AGEMA_signal_13037, new_AGEMA_signal_13036, KeyExpansionIns_tmp[7]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S1_U1 ( .a ({new_AGEMA_signal_12405, new_AGEMA_signal_12404, new_AGEMA_signal_12403, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L16}), .b ({new_AGEMA_signal_12420, new_AGEMA_signal_12419, new_AGEMA_signal_12418, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L26}), .c ({new_AGEMA_signal_13041, new_AGEMA_signal_13040, new_AGEMA_signal_13039, KeyExpansionIns_tmp[6]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S2_U1 ( .a ({new_AGEMA_signal_11862, new_AGEMA_signal_11861, new_AGEMA_signal_11860, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L19}), .b ({new_AGEMA_signal_12426, new_AGEMA_signal_12425, new_AGEMA_signal_12424, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L28}), .c ({new_AGEMA_signal_13044, new_AGEMA_signal_13043, new_AGEMA_signal_13042, KeyExpansionIns_tmp[5]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S3_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_12411, new_AGEMA_signal_12410, new_AGEMA_signal_12409, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L21}), .c ({new_AGEMA_signal_13047, new_AGEMA_signal_13046, new_AGEMA_signal_13045, KeyExpansionIns_tmp[4]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S4_U1 ( .a ({new_AGEMA_signal_12408, new_AGEMA_signal_12407, new_AGEMA_signal_12406, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L20}), .b ({new_AGEMA_signal_11865, new_AGEMA_signal_11864, new_AGEMA_signal_11863, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L22}), .c ({new_AGEMA_signal_13050, new_AGEMA_signal_13049, new_AGEMA_signal_13048, KeyExpansionIns_tmp[3]}) ) ;
    xor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S5_U1 ( .a ({new_AGEMA_signal_12417, new_AGEMA_signal_12416, new_AGEMA_signal_12415, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L25}), .b ({new_AGEMA_signal_12429, new_AGEMA_signal_12428, new_AGEMA_signal_12427, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L29}), .c ({new_AGEMA_signal_13053, new_AGEMA_signal_13052, new_AGEMA_signal_13051, KeyExpansionIns_tmp[2]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S6_U1 ( .a ({new_AGEMA_signal_12402, new_AGEMA_signal_12401, new_AGEMA_signal_12400, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L13}), .b ({new_AGEMA_signal_12423, new_AGEMA_signal_12422, new_AGEMA_signal_12421, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L27}), .c ({new_AGEMA_signal_13056, new_AGEMA_signal_13055, new_AGEMA_signal_13054, KeyExpansionIns_tmp[1]}) ) ;
    xnor_HPC2 #(.security_order(3), .pipeline(0)) KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_XOR_S7_U1 ( .a ({new_AGEMA_signal_11847, new_AGEMA_signal_11846, new_AGEMA_signal_11845, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L6}), .b ({new_AGEMA_signal_11868, new_AGEMA_signal_11867, new_AGEMA_signal_11866, KeyExpansionIns_KeySchedCoreInst_Inst_Sbox_3_L23}), .c ({new_AGEMA_signal_12432, new_AGEMA_signal_12431, new_AGEMA_signal_12430, KeyExpansionIns_tmp[0]}) ) ;

    /* register cells */
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16200, new_AGEMA_signal_16199, new_AGEMA_signal_16198, RoundReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, new_AGEMA_signal_4549, RoundInput[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16722, new_AGEMA_signal_16721, new_AGEMA_signal_16720, RoundReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4902, new_AGEMA_signal_4901, new_AGEMA_signal_4900, RoundInput[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16206, new_AGEMA_signal_16205, new_AGEMA_signal_16204, RoundReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, new_AGEMA_signal_4999, RoundInput[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16728, new_AGEMA_signal_16727, new_AGEMA_signal_16726, RoundReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_5100, new_AGEMA_signal_5099, new_AGEMA_signal_5098, RoundInput[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16734, new_AGEMA_signal_16733, new_AGEMA_signal_16732, RoundReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_5199, new_AGEMA_signal_5198, new_AGEMA_signal_5197, RoundInput[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16212, new_AGEMA_signal_16211, new_AGEMA_signal_16210, RoundReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5298, new_AGEMA_signal_5297, new_AGEMA_signal_5296, RoundInput[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16218, new_AGEMA_signal_16217, new_AGEMA_signal_16216, RoundReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5397, new_AGEMA_signal_5396, new_AGEMA_signal_5395, RoundInput[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16224, new_AGEMA_signal_16223, new_AGEMA_signal_16222, RoundReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5496, new_AGEMA_signal_5495, new_AGEMA_signal_5494, RoundInput[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16230, new_AGEMA_signal_16229, new_AGEMA_signal_16228, RoundReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5595, new_AGEMA_signal_5594, new_AGEMA_signal_5593, RoundInput[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16740, new_AGEMA_signal_16739, new_AGEMA_signal_16738, RoundReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5694, new_AGEMA_signal_5693, new_AGEMA_signal_5692, RoundInput[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16236, new_AGEMA_signal_16235, new_AGEMA_signal_16234, RoundReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4650, new_AGEMA_signal_4649, new_AGEMA_signal_4648, RoundInput[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16746, new_AGEMA_signal_16745, new_AGEMA_signal_16744, RoundReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, new_AGEMA_signal_4747, RoundInput[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16752, new_AGEMA_signal_16751, new_AGEMA_signal_16750, RoundReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4830, new_AGEMA_signal_4829, new_AGEMA_signal_4828, RoundInput[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16242, new_AGEMA_signal_16241, new_AGEMA_signal_16240, RoundReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, new_AGEMA_signal_4837, RoundInput[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16248, new_AGEMA_signal_16247, new_AGEMA_signal_16246, RoundReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4848, new_AGEMA_signal_4847, new_AGEMA_signal_4846, RoundInput[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16254, new_AGEMA_signal_16253, new_AGEMA_signal_16252, RoundReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, new_AGEMA_signal_4855, RoundInput[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16260, new_AGEMA_signal_16259, new_AGEMA_signal_16258, RoundReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4866, new_AGEMA_signal_4865, new_AGEMA_signal_4864, RoundInput[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16758, new_AGEMA_signal_16757, new_AGEMA_signal_16756, RoundReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, new_AGEMA_signal_4873, RoundInput[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16266, new_AGEMA_signal_16265, new_AGEMA_signal_16264, RoundReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4884, new_AGEMA_signal_4883, new_AGEMA_signal_4882, RoundInput[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16764, new_AGEMA_signal_16763, new_AGEMA_signal_16762, RoundReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, new_AGEMA_signal_4891, RoundInput[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16770, new_AGEMA_signal_16769, new_AGEMA_signal_16768, RoundReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, new_AGEMA_signal_4909, RoundInput[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16272, new_AGEMA_signal_16271, new_AGEMA_signal_16270, RoundReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4920, new_AGEMA_signal_4919, new_AGEMA_signal_4918, RoundInput[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16278, new_AGEMA_signal_16277, new_AGEMA_signal_16276, RoundReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, new_AGEMA_signal_4927, RoundInput[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16284, new_AGEMA_signal_16283, new_AGEMA_signal_16282, RoundReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4938, new_AGEMA_signal_4937, new_AGEMA_signal_4936, RoundInput[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16290, new_AGEMA_signal_16289, new_AGEMA_signal_16288, RoundReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, new_AGEMA_signal_4945, RoundInput[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16776, new_AGEMA_signal_16775, new_AGEMA_signal_16774, RoundReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4956, new_AGEMA_signal_4955, new_AGEMA_signal_4954, RoundInput[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16296, new_AGEMA_signal_16295, new_AGEMA_signal_16294, RoundReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, new_AGEMA_signal_4963, RoundInput[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16782, new_AGEMA_signal_16781, new_AGEMA_signal_16780, RoundReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4974, new_AGEMA_signal_4973, new_AGEMA_signal_4972, RoundInput[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16788, new_AGEMA_signal_16787, new_AGEMA_signal_16786, RoundReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, new_AGEMA_signal_4981, RoundInput[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16302, new_AGEMA_signal_16301, new_AGEMA_signal_16300, RoundReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4992, new_AGEMA_signal_4991, new_AGEMA_signal_4990, RoundInput[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16308, new_AGEMA_signal_16307, new_AGEMA_signal_16306, RoundReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_5010, new_AGEMA_signal_5009, new_AGEMA_signal_5008, RoundInput[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16314, new_AGEMA_signal_16313, new_AGEMA_signal_16312, RoundReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, new_AGEMA_signal_5017, RoundInput[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16320, new_AGEMA_signal_16319, new_AGEMA_signal_16318, RoundReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_5028, new_AGEMA_signal_5027, new_AGEMA_signal_5026, RoundInput[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16794, new_AGEMA_signal_16793, new_AGEMA_signal_16792, RoundReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, new_AGEMA_signal_5035, RoundInput[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16326, new_AGEMA_signal_16325, new_AGEMA_signal_16324, RoundReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_5046, new_AGEMA_signal_5045, new_AGEMA_signal_5044, RoundInput[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16800, new_AGEMA_signal_16799, new_AGEMA_signal_16798, RoundReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, new_AGEMA_signal_5053, RoundInput[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16806, new_AGEMA_signal_16805, new_AGEMA_signal_16804, RoundReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_5064, new_AGEMA_signal_5063, new_AGEMA_signal_5062, RoundInput[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16332, new_AGEMA_signal_16331, new_AGEMA_signal_16330, RoundReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, new_AGEMA_signal_5071, RoundInput[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16338, new_AGEMA_signal_16337, new_AGEMA_signal_16336, RoundReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_5082, new_AGEMA_signal_5081, new_AGEMA_signal_5080, RoundInput[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16344, new_AGEMA_signal_16343, new_AGEMA_signal_16342, RoundReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, new_AGEMA_signal_5089, RoundInput[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16350, new_AGEMA_signal_16349, new_AGEMA_signal_16348, RoundReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, new_AGEMA_signal_5107, RoundInput[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16812, new_AGEMA_signal_16811, new_AGEMA_signal_16810, RoundReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_5118, new_AGEMA_signal_5117, new_AGEMA_signal_5116, RoundInput[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16356, new_AGEMA_signal_16355, new_AGEMA_signal_16354, RoundReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, new_AGEMA_signal_5125, RoundInput[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16818, new_AGEMA_signal_16817, new_AGEMA_signal_16816, RoundReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_5136, new_AGEMA_signal_5135, new_AGEMA_signal_5134, RoundInput[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16824, new_AGEMA_signal_16823, new_AGEMA_signal_16822, RoundReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, new_AGEMA_signal_5143, RoundInput[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16362, new_AGEMA_signal_16361, new_AGEMA_signal_16360, RoundReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_5154, new_AGEMA_signal_5153, new_AGEMA_signal_5152, RoundInput[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16368, new_AGEMA_signal_16367, new_AGEMA_signal_16366, RoundReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, new_AGEMA_signal_5161, RoundInput[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16374, new_AGEMA_signal_16373, new_AGEMA_signal_16372, RoundReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_5172, new_AGEMA_signal_5171, new_AGEMA_signal_5170, RoundInput[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16380, new_AGEMA_signal_16379, new_AGEMA_signal_16378, RoundReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, new_AGEMA_signal_5179, RoundInput[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16830, new_AGEMA_signal_16829, new_AGEMA_signal_16828, RoundReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_5190, new_AGEMA_signal_5189, new_AGEMA_signal_5188, RoundInput[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16386, new_AGEMA_signal_16385, new_AGEMA_signal_16384, RoundReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_5208, new_AGEMA_signal_5207, new_AGEMA_signal_5206, RoundInput[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16836, new_AGEMA_signal_16835, new_AGEMA_signal_16834, RoundReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_5217, new_AGEMA_signal_5216, new_AGEMA_signal_5215, RoundInput[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16842, new_AGEMA_signal_16841, new_AGEMA_signal_16840, RoundReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5226, new_AGEMA_signal_5225, new_AGEMA_signal_5224, RoundInput[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16392, new_AGEMA_signal_16391, new_AGEMA_signal_16390, RoundReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5235, new_AGEMA_signal_5234, new_AGEMA_signal_5233, RoundInput[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16398, new_AGEMA_signal_16397, new_AGEMA_signal_16396, RoundReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5244, new_AGEMA_signal_5243, new_AGEMA_signal_5242, RoundInput[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16404, new_AGEMA_signal_16403, new_AGEMA_signal_16402, RoundReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5253, new_AGEMA_signal_5252, new_AGEMA_signal_5251, RoundInput[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16410, new_AGEMA_signal_16409, new_AGEMA_signal_16408, RoundReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5262, new_AGEMA_signal_5261, new_AGEMA_signal_5260, RoundInput[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16848, new_AGEMA_signal_16847, new_AGEMA_signal_16846, RoundReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5271, new_AGEMA_signal_5270, new_AGEMA_signal_5269, RoundInput[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16416, new_AGEMA_signal_16415, new_AGEMA_signal_16414, RoundReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5280, new_AGEMA_signal_5279, new_AGEMA_signal_5278, RoundInput[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16854, new_AGEMA_signal_16853, new_AGEMA_signal_16852, RoundReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5289, new_AGEMA_signal_5288, new_AGEMA_signal_5287, RoundInput[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16860, new_AGEMA_signal_16859, new_AGEMA_signal_16858, RoundReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5307, new_AGEMA_signal_5306, new_AGEMA_signal_5305, RoundInput[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16422, new_AGEMA_signal_16421, new_AGEMA_signal_16420, RoundReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5316, new_AGEMA_signal_5315, new_AGEMA_signal_5314, RoundInput[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16428, new_AGEMA_signal_16427, new_AGEMA_signal_16426, RoundReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5325, new_AGEMA_signal_5324, new_AGEMA_signal_5323, RoundInput[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16434, new_AGEMA_signal_16433, new_AGEMA_signal_16432, RoundReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5334, new_AGEMA_signal_5333, new_AGEMA_signal_5332, RoundInput[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16440, new_AGEMA_signal_16439, new_AGEMA_signal_16438, RoundReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5343, new_AGEMA_signal_5342, new_AGEMA_signal_5341, RoundInput[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16866, new_AGEMA_signal_16865, new_AGEMA_signal_16864, RoundReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5352, new_AGEMA_signal_5351, new_AGEMA_signal_5350, RoundInput[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16446, new_AGEMA_signal_16445, new_AGEMA_signal_16444, RoundReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5361, new_AGEMA_signal_5360, new_AGEMA_signal_5359, RoundInput[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16872, new_AGEMA_signal_16871, new_AGEMA_signal_16870, RoundReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5370, new_AGEMA_signal_5369, new_AGEMA_signal_5368, RoundInput[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16878, new_AGEMA_signal_16877, new_AGEMA_signal_16876, RoundReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5379, new_AGEMA_signal_5378, new_AGEMA_signal_5377, RoundInput[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16452, new_AGEMA_signal_16451, new_AGEMA_signal_16450, RoundReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5388, new_AGEMA_signal_5387, new_AGEMA_signal_5386, RoundInput[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16458, new_AGEMA_signal_16457, new_AGEMA_signal_16456, RoundReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5406, new_AGEMA_signal_5405, new_AGEMA_signal_5404, RoundInput[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16464, new_AGEMA_signal_16463, new_AGEMA_signal_16462, RoundReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5415, new_AGEMA_signal_5414, new_AGEMA_signal_5413, RoundInput[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16470, new_AGEMA_signal_16469, new_AGEMA_signal_16468, RoundReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5424, new_AGEMA_signal_5423, new_AGEMA_signal_5422, RoundInput[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16884, new_AGEMA_signal_16883, new_AGEMA_signal_16882, RoundReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5433, new_AGEMA_signal_5432, new_AGEMA_signal_5431, RoundInput[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16476, new_AGEMA_signal_16475, new_AGEMA_signal_16474, RoundReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5442, new_AGEMA_signal_5441, new_AGEMA_signal_5440, RoundInput[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16890, new_AGEMA_signal_16889, new_AGEMA_signal_16888, RoundReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5451, new_AGEMA_signal_5450, new_AGEMA_signal_5449, RoundInput[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16896, new_AGEMA_signal_16895, new_AGEMA_signal_16894, RoundReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5460, new_AGEMA_signal_5459, new_AGEMA_signal_5458, RoundInput[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16482, new_AGEMA_signal_16481, new_AGEMA_signal_16480, RoundReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5469, new_AGEMA_signal_5468, new_AGEMA_signal_5467, RoundInput[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16488, new_AGEMA_signal_16487, new_AGEMA_signal_16486, RoundReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5478, new_AGEMA_signal_5477, new_AGEMA_signal_5476, RoundInput[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16494, new_AGEMA_signal_16493, new_AGEMA_signal_16492, RoundReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5487, new_AGEMA_signal_5486, new_AGEMA_signal_5485, RoundInput[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16500, new_AGEMA_signal_16499, new_AGEMA_signal_16498, RoundReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5505, new_AGEMA_signal_5504, new_AGEMA_signal_5503, RoundInput[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16902, new_AGEMA_signal_16901, new_AGEMA_signal_16900, RoundReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5514, new_AGEMA_signal_5513, new_AGEMA_signal_5512, RoundInput[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16506, new_AGEMA_signal_16505, new_AGEMA_signal_16504, RoundReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5523, new_AGEMA_signal_5522, new_AGEMA_signal_5521, RoundInput[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16908, new_AGEMA_signal_16907, new_AGEMA_signal_16906, RoundReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5532, new_AGEMA_signal_5531, new_AGEMA_signal_5530, RoundInput[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16914, new_AGEMA_signal_16913, new_AGEMA_signal_16912, RoundReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5541, new_AGEMA_signal_5540, new_AGEMA_signal_5539, RoundInput[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16512, new_AGEMA_signal_16511, new_AGEMA_signal_16510, RoundReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5550, new_AGEMA_signal_5549, new_AGEMA_signal_5548, RoundInput[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16518, new_AGEMA_signal_16517, new_AGEMA_signal_16516, RoundReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5559, new_AGEMA_signal_5558, new_AGEMA_signal_5557, RoundInput[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16524, new_AGEMA_signal_16523, new_AGEMA_signal_16522, RoundReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5568, new_AGEMA_signal_5567, new_AGEMA_signal_5566, RoundInput[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16530, new_AGEMA_signal_16529, new_AGEMA_signal_16528, RoundReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5577, new_AGEMA_signal_5576, new_AGEMA_signal_5575, RoundInput[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16920, new_AGEMA_signal_16919, new_AGEMA_signal_16918, RoundReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5586, new_AGEMA_signal_5585, new_AGEMA_signal_5584, RoundInput[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16536, new_AGEMA_signal_16535, new_AGEMA_signal_16534, RoundReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5604, new_AGEMA_signal_5603, new_AGEMA_signal_5602, RoundInput[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16926, new_AGEMA_signal_16925, new_AGEMA_signal_16924, RoundReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5613, new_AGEMA_signal_5612, new_AGEMA_signal_5611, RoundInput[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16932, new_AGEMA_signal_16931, new_AGEMA_signal_16930, RoundReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5622, new_AGEMA_signal_5621, new_AGEMA_signal_5620, RoundInput[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16542, new_AGEMA_signal_16541, new_AGEMA_signal_16540, RoundReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5631, new_AGEMA_signal_5630, new_AGEMA_signal_5629, RoundInput[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16548, new_AGEMA_signal_16547, new_AGEMA_signal_16546, RoundReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5640, new_AGEMA_signal_5639, new_AGEMA_signal_5638, RoundInput[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16554, new_AGEMA_signal_16553, new_AGEMA_signal_16552, RoundReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5649, new_AGEMA_signal_5648, new_AGEMA_signal_5647, RoundInput[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16560, new_AGEMA_signal_16559, new_AGEMA_signal_16558, RoundReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5658, new_AGEMA_signal_5657, new_AGEMA_signal_5656, RoundInput[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16938, new_AGEMA_signal_16937, new_AGEMA_signal_16936, RoundReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5667, new_AGEMA_signal_5666, new_AGEMA_signal_5665, RoundInput[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16566, new_AGEMA_signal_16565, new_AGEMA_signal_16564, RoundReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5676, new_AGEMA_signal_5675, new_AGEMA_signal_5674, RoundInput[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16944, new_AGEMA_signal_16943, new_AGEMA_signal_16942, RoundReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5685, new_AGEMA_signal_5684, new_AGEMA_signal_5683, RoundInput[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16950, new_AGEMA_signal_16949, new_AGEMA_signal_16948, RoundReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4560, new_AGEMA_signal_4559, new_AGEMA_signal_4558, RoundInput[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16572, new_AGEMA_signal_16571, new_AGEMA_signal_16570, RoundReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, new_AGEMA_signal_4567, RoundInput[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16578, new_AGEMA_signal_16577, new_AGEMA_signal_16576, RoundReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4578, new_AGEMA_signal_4577, new_AGEMA_signal_4576, RoundInput[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16584, new_AGEMA_signal_16583, new_AGEMA_signal_16582, RoundReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, new_AGEMA_signal_4585, RoundInput[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16590, new_AGEMA_signal_16589, new_AGEMA_signal_16588, RoundReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4596, new_AGEMA_signal_4595, new_AGEMA_signal_4594, RoundInput[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16956, new_AGEMA_signal_16955, new_AGEMA_signal_16954, RoundReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, new_AGEMA_signal_4603, RoundInput[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16596, new_AGEMA_signal_16595, new_AGEMA_signal_16594, RoundReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4614, new_AGEMA_signal_4613, new_AGEMA_signal_4612, RoundInput[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16962, new_AGEMA_signal_16961, new_AGEMA_signal_16960, RoundReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, new_AGEMA_signal_4621, RoundInput[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16968, new_AGEMA_signal_16967, new_AGEMA_signal_16966, RoundReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4632, new_AGEMA_signal_4631, new_AGEMA_signal_4630, RoundInput[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16602, new_AGEMA_signal_16601, new_AGEMA_signal_16600, RoundReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, new_AGEMA_signal_4639, RoundInput[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16608, new_AGEMA_signal_16607, new_AGEMA_signal_16606, RoundReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, new_AGEMA_signal_4657, RoundInput[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16614, new_AGEMA_signal_16613, new_AGEMA_signal_16612, RoundReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4668, new_AGEMA_signal_4667, new_AGEMA_signal_4666, RoundInput[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16620, new_AGEMA_signal_16619, new_AGEMA_signal_16618, RoundReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, new_AGEMA_signal_4675, RoundInput[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16974, new_AGEMA_signal_16973, new_AGEMA_signal_16972, RoundReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4686, new_AGEMA_signal_4685, new_AGEMA_signal_4684, RoundInput[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16626, new_AGEMA_signal_16625, new_AGEMA_signal_16624, RoundReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, new_AGEMA_signal_4693, RoundInput[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16980, new_AGEMA_signal_16979, new_AGEMA_signal_16978, RoundReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4704, new_AGEMA_signal_4703, new_AGEMA_signal_4702, RoundInput[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16986, new_AGEMA_signal_16985, new_AGEMA_signal_16984, RoundReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, new_AGEMA_signal_4711, RoundInput[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16632, new_AGEMA_signal_16631, new_AGEMA_signal_16630, RoundReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4722, new_AGEMA_signal_4721, new_AGEMA_signal_4720, RoundInput[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16638, new_AGEMA_signal_16637, new_AGEMA_signal_16636, RoundReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, new_AGEMA_signal_4729, RoundInput[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16644, new_AGEMA_signal_16643, new_AGEMA_signal_16642, RoundReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4740, new_AGEMA_signal_4739, new_AGEMA_signal_4738, RoundInput[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16650, new_AGEMA_signal_16649, new_AGEMA_signal_16648, RoundReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4758, new_AGEMA_signal_4757, new_AGEMA_signal_4756, RoundInput[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16992, new_AGEMA_signal_16991, new_AGEMA_signal_16990, RoundReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, new_AGEMA_signal_4765, RoundInput[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16656, new_AGEMA_signal_16655, new_AGEMA_signal_16654, RoundReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4776, new_AGEMA_signal_4775, new_AGEMA_signal_4774, RoundInput[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16998, new_AGEMA_signal_16997, new_AGEMA_signal_16996, RoundReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, new_AGEMA_signal_4783, RoundInput[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_17004, new_AGEMA_signal_17003, new_AGEMA_signal_17002, RoundReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4794, new_AGEMA_signal_4793, new_AGEMA_signal_4792, RoundInput[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16662, new_AGEMA_signal_16661, new_AGEMA_signal_16660, RoundReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, new_AGEMA_signal_4801, RoundInput[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16668, new_AGEMA_signal_16667, new_AGEMA_signal_16666, RoundReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4812, new_AGEMA_signal_4811, new_AGEMA_signal_4810, RoundInput[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) RoundReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16674, new_AGEMA_signal_16673, new_AGEMA_signal_16672, RoundReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, new_AGEMA_signal_4819, RoundInput[127]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_0_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15198, new_AGEMA_signal_15197, new_AGEMA_signal_15196, KeyReg_Inst_ff_SDE_0_next_state}), .Q ({new_AGEMA_signal_4554, new_AGEMA_signal_4553, new_AGEMA_signal_4552, RoundKey[0]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_1_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15861, new_AGEMA_signal_15860, new_AGEMA_signal_15859, KeyReg_Inst_ff_SDE_1_next_state}), .Q ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, new_AGEMA_signal_4903, RoundKey[1]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_2_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15867, new_AGEMA_signal_15866, new_AGEMA_signal_15865, KeyReg_Inst_ff_SDE_2_next_state}), .Q ({new_AGEMA_signal_5004, new_AGEMA_signal_5003, new_AGEMA_signal_5002, RoundKey[2]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_3_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15873, new_AGEMA_signal_15872, new_AGEMA_signal_15871, KeyReg_Inst_ff_SDE_3_next_state}), .Q ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, new_AGEMA_signal_5101, RoundKey[3]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_4_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15879, new_AGEMA_signal_15878, new_AGEMA_signal_15877, KeyReg_Inst_ff_SDE_4_next_state}), .Q ({new_AGEMA_signal_5202, new_AGEMA_signal_5201, new_AGEMA_signal_5200, RoundKey[4]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_5_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15885, new_AGEMA_signal_15884, new_AGEMA_signal_15883, KeyReg_Inst_ff_SDE_5_next_state}), .Q ({new_AGEMA_signal_5301, new_AGEMA_signal_5300, new_AGEMA_signal_5299, RoundKey[5]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_6_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15891, new_AGEMA_signal_15890, new_AGEMA_signal_15889, KeyReg_Inst_ff_SDE_6_next_state}), .Q ({new_AGEMA_signal_5400, new_AGEMA_signal_5399, new_AGEMA_signal_5398, RoundKey[6]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_7_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15897, new_AGEMA_signal_15896, new_AGEMA_signal_15895, KeyReg_Inst_ff_SDE_7_next_state}), .Q ({new_AGEMA_signal_5499, new_AGEMA_signal_5498, new_AGEMA_signal_5497, RoundKey[7]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_8_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15204, new_AGEMA_signal_15203, new_AGEMA_signal_15202, KeyReg_Inst_ff_SDE_8_next_state}), .Q ({new_AGEMA_signal_5598, new_AGEMA_signal_5597, new_AGEMA_signal_5596, RoundKey[8]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_9_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15903, new_AGEMA_signal_15902, new_AGEMA_signal_15901, KeyReg_Inst_ff_SDE_9_next_state}), .Q ({new_AGEMA_signal_5697, new_AGEMA_signal_5696, new_AGEMA_signal_5695, RoundKey[9]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_10_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15909, new_AGEMA_signal_15908, new_AGEMA_signal_15907, KeyReg_Inst_ff_SDE_10_next_state}), .Q ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, new_AGEMA_signal_4651, RoundKey[10]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_11_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15915, new_AGEMA_signal_15914, new_AGEMA_signal_15913, KeyReg_Inst_ff_SDE_11_next_state}), .Q ({new_AGEMA_signal_4752, new_AGEMA_signal_4751, new_AGEMA_signal_4750, RoundKey[11]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_12_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15921, new_AGEMA_signal_15920, new_AGEMA_signal_15919, KeyReg_Inst_ff_SDE_12_next_state}), .Q ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, new_AGEMA_signal_4831, RoundKey[12]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_13_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15927, new_AGEMA_signal_15926, new_AGEMA_signal_15925, KeyReg_Inst_ff_SDE_13_next_state}), .Q ({new_AGEMA_signal_4842, new_AGEMA_signal_4841, new_AGEMA_signal_4840, RoundKey[13]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_14_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15933, new_AGEMA_signal_15932, new_AGEMA_signal_15931, KeyReg_Inst_ff_SDE_14_next_state}), .Q ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, new_AGEMA_signal_4849, RoundKey[14]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_15_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15939, new_AGEMA_signal_15938, new_AGEMA_signal_15937, KeyReg_Inst_ff_SDE_15_next_state}), .Q ({new_AGEMA_signal_4860, new_AGEMA_signal_4859, new_AGEMA_signal_4858, RoundKey[15]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_16_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15210, new_AGEMA_signal_15209, new_AGEMA_signal_15208, KeyReg_Inst_ff_SDE_16_next_state}), .Q ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, new_AGEMA_signal_4867, RoundKey[16]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_17_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15945, new_AGEMA_signal_15944, new_AGEMA_signal_15943, KeyReg_Inst_ff_SDE_17_next_state}), .Q ({new_AGEMA_signal_4878, new_AGEMA_signal_4877, new_AGEMA_signal_4876, RoundKey[17]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_18_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15951, new_AGEMA_signal_15950, new_AGEMA_signal_15949, KeyReg_Inst_ff_SDE_18_next_state}), .Q ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, new_AGEMA_signal_4885, RoundKey[18]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_19_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15957, new_AGEMA_signal_15956, new_AGEMA_signal_15955, KeyReg_Inst_ff_SDE_19_next_state}), .Q ({new_AGEMA_signal_4896, new_AGEMA_signal_4895, new_AGEMA_signal_4894, RoundKey[19]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_20_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15963, new_AGEMA_signal_15962, new_AGEMA_signal_15961, KeyReg_Inst_ff_SDE_20_next_state}), .Q ({new_AGEMA_signal_4914, new_AGEMA_signal_4913, new_AGEMA_signal_4912, RoundKey[20]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_21_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15969, new_AGEMA_signal_15968, new_AGEMA_signal_15967, KeyReg_Inst_ff_SDE_21_next_state}), .Q ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, new_AGEMA_signal_4921, RoundKey[21]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_22_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15975, new_AGEMA_signal_15974, new_AGEMA_signal_15973, KeyReg_Inst_ff_SDE_22_next_state}), .Q ({new_AGEMA_signal_4932, new_AGEMA_signal_4931, new_AGEMA_signal_4930, RoundKey[22]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_23_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15981, new_AGEMA_signal_15980, new_AGEMA_signal_15979, KeyReg_Inst_ff_SDE_23_next_state}), .Q ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, new_AGEMA_signal_4939, RoundKey[23]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_24_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15987, new_AGEMA_signal_15986, new_AGEMA_signal_15985, KeyReg_Inst_ff_SDE_24_next_state}), .Q ({new_AGEMA_signal_4950, new_AGEMA_signal_4949, new_AGEMA_signal_4948, RoundKey[24]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_25_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16680, new_AGEMA_signal_16679, new_AGEMA_signal_16678, KeyReg_Inst_ff_SDE_25_next_state}), .Q ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, new_AGEMA_signal_4957, RoundKey[25]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_26_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16686, new_AGEMA_signal_16685, new_AGEMA_signal_16684, KeyReg_Inst_ff_SDE_26_next_state}), .Q ({new_AGEMA_signal_4968, new_AGEMA_signal_4967, new_AGEMA_signal_4966, RoundKey[26]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_27_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16692, new_AGEMA_signal_16691, new_AGEMA_signal_16690, KeyReg_Inst_ff_SDE_27_next_state}), .Q ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, new_AGEMA_signal_4975, RoundKey[27]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_28_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16698, new_AGEMA_signal_16697, new_AGEMA_signal_16696, KeyReg_Inst_ff_SDE_28_next_state}), .Q ({new_AGEMA_signal_4986, new_AGEMA_signal_4985, new_AGEMA_signal_4984, RoundKey[28]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_29_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16704, new_AGEMA_signal_16703, new_AGEMA_signal_16702, KeyReg_Inst_ff_SDE_29_next_state}), .Q ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, new_AGEMA_signal_4993, RoundKey[29]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_30_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16710, new_AGEMA_signal_16709, new_AGEMA_signal_16708, KeyReg_Inst_ff_SDE_30_next_state}), .Q ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, new_AGEMA_signal_5011, RoundKey[30]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_31_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16716, new_AGEMA_signal_16715, new_AGEMA_signal_16714, KeyReg_Inst_ff_SDE_31_next_state}), .Q ({new_AGEMA_signal_5022, new_AGEMA_signal_5021, new_AGEMA_signal_5020, RoundKey[31]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_32_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14526, new_AGEMA_signal_14525, new_AGEMA_signal_14524, KeyReg_Inst_ff_SDE_32_next_state}), .Q ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, new_AGEMA_signal_5029, RoundKey[32]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_33_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15216, new_AGEMA_signal_15215, new_AGEMA_signal_15214, KeyReg_Inst_ff_SDE_33_next_state}), .Q ({new_AGEMA_signal_5040, new_AGEMA_signal_5039, new_AGEMA_signal_5038, RoundKey[33]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_34_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15222, new_AGEMA_signal_15221, new_AGEMA_signal_15220, KeyReg_Inst_ff_SDE_34_next_state}), .Q ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, new_AGEMA_signal_5047, RoundKey[34]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_35_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15228, new_AGEMA_signal_15227, new_AGEMA_signal_15226, KeyReg_Inst_ff_SDE_35_next_state}), .Q ({new_AGEMA_signal_5058, new_AGEMA_signal_5057, new_AGEMA_signal_5056, RoundKey[35]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_36_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15234, new_AGEMA_signal_15233, new_AGEMA_signal_15232, KeyReg_Inst_ff_SDE_36_next_state}), .Q ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, new_AGEMA_signal_5065, RoundKey[36]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_37_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15240, new_AGEMA_signal_15239, new_AGEMA_signal_15238, KeyReg_Inst_ff_SDE_37_next_state}), .Q ({new_AGEMA_signal_5076, new_AGEMA_signal_5075, new_AGEMA_signal_5074, RoundKey[37]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_38_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15246, new_AGEMA_signal_15245, new_AGEMA_signal_15244, KeyReg_Inst_ff_SDE_38_next_state}), .Q ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, new_AGEMA_signal_5083, RoundKey[38]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_39_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15252, new_AGEMA_signal_15251, new_AGEMA_signal_15250, KeyReg_Inst_ff_SDE_39_next_state}), .Q ({new_AGEMA_signal_5094, new_AGEMA_signal_5093, new_AGEMA_signal_5092, RoundKey[39]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_40_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14532, new_AGEMA_signal_14531, new_AGEMA_signal_14530, KeyReg_Inst_ff_SDE_40_next_state}), .Q ({new_AGEMA_signal_5112, new_AGEMA_signal_5111, new_AGEMA_signal_5110, RoundKey[40]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_41_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15258, new_AGEMA_signal_15257, new_AGEMA_signal_15256, KeyReg_Inst_ff_SDE_41_next_state}), .Q ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, new_AGEMA_signal_5119, RoundKey[41]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_42_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15264, new_AGEMA_signal_15263, new_AGEMA_signal_15262, KeyReg_Inst_ff_SDE_42_next_state}), .Q ({new_AGEMA_signal_5130, new_AGEMA_signal_5129, new_AGEMA_signal_5128, RoundKey[42]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_43_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15270, new_AGEMA_signal_15269, new_AGEMA_signal_15268, KeyReg_Inst_ff_SDE_43_next_state}), .Q ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, new_AGEMA_signal_5137, RoundKey[43]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_44_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15276, new_AGEMA_signal_15275, new_AGEMA_signal_15274, KeyReg_Inst_ff_SDE_44_next_state}), .Q ({new_AGEMA_signal_5148, new_AGEMA_signal_5147, new_AGEMA_signal_5146, RoundKey[44]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_45_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15282, new_AGEMA_signal_15281, new_AGEMA_signal_15280, KeyReg_Inst_ff_SDE_45_next_state}), .Q ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, new_AGEMA_signal_5155, RoundKey[45]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_46_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15288, new_AGEMA_signal_15287, new_AGEMA_signal_15286, KeyReg_Inst_ff_SDE_46_next_state}), .Q ({new_AGEMA_signal_5166, new_AGEMA_signal_5165, new_AGEMA_signal_5164, RoundKey[46]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_47_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15294, new_AGEMA_signal_15293, new_AGEMA_signal_15292, KeyReg_Inst_ff_SDE_47_next_state}), .Q ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, new_AGEMA_signal_5173, RoundKey[47]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_48_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14538, new_AGEMA_signal_14537, new_AGEMA_signal_14536, KeyReg_Inst_ff_SDE_48_next_state}), .Q ({new_AGEMA_signal_5184, new_AGEMA_signal_5183, new_AGEMA_signal_5182, RoundKey[48]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_49_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15300, new_AGEMA_signal_15299, new_AGEMA_signal_15298, KeyReg_Inst_ff_SDE_49_next_state}), .Q ({new_AGEMA_signal_5193, new_AGEMA_signal_5192, new_AGEMA_signal_5191, RoundKey[49]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_50_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15306, new_AGEMA_signal_15305, new_AGEMA_signal_15304, KeyReg_Inst_ff_SDE_50_next_state}), .Q ({new_AGEMA_signal_5211, new_AGEMA_signal_5210, new_AGEMA_signal_5209, RoundKey[50]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_51_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15312, new_AGEMA_signal_15311, new_AGEMA_signal_15310, KeyReg_Inst_ff_SDE_51_next_state}), .Q ({new_AGEMA_signal_5220, new_AGEMA_signal_5219, new_AGEMA_signal_5218, RoundKey[51]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_52_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15318, new_AGEMA_signal_15317, new_AGEMA_signal_15316, KeyReg_Inst_ff_SDE_52_next_state}), .Q ({new_AGEMA_signal_5229, new_AGEMA_signal_5228, new_AGEMA_signal_5227, RoundKey[52]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_53_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15324, new_AGEMA_signal_15323, new_AGEMA_signal_15322, KeyReg_Inst_ff_SDE_53_next_state}), .Q ({new_AGEMA_signal_5238, new_AGEMA_signal_5237, new_AGEMA_signal_5236, RoundKey[53]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_54_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15330, new_AGEMA_signal_15329, new_AGEMA_signal_15328, KeyReg_Inst_ff_SDE_54_next_state}), .Q ({new_AGEMA_signal_5247, new_AGEMA_signal_5246, new_AGEMA_signal_5245, RoundKey[54]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_55_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15336, new_AGEMA_signal_15335, new_AGEMA_signal_15334, KeyReg_Inst_ff_SDE_55_next_state}), .Q ({new_AGEMA_signal_5256, new_AGEMA_signal_5255, new_AGEMA_signal_5254, RoundKey[55]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_56_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15342, new_AGEMA_signal_15341, new_AGEMA_signal_15340, KeyReg_Inst_ff_SDE_56_next_state}), .Q ({new_AGEMA_signal_5265, new_AGEMA_signal_5264, new_AGEMA_signal_5263, RoundKey[56]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_57_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15993, new_AGEMA_signal_15992, new_AGEMA_signal_15991, KeyReg_Inst_ff_SDE_57_next_state}), .Q ({new_AGEMA_signal_5274, new_AGEMA_signal_5273, new_AGEMA_signal_5272, RoundKey[57]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_58_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15999, new_AGEMA_signal_15998, new_AGEMA_signal_15997, KeyReg_Inst_ff_SDE_58_next_state}), .Q ({new_AGEMA_signal_5283, new_AGEMA_signal_5282, new_AGEMA_signal_5281, RoundKey[58]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_59_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16005, new_AGEMA_signal_16004, new_AGEMA_signal_16003, KeyReg_Inst_ff_SDE_59_next_state}), .Q ({new_AGEMA_signal_5292, new_AGEMA_signal_5291, new_AGEMA_signal_5290, RoundKey[59]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_60_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16011, new_AGEMA_signal_16010, new_AGEMA_signal_16009, KeyReg_Inst_ff_SDE_60_next_state}), .Q ({new_AGEMA_signal_5310, new_AGEMA_signal_5309, new_AGEMA_signal_5308, RoundKey[60]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_61_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16017, new_AGEMA_signal_16016, new_AGEMA_signal_16015, KeyReg_Inst_ff_SDE_61_next_state}), .Q ({new_AGEMA_signal_5319, new_AGEMA_signal_5318, new_AGEMA_signal_5317, RoundKey[61]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_62_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16023, new_AGEMA_signal_16022, new_AGEMA_signal_16021, KeyReg_Inst_ff_SDE_62_next_state}), .Q ({new_AGEMA_signal_5328, new_AGEMA_signal_5327, new_AGEMA_signal_5326, RoundKey[62]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_63_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_16029, new_AGEMA_signal_16028, new_AGEMA_signal_16027, KeyReg_Inst_ff_SDE_63_next_state}), .Q ({new_AGEMA_signal_5337, new_AGEMA_signal_5336, new_AGEMA_signal_5335, RoundKey[63]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_64_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13896, new_AGEMA_signal_13895, new_AGEMA_signal_13894, KeyReg_Inst_ff_SDE_64_next_state}), .Q ({new_AGEMA_signal_5346, new_AGEMA_signal_5345, new_AGEMA_signal_5344, RoundKey[64]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_65_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14544, new_AGEMA_signal_14543, new_AGEMA_signal_14542, KeyReg_Inst_ff_SDE_65_next_state}), .Q ({new_AGEMA_signal_5355, new_AGEMA_signal_5354, new_AGEMA_signal_5353, RoundKey[65]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_66_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14550, new_AGEMA_signal_14549, new_AGEMA_signal_14548, KeyReg_Inst_ff_SDE_66_next_state}), .Q ({new_AGEMA_signal_5364, new_AGEMA_signal_5363, new_AGEMA_signal_5362, RoundKey[66]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_67_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14556, new_AGEMA_signal_14555, new_AGEMA_signal_14554, KeyReg_Inst_ff_SDE_67_next_state}), .Q ({new_AGEMA_signal_5373, new_AGEMA_signal_5372, new_AGEMA_signal_5371, RoundKey[67]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_68_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14562, new_AGEMA_signal_14561, new_AGEMA_signal_14560, KeyReg_Inst_ff_SDE_68_next_state}), .Q ({new_AGEMA_signal_5382, new_AGEMA_signal_5381, new_AGEMA_signal_5380, RoundKey[68]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_69_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14568, new_AGEMA_signal_14567, new_AGEMA_signal_14566, KeyReg_Inst_ff_SDE_69_next_state}), .Q ({new_AGEMA_signal_5391, new_AGEMA_signal_5390, new_AGEMA_signal_5389, RoundKey[69]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_70_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14574, new_AGEMA_signal_14573, new_AGEMA_signal_14572, KeyReg_Inst_ff_SDE_70_next_state}), .Q ({new_AGEMA_signal_5409, new_AGEMA_signal_5408, new_AGEMA_signal_5407, RoundKey[70]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_71_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14580, new_AGEMA_signal_14579, new_AGEMA_signal_14578, KeyReg_Inst_ff_SDE_71_next_state}), .Q ({new_AGEMA_signal_5418, new_AGEMA_signal_5417, new_AGEMA_signal_5416, RoundKey[71]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_72_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13902, new_AGEMA_signal_13901, new_AGEMA_signal_13900, KeyReg_Inst_ff_SDE_72_next_state}), .Q ({new_AGEMA_signal_5427, new_AGEMA_signal_5426, new_AGEMA_signal_5425, RoundKey[72]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_73_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14586, new_AGEMA_signal_14585, new_AGEMA_signal_14584, KeyReg_Inst_ff_SDE_73_next_state}), .Q ({new_AGEMA_signal_5436, new_AGEMA_signal_5435, new_AGEMA_signal_5434, RoundKey[73]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_74_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14592, new_AGEMA_signal_14591, new_AGEMA_signal_14590, KeyReg_Inst_ff_SDE_74_next_state}), .Q ({new_AGEMA_signal_5445, new_AGEMA_signal_5444, new_AGEMA_signal_5443, RoundKey[74]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_75_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14598, new_AGEMA_signal_14597, new_AGEMA_signal_14596, KeyReg_Inst_ff_SDE_75_next_state}), .Q ({new_AGEMA_signal_5454, new_AGEMA_signal_5453, new_AGEMA_signal_5452, RoundKey[75]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_76_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14604, new_AGEMA_signal_14603, new_AGEMA_signal_14602, KeyReg_Inst_ff_SDE_76_next_state}), .Q ({new_AGEMA_signal_5463, new_AGEMA_signal_5462, new_AGEMA_signal_5461, RoundKey[76]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_77_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14610, new_AGEMA_signal_14609, new_AGEMA_signal_14608, KeyReg_Inst_ff_SDE_77_next_state}), .Q ({new_AGEMA_signal_5472, new_AGEMA_signal_5471, new_AGEMA_signal_5470, RoundKey[77]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_78_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14616, new_AGEMA_signal_14615, new_AGEMA_signal_14614, KeyReg_Inst_ff_SDE_78_next_state}), .Q ({new_AGEMA_signal_5481, new_AGEMA_signal_5480, new_AGEMA_signal_5479, RoundKey[78]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_79_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14622, new_AGEMA_signal_14621, new_AGEMA_signal_14620, KeyReg_Inst_ff_SDE_79_next_state}), .Q ({new_AGEMA_signal_5490, new_AGEMA_signal_5489, new_AGEMA_signal_5488, RoundKey[79]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_80_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13908, new_AGEMA_signal_13907, new_AGEMA_signal_13906, KeyReg_Inst_ff_SDE_80_next_state}), .Q ({new_AGEMA_signal_5508, new_AGEMA_signal_5507, new_AGEMA_signal_5506, RoundKey[80]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_81_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14628, new_AGEMA_signal_14627, new_AGEMA_signal_14626, KeyReg_Inst_ff_SDE_81_next_state}), .Q ({new_AGEMA_signal_5517, new_AGEMA_signal_5516, new_AGEMA_signal_5515, RoundKey[81]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_82_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14634, new_AGEMA_signal_14633, new_AGEMA_signal_14632, KeyReg_Inst_ff_SDE_82_next_state}), .Q ({new_AGEMA_signal_5526, new_AGEMA_signal_5525, new_AGEMA_signal_5524, RoundKey[82]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_83_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14640, new_AGEMA_signal_14639, new_AGEMA_signal_14638, KeyReg_Inst_ff_SDE_83_next_state}), .Q ({new_AGEMA_signal_5535, new_AGEMA_signal_5534, new_AGEMA_signal_5533, RoundKey[83]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_84_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14646, new_AGEMA_signal_14645, new_AGEMA_signal_14644, KeyReg_Inst_ff_SDE_84_next_state}), .Q ({new_AGEMA_signal_5544, new_AGEMA_signal_5543, new_AGEMA_signal_5542, RoundKey[84]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_85_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14652, new_AGEMA_signal_14651, new_AGEMA_signal_14650, KeyReg_Inst_ff_SDE_85_next_state}), .Q ({new_AGEMA_signal_5553, new_AGEMA_signal_5552, new_AGEMA_signal_5551, RoundKey[85]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_86_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14658, new_AGEMA_signal_14657, new_AGEMA_signal_14656, KeyReg_Inst_ff_SDE_86_next_state}), .Q ({new_AGEMA_signal_5562, new_AGEMA_signal_5561, new_AGEMA_signal_5560, RoundKey[86]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_87_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14664, new_AGEMA_signal_14663, new_AGEMA_signal_14662, KeyReg_Inst_ff_SDE_87_next_state}), .Q ({new_AGEMA_signal_5571, new_AGEMA_signal_5570, new_AGEMA_signal_5569, RoundKey[87]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_88_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14670, new_AGEMA_signal_14669, new_AGEMA_signal_14668, KeyReg_Inst_ff_SDE_88_next_state}), .Q ({new_AGEMA_signal_5580, new_AGEMA_signal_5579, new_AGEMA_signal_5578, RoundKey[88]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_89_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15348, new_AGEMA_signal_15347, new_AGEMA_signal_15346, KeyReg_Inst_ff_SDE_89_next_state}), .Q ({new_AGEMA_signal_5589, new_AGEMA_signal_5588, new_AGEMA_signal_5587, RoundKey[89]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_90_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15354, new_AGEMA_signal_15353, new_AGEMA_signal_15352, KeyReg_Inst_ff_SDE_90_next_state}), .Q ({new_AGEMA_signal_5607, new_AGEMA_signal_5606, new_AGEMA_signal_5605, RoundKey[90]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_91_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15360, new_AGEMA_signal_15359, new_AGEMA_signal_15358, KeyReg_Inst_ff_SDE_91_next_state}), .Q ({new_AGEMA_signal_5616, new_AGEMA_signal_5615, new_AGEMA_signal_5614, RoundKey[91]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_92_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15366, new_AGEMA_signal_15365, new_AGEMA_signal_15364, KeyReg_Inst_ff_SDE_92_next_state}), .Q ({new_AGEMA_signal_5625, new_AGEMA_signal_5624, new_AGEMA_signal_5623, RoundKey[92]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_93_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15372, new_AGEMA_signal_15371, new_AGEMA_signal_15370, KeyReg_Inst_ff_SDE_93_next_state}), .Q ({new_AGEMA_signal_5634, new_AGEMA_signal_5633, new_AGEMA_signal_5632, RoundKey[93]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_94_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15378, new_AGEMA_signal_15377, new_AGEMA_signal_15376, KeyReg_Inst_ff_SDE_94_next_state}), .Q ({new_AGEMA_signal_5643, new_AGEMA_signal_5642, new_AGEMA_signal_5641, RoundKey[94]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_95_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_15384, new_AGEMA_signal_15383, new_AGEMA_signal_15382, KeyReg_Inst_ff_SDE_95_next_state}), .Q ({new_AGEMA_signal_5652, new_AGEMA_signal_5651, new_AGEMA_signal_5650, RoundKey[95]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_96_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13398, new_AGEMA_signal_13397, new_AGEMA_signal_13396, KeyReg_Inst_ff_SDE_96_next_state}), .Q ({new_AGEMA_signal_5661, new_AGEMA_signal_5660, new_AGEMA_signal_5659, RoundKey[96]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_97_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13914, new_AGEMA_signal_13913, new_AGEMA_signal_13912, KeyReg_Inst_ff_SDE_97_next_state}), .Q ({new_AGEMA_signal_5670, new_AGEMA_signal_5669, new_AGEMA_signal_5668, RoundKey[97]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_98_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13920, new_AGEMA_signal_13919, new_AGEMA_signal_13918, KeyReg_Inst_ff_SDE_98_next_state}), .Q ({new_AGEMA_signal_5679, new_AGEMA_signal_5678, new_AGEMA_signal_5677, RoundKey[98]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_99_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13926, new_AGEMA_signal_13925, new_AGEMA_signal_13924, KeyReg_Inst_ff_SDE_99_next_state}), .Q ({new_AGEMA_signal_5688, new_AGEMA_signal_5687, new_AGEMA_signal_5686, RoundKey[99]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_100_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13932, new_AGEMA_signal_13931, new_AGEMA_signal_13930, KeyReg_Inst_ff_SDE_100_next_state}), .Q ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, new_AGEMA_signal_4561, RoundKey[100]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_101_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13938, new_AGEMA_signal_13937, new_AGEMA_signal_13936, KeyReg_Inst_ff_SDE_101_next_state}), .Q ({new_AGEMA_signal_4572, new_AGEMA_signal_4571, new_AGEMA_signal_4570, RoundKey[101]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_102_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13944, new_AGEMA_signal_13943, new_AGEMA_signal_13942, KeyReg_Inst_ff_SDE_102_next_state}), .Q ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, new_AGEMA_signal_4579, RoundKey[102]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_103_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13950, new_AGEMA_signal_13949, new_AGEMA_signal_13948, KeyReg_Inst_ff_SDE_103_next_state}), .Q ({new_AGEMA_signal_4590, new_AGEMA_signal_4589, new_AGEMA_signal_4588, RoundKey[103]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_104_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13404, new_AGEMA_signal_13403, new_AGEMA_signal_13402, KeyReg_Inst_ff_SDE_104_next_state}), .Q ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, new_AGEMA_signal_4597, RoundKey[104]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_105_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13956, new_AGEMA_signal_13955, new_AGEMA_signal_13954, KeyReg_Inst_ff_SDE_105_next_state}), .Q ({new_AGEMA_signal_4608, new_AGEMA_signal_4607, new_AGEMA_signal_4606, RoundKey[105]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_106_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13962, new_AGEMA_signal_13961, new_AGEMA_signal_13960, KeyReg_Inst_ff_SDE_106_next_state}), .Q ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, new_AGEMA_signal_4615, RoundKey[106]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_107_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13968, new_AGEMA_signal_13967, new_AGEMA_signal_13966, KeyReg_Inst_ff_SDE_107_next_state}), .Q ({new_AGEMA_signal_4626, new_AGEMA_signal_4625, new_AGEMA_signal_4624, RoundKey[107]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_108_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13974, new_AGEMA_signal_13973, new_AGEMA_signal_13972, KeyReg_Inst_ff_SDE_108_next_state}), .Q ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, new_AGEMA_signal_4633, RoundKey[108]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_109_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13980, new_AGEMA_signal_13979, new_AGEMA_signal_13978, KeyReg_Inst_ff_SDE_109_next_state}), .Q ({new_AGEMA_signal_4644, new_AGEMA_signal_4643, new_AGEMA_signal_4642, RoundKey[109]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_110_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13986, new_AGEMA_signal_13985, new_AGEMA_signal_13984, KeyReg_Inst_ff_SDE_110_next_state}), .Q ({new_AGEMA_signal_4662, new_AGEMA_signal_4661, new_AGEMA_signal_4660, RoundKey[110]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_111_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13992, new_AGEMA_signal_13991, new_AGEMA_signal_13990, KeyReg_Inst_ff_SDE_111_next_state}), .Q ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, new_AGEMA_signal_4669, RoundKey[111]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_112_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13410, new_AGEMA_signal_13409, new_AGEMA_signal_13408, KeyReg_Inst_ff_SDE_112_next_state}), .Q ({new_AGEMA_signal_4680, new_AGEMA_signal_4679, new_AGEMA_signal_4678, RoundKey[112]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_113_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_13998, new_AGEMA_signal_13997, new_AGEMA_signal_13996, KeyReg_Inst_ff_SDE_113_next_state}), .Q ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, new_AGEMA_signal_4687, RoundKey[113]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_114_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14004, new_AGEMA_signal_14003, new_AGEMA_signal_14002, KeyReg_Inst_ff_SDE_114_next_state}), .Q ({new_AGEMA_signal_4698, new_AGEMA_signal_4697, new_AGEMA_signal_4696, RoundKey[114]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_115_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14010, new_AGEMA_signal_14009, new_AGEMA_signal_14008, KeyReg_Inst_ff_SDE_115_next_state}), .Q ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, new_AGEMA_signal_4705, RoundKey[115]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_116_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14016, new_AGEMA_signal_14015, new_AGEMA_signal_14014, KeyReg_Inst_ff_SDE_116_next_state}), .Q ({new_AGEMA_signal_4716, new_AGEMA_signal_4715, new_AGEMA_signal_4714, RoundKey[116]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_117_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14022, new_AGEMA_signal_14021, new_AGEMA_signal_14020, KeyReg_Inst_ff_SDE_117_next_state}), .Q ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, new_AGEMA_signal_4723, RoundKey[117]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_118_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14028, new_AGEMA_signal_14027, new_AGEMA_signal_14026, KeyReg_Inst_ff_SDE_118_next_state}), .Q ({new_AGEMA_signal_4734, new_AGEMA_signal_4733, new_AGEMA_signal_4732, RoundKey[118]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_119_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14034, new_AGEMA_signal_14033, new_AGEMA_signal_14032, KeyReg_Inst_ff_SDE_119_next_state}), .Q ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, new_AGEMA_signal_4741, RoundKey[119]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_120_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14040, new_AGEMA_signal_14039, new_AGEMA_signal_14038, KeyReg_Inst_ff_SDE_120_next_state}), .Q ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, new_AGEMA_signal_4759, RoundKey[120]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_121_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14676, new_AGEMA_signal_14675, new_AGEMA_signal_14674, KeyReg_Inst_ff_SDE_121_next_state}), .Q ({new_AGEMA_signal_4770, new_AGEMA_signal_4769, new_AGEMA_signal_4768, RoundKey[121]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_122_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14682, new_AGEMA_signal_14681, new_AGEMA_signal_14680, KeyReg_Inst_ff_SDE_122_next_state}), .Q ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, new_AGEMA_signal_4777, RoundKey[122]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_123_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14688, new_AGEMA_signal_14687, new_AGEMA_signal_14686, KeyReg_Inst_ff_SDE_123_next_state}), .Q ({new_AGEMA_signal_4788, new_AGEMA_signal_4787, new_AGEMA_signal_4786, RoundKey[123]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_124_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14694, new_AGEMA_signal_14693, new_AGEMA_signal_14692, KeyReg_Inst_ff_SDE_124_next_state}), .Q ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, new_AGEMA_signal_4795, RoundKey[124]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_125_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14700, new_AGEMA_signal_14699, new_AGEMA_signal_14698, KeyReg_Inst_ff_SDE_125_next_state}), .Q ({new_AGEMA_signal_4806, new_AGEMA_signal_4805, new_AGEMA_signal_4804, RoundKey[125]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_126_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14706, new_AGEMA_signal_14705, new_AGEMA_signal_14704, KeyReg_Inst_ff_SDE_126_next_state}), .Q ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, new_AGEMA_signal_4813, RoundKey[126]}) ) ;
    reg_masked #(.security_order(3), .pipeline(0)) KeyReg_Inst_ff_SDE_127_current_state_reg_FF_FF ( .clk (clk_gated), .D ({new_AGEMA_signal_14712, new_AGEMA_signal_14711, new_AGEMA_signal_14710, KeyReg_Inst_ff_SDE_127_next_state}), .Q ({new_AGEMA_signal_4824, new_AGEMA_signal_4823, new_AGEMA_signal_4822, RoundKey[127]}) ) ;
    DFF_X1 RoundCounterIns_count_reg_0__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N7), .Q (RoundCounter[0]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_1__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N8), .Q (RoundCounter[1]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_2__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_n1), .Q (RoundCounter[2]), .QN () ) ;
    DFF_X1 RoundCounterIns_count_reg_3__FF_FF ( .CK (clk_gated), .D (RoundCounterIns_N10), .Q (RoundCounter[3]), .QN () ) ;
endmodule
