module Reg1(x, y);
 input [135:0] x;
 output [134:0] y;

  assign y[0] = x[135];
  register_stage #(.WIDTH(134)) inst_0(.clk(x[134]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[17],x[28],x[39],x[50],x[61],x[66],x[67],x[68],x[69],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[62],x[63],x[64],x[65],x[70],x[81],x[92],x[103],x[114],x[125],x[130],x[131],x[132],x[133],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[126],x[127],x[128],x[129]}), .Q({y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134]}));
endmodule

module Reg2(x, y);
 input [273:0] x;
 output [272:0] y;

  assign y[0] = x[267];
  assign y[1] = x[268];
  assign y[2] = x[269];
  assign y[3] = x[270];
  assign y[4] = x[271];
  assign y[5] = x[272];
  assign y[6] = x[273];
  register_stage #(.WIDTH(266)) inst_0(.clk(x[266]), .D({x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[259],x[260],x[261],x[262],x[263],x[264],x[265],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[205],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258]}), .Q({y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265],y[266],y[267],y[268],y[269],y[270],y[271],y[272]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx5(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx6(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx12(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx13(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx19(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx20(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx26(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx27(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx33(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx34(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx40(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx41(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx47(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx48(x, y);
 input x;
 output y;

 wire t;
  assign t = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign y = t ^ x;
endmodule

module Fx49(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx50(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx51(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx52(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx53(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx54(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx55(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx56(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx57(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx58(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx59(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx60(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx61(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx62(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx63(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx64(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx65(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx66(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx67(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx68(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx69(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx70(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx71(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx72(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx73(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx74(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx75(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx76(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx77(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx78(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx79(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx80(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx81(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx82(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx83(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx84(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx85(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx86(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx87(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx88(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx89(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx90(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx91(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx92(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx93(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx94(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx95(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx96(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx97(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx98(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx99(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx100(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx101(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx102(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx103(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx104(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx105(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx106(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx107(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx108(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx109(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx110(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx111(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx112(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx113(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx114(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx115(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx116(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx117(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx118(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx119(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx120(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx121(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx122(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx123(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx124(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx125(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx126(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx127(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx128(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx129(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx130(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx131(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx132(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx133(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx134(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx135(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx136(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx137(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx138(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx139(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx140(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx141(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx142(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx143(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx144(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx145(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx146(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx147(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx148(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx149(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx150(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx151(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx152(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx153(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx154(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx155(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx156(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx157(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx158(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx159(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx160(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx161(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx162(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx163(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx164(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx165(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx166(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx167(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx168(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx169(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx170(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx171(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx172(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx173(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx174(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx175(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx176(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx177(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx178(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx179(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx180(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx181(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx182(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx183(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx184(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx185(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx186(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx187(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx188(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx189(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx190(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx191(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx192(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx193(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx194(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx195(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx196(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx197(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx198(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx199(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx200(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx201(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx202(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx203(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx204(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx205(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx206(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx207(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx208(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx209(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx210(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx211(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx212(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx213(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx214(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx215(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx216(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx217(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx218(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx219(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx220(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx221(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx222(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx223(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx224(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx225(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx226(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx227(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx228(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx229(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx230(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx231(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx232(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx233(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx234(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx235(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx236(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx237(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx238(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx239(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx240(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx241(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx242(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx243(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx244(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx245(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx246(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx247(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx248(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx249(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx250(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx251(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx252(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx253(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx254(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx255(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx256(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx257(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx258(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx259(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx260(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx261(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx262(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx263(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx264(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx265(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx266(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx267(x, y);
 input [3:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2]) | (~x[0] & x[1] & ~x[2]) | (~x[0] & ~x[1] & x[2]) | (x[0] & x[1] & x[2]);
  assign y = t ^ x[3];
endmodule

module Fx268(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx269(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx270(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx271(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module Fx272(x, y);
 input [2:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1]) | (~x[0] & x[1]);
  assign y = t ^ x[2];
endmodule

module FX(x, y);
 input [407:0] x;
 output [272:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[3], x[0]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[4], x[0]}), .y(y[3]));
  Fx4 Fx4_inst(.x(x[5]), .y(y[4]));
  Fx5 Fx5_inst(.x(x[6]), .y(y[5]));
  Fx6 Fx6_inst(.x(x[7]), .y(y[6]));
  Fx7 Fx7_inst(.x({x[9], x[8]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[10], x[8]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[11], x[8]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[12], x[8]}), .y(y[10]));
  Fx11 Fx11_inst(.x(x[13]), .y(y[11]));
  Fx12 Fx12_inst(.x(x[14]), .y(y[12]));
  Fx13 Fx13_inst(.x(x[15]), .y(y[13]));
  Fx14 Fx14_inst(.x({x[17], x[16]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[18], x[16]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[19], x[16]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[20], x[16]}), .y(y[17]));
  Fx18 Fx18_inst(.x(x[21]), .y(y[18]));
  Fx19 Fx19_inst(.x(x[22]), .y(y[19]));
  Fx20 Fx20_inst(.x(x[23]), .y(y[20]));
  Fx21 Fx21_inst(.x({x[25], x[24]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[26], x[24]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[27], x[24]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[28], x[24]}), .y(y[24]));
  Fx25 Fx25_inst(.x(x[29]), .y(y[25]));
  Fx26 Fx26_inst(.x(x[30]), .y(y[26]));
  Fx27 Fx27_inst(.x(x[31]), .y(y[27]));
  Fx28 Fx28_inst(.x({x[33], x[32]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[34], x[32]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[35], x[32]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[36], x[32]}), .y(y[31]));
  Fx32 Fx32_inst(.x(x[37]), .y(y[32]));
  Fx33 Fx33_inst(.x(x[38]), .y(y[33]));
  Fx34 Fx34_inst(.x(x[39]), .y(y[34]));
  Fx35 Fx35_inst(.x({x[41], x[40]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[42], x[40]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[43], x[40]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[44], x[40]}), .y(y[38]));
  Fx39 Fx39_inst(.x(x[45]), .y(y[39]));
  Fx40 Fx40_inst(.x(x[46]), .y(y[40]));
  Fx41 Fx41_inst(.x(x[47]), .y(y[41]));
  Fx42 Fx42_inst(.x({x[49], x[48]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[50], x[48]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[51], x[48]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[52], x[48]}), .y(y[45]));
  Fx46 Fx46_inst(.x(x[53]), .y(y[46]));
  Fx47 Fx47_inst(.x(x[54]), .y(y[47]));
  Fx48 Fx48_inst(.x(x[55]), .y(y[48]));
  Fx49 Fx49_inst(.x({x[59], x[58], x[57], x[56]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[61], x[60], x[57], x[56]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[62], x[58], x[56]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[63], x[60], x[56]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[64], x[58], x[57]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[65], x[60], x[57]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[66], x[60], x[58]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[70], x[69], x[68], x[67]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[72], x[71], x[68], x[67]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[73], x[69], x[67]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[74], x[71], x[67]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[75], x[69], x[68]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[76], x[71], x[68]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[77], x[71], x[69]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[81], x[80], x[79], x[78]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[83], x[82], x[79], x[78]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[84], x[80], x[78]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[85], x[82], x[78]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[86], x[80], x[79]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[87], x[82], x[79]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[88], x[82], x[80]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[92], x[91], x[90], x[89]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[94], x[93], x[90], x[89]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[95], x[91], x[89]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[96], x[93], x[89]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[97], x[91], x[90]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[98], x[93], x[90]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[99], x[93], x[91]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[103], x[102], x[101], x[100]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[105], x[104], x[101], x[100]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[106], x[102], x[100]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[107], x[104], x[100]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[108], x[102], x[101]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[109], x[104], x[101]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[110], x[104], x[102]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[114], x[113], x[112], x[111]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[116], x[115], x[112], x[111]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[117], x[113], x[111]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[118], x[115], x[111]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[119], x[113], x[112]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[120], x[115], x[112]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[121], x[115], x[113]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[125], x[124], x[123], x[122]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[127], x[126], x[123], x[122]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[128], x[124], x[122]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[129], x[126], x[122]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[130], x[124], x[123]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[131], x[126], x[123]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[132], x[126], x[124]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[136], x[135], x[134], x[133]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[138], x[137], x[134], x[133]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[139], x[135], x[133]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[140], x[137], x[133]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[141], x[135], x[134]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[142], x[137], x[134]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[143], x[137], x[135]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[147], x[146], x[145], x[144]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[149], x[148], x[145], x[144]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[150], x[146], x[144]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[151], x[148], x[144]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[152], x[146], x[145]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[153], x[148], x[145]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[154], x[148], x[146]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[158], x[157], x[156], x[155]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[160], x[159], x[156], x[155]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[161], x[157], x[155]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[162], x[159], x[155]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[163], x[157], x[156]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[164], x[159], x[156]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[165], x[159], x[157]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[169], x[168], x[167], x[166]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[171], x[170], x[167], x[166]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[172], x[168], x[166]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[173], x[170], x[166]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[174], x[168], x[167]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[175], x[170], x[167]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[176], x[170], x[168]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[180], x[179], x[178], x[177]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[182], x[181], x[178], x[177]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[183], x[179], x[177]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[184], x[181], x[177]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[185], x[179], x[178]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[186], x[181], x[178]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[187], x[181], x[179]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[191], x[190], x[189], x[188]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[193], x[192], x[189], x[188]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[194], x[190], x[188]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[195], x[192], x[188]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[196], x[190], x[189]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[197], x[192], x[189]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[198], x[192], x[190]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[202], x[201], x[200], x[199]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[204], x[203], x[200], x[199]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[205], x[201], x[199]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[206], x[203], x[199]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[207], x[201], x[200]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[208], x[203], x[200]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[209], x[203], x[201]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[213], x[212], x[211], x[210]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[215], x[214], x[211], x[210]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[216], x[212], x[210]}), .y(y[149]));
  Fx150 Fx150_inst(.x({x[217], x[214], x[210]}), .y(y[150]));
  Fx151 Fx151_inst(.x({x[218], x[212], x[211]}), .y(y[151]));
  Fx152 Fx152_inst(.x({x[219], x[214], x[211]}), .y(y[152]));
  Fx153 Fx153_inst(.x({x[220], x[214], x[212]}), .y(y[153]));
  Fx154 Fx154_inst(.x({x[224], x[223], x[222], x[221]}), .y(y[154]));
  Fx155 Fx155_inst(.x({x[226], x[225], x[222], x[221]}), .y(y[155]));
  Fx156 Fx156_inst(.x({x[227], x[223], x[221]}), .y(y[156]));
  Fx157 Fx157_inst(.x({x[228], x[225], x[221]}), .y(y[157]));
  Fx158 Fx158_inst(.x({x[229], x[223], x[222]}), .y(y[158]));
  Fx159 Fx159_inst(.x({x[230], x[225], x[222]}), .y(y[159]));
  Fx160 Fx160_inst(.x({x[231], x[225], x[223]}), .y(y[160]));
  Fx161 Fx161_inst(.x({x[235], x[234], x[233], x[232]}), .y(y[161]));
  Fx162 Fx162_inst(.x({x[237], x[236], x[233], x[232]}), .y(y[162]));
  Fx163 Fx163_inst(.x({x[238], x[234], x[232]}), .y(y[163]));
  Fx164 Fx164_inst(.x({x[239], x[236], x[232]}), .y(y[164]));
  Fx165 Fx165_inst(.x({x[240], x[234], x[233]}), .y(y[165]));
  Fx166 Fx166_inst(.x({x[241], x[236], x[233]}), .y(y[166]));
  Fx167 Fx167_inst(.x({x[242], x[236], x[234]}), .y(y[167]));
  Fx168 Fx168_inst(.x({x[246], x[245], x[244], x[243]}), .y(y[168]));
  Fx169 Fx169_inst(.x({x[248], x[247], x[244], x[243]}), .y(y[169]));
  Fx170 Fx170_inst(.x({x[249], x[245], x[243]}), .y(y[170]));
  Fx171 Fx171_inst(.x({x[250], x[247], x[243]}), .y(y[171]));
  Fx172 Fx172_inst(.x({x[251], x[245], x[244]}), .y(y[172]));
  Fx173 Fx173_inst(.x({x[252], x[247], x[244]}), .y(y[173]));
  Fx174 Fx174_inst(.x({x[253], x[247], x[245]}), .y(y[174]));
  Fx175 Fx175_inst(.x({x[257], x[256], x[255], x[254]}), .y(y[175]));
  Fx176 Fx176_inst(.x({x[259], x[258], x[255], x[254]}), .y(y[176]));
  Fx177 Fx177_inst(.x({x[260], x[256], x[254]}), .y(y[177]));
  Fx178 Fx178_inst(.x({x[261], x[258], x[254]}), .y(y[178]));
  Fx179 Fx179_inst(.x({x[262], x[256], x[255]}), .y(y[179]));
  Fx180 Fx180_inst(.x({x[263], x[258], x[255]}), .y(y[180]));
  Fx181 Fx181_inst(.x({x[264], x[258], x[256]}), .y(y[181]));
  Fx182 Fx182_inst(.x({x[268], x[267], x[266], x[265]}), .y(y[182]));
  Fx183 Fx183_inst(.x({x[270], x[269], x[266], x[265]}), .y(y[183]));
  Fx184 Fx184_inst(.x({x[271], x[267], x[265]}), .y(y[184]));
  Fx185 Fx185_inst(.x({x[272], x[269], x[265]}), .y(y[185]));
  Fx186 Fx186_inst(.x({x[273], x[267], x[266]}), .y(y[186]));
  Fx187 Fx187_inst(.x({x[274], x[269], x[266]}), .y(y[187]));
  Fx188 Fx188_inst(.x({x[275], x[269], x[267]}), .y(y[188]));
  Fx189 Fx189_inst(.x({x[279], x[278], x[277], x[276]}), .y(y[189]));
  Fx190 Fx190_inst(.x({x[281], x[280], x[277], x[276]}), .y(y[190]));
  Fx191 Fx191_inst(.x({x[282], x[278], x[276]}), .y(y[191]));
  Fx192 Fx192_inst(.x({x[283], x[280], x[276]}), .y(y[192]));
  Fx193 Fx193_inst(.x({x[284], x[278], x[277]}), .y(y[193]));
  Fx194 Fx194_inst(.x({x[285], x[280], x[277]}), .y(y[194]));
  Fx195 Fx195_inst(.x({x[286], x[280], x[278]}), .y(y[195]));
  Fx196 Fx196_inst(.x({x[290], x[289], x[288], x[287]}), .y(y[196]));
  Fx197 Fx197_inst(.x({x[292], x[291], x[288], x[287]}), .y(y[197]));
  Fx198 Fx198_inst(.x({x[293], x[289], x[287]}), .y(y[198]));
  Fx199 Fx199_inst(.x({x[294], x[291], x[287]}), .y(y[199]));
  Fx200 Fx200_inst(.x({x[295], x[289], x[288]}), .y(y[200]));
  Fx201 Fx201_inst(.x({x[296], x[291], x[288]}), .y(y[201]));
  Fx202 Fx202_inst(.x({x[297], x[291], x[289]}), .y(y[202]));
  Fx203 Fx203_inst(.x({x[301], x[300], x[299], x[298]}), .y(y[203]));
  Fx204 Fx204_inst(.x({x[303], x[302], x[299], x[298]}), .y(y[204]));
  Fx205 Fx205_inst(.x({x[304], x[300], x[298]}), .y(y[205]));
  Fx206 Fx206_inst(.x({x[305], x[302], x[298]}), .y(y[206]));
  Fx207 Fx207_inst(.x({x[306], x[300], x[299]}), .y(y[207]));
  Fx208 Fx208_inst(.x({x[307], x[302], x[299]}), .y(y[208]));
  Fx209 Fx209_inst(.x({x[308], x[302], x[300]}), .y(y[209]));
  Fx210 Fx210_inst(.x({x[312], x[311], x[310], x[309]}), .y(y[210]));
  Fx211 Fx211_inst(.x({x[314], x[313], x[310], x[309]}), .y(y[211]));
  Fx212 Fx212_inst(.x({x[315], x[311], x[309]}), .y(y[212]));
  Fx213 Fx213_inst(.x({x[316], x[313], x[309]}), .y(y[213]));
  Fx214 Fx214_inst(.x({x[317], x[311], x[310]}), .y(y[214]));
  Fx215 Fx215_inst(.x({x[318], x[313], x[310]}), .y(y[215]));
  Fx216 Fx216_inst(.x({x[319], x[313], x[311]}), .y(y[216]));
  Fx217 Fx217_inst(.x({x[323], x[322], x[321], x[320]}), .y(y[217]));
  Fx218 Fx218_inst(.x({x[325], x[324], x[321], x[320]}), .y(y[218]));
  Fx219 Fx219_inst(.x({x[326], x[322], x[320]}), .y(y[219]));
  Fx220 Fx220_inst(.x({x[327], x[324], x[320]}), .y(y[220]));
  Fx221 Fx221_inst(.x({x[328], x[322], x[321]}), .y(y[221]));
  Fx222 Fx222_inst(.x({x[329], x[324], x[321]}), .y(y[222]));
  Fx223 Fx223_inst(.x({x[330], x[324], x[322]}), .y(y[223]));
  Fx224 Fx224_inst(.x({x[334], x[333], x[332], x[331]}), .y(y[224]));
  Fx225 Fx225_inst(.x({x[336], x[335], x[332], x[331]}), .y(y[225]));
  Fx226 Fx226_inst(.x({x[337], x[333], x[331]}), .y(y[226]));
  Fx227 Fx227_inst(.x({x[338], x[335], x[331]}), .y(y[227]));
  Fx228 Fx228_inst(.x({x[339], x[333], x[332]}), .y(y[228]));
  Fx229 Fx229_inst(.x({x[340], x[335], x[332]}), .y(y[229]));
  Fx230 Fx230_inst(.x({x[341], x[335], x[333]}), .y(y[230]));
  Fx231 Fx231_inst(.x({x[345], x[344], x[343], x[342]}), .y(y[231]));
  Fx232 Fx232_inst(.x({x[347], x[346], x[343], x[342]}), .y(y[232]));
  Fx233 Fx233_inst(.x({x[348], x[344], x[342]}), .y(y[233]));
  Fx234 Fx234_inst(.x({x[349], x[346], x[342]}), .y(y[234]));
  Fx235 Fx235_inst(.x({x[350], x[344], x[343]}), .y(y[235]));
  Fx236 Fx236_inst(.x({x[351], x[346], x[343]}), .y(y[236]));
  Fx237 Fx237_inst(.x({x[352], x[346], x[344]}), .y(y[237]));
  Fx238 Fx238_inst(.x({x[356], x[355], x[354], x[353]}), .y(y[238]));
  Fx239 Fx239_inst(.x({x[358], x[357], x[354], x[353]}), .y(y[239]));
  Fx240 Fx240_inst(.x({x[359], x[355], x[353]}), .y(y[240]));
  Fx241 Fx241_inst(.x({x[360], x[357], x[353]}), .y(y[241]));
  Fx242 Fx242_inst(.x({x[361], x[355], x[354]}), .y(y[242]));
  Fx243 Fx243_inst(.x({x[362], x[357], x[354]}), .y(y[243]));
  Fx244 Fx244_inst(.x({x[363], x[357], x[355]}), .y(y[244]));
  Fx245 Fx245_inst(.x({x[367], x[366], x[365], x[364]}), .y(y[245]));
  Fx246 Fx246_inst(.x({x[369], x[368], x[365], x[364]}), .y(y[246]));
  Fx247 Fx247_inst(.x({x[370], x[366], x[364]}), .y(y[247]));
  Fx248 Fx248_inst(.x({x[371], x[368], x[364]}), .y(y[248]));
  Fx249 Fx249_inst(.x({x[372], x[366], x[365]}), .y(y[249]));
  Fx250 Fx250_inst(.x({x[373], x[368], x[365]}), .y(y[250]));
  Fx251 Fx251_inst(.x({x[374], x[368], x[366]}), .y(y[251]));
  Fx252 Fx252_inst(.x({x[378], x[377], x[376], x[375]}), .y(y[252]));
  Fx253 Fx253_inst(.x({x[380], x[379], x[376], x[375]}), .y(y[253]));
  Fx254 Fx254_inst(.x({x[381], x[377], x[375]}), .y(y[254]));
  Fx255 Fx255_inst(.x({x[382], x[379], x[375]}), .y(y[255]));
  Fx256 Fx256_inst(.x({x[383], x[377], x[376]}), .y(y[256]));
  Fx257 Fx257_inst(.x({x[384], x[379], x[376]}), .y(y[257]));
  Fx258 Fx258_inst(.x({x[385], x[379], x[377]}), .y(y[258]));
  Fx259 Fx259_inst(.x({x[389], x[388], x[387], x[386]}), .y(y[259]));
  Fx260 Fx260_inst(.x({x[391], x[390], x[387], x[386]}), .y(y[260]));
  Fx261 Fx261_inst(.x({x[392], x[388], x[386]}), .y(y[261]));
  Fx262 Fx262_inst(.x({x[393], x[390], x[386]}), .y(y[262]));
  Fx263 Fx263_inst(.x({x[394], x[388], x[387]}), .y(y[263]));
  Fx264 Fx264_inst(.x({x[395], x[390], x[387]}), .y(y[264]));
  Fx265 Fx265_inst(.x({x[396], x[390], x[388]}), .y(y[265]));
  Fx266 Fx266_inst(.x({x[400], x[399], x[398], x[397]}), .y(y[266]));
  Fx267 Fx267_inst(.x({x[402], x[401], x[398], x[397]}), .y(y[267]));
  Fx268 Fx268_inst(.x({x[403], x[399], x[397]}), .y(y[268]));
  Fx269 Fx269_inst(.x({x[404], x[401], x[397]}), .y(y[269]));
  Fx270 Fx270_inst(.x({x[405], x[399], x[398]}), .y(y[270]));
  Fx271 Fx271_inst(.x({x[406], x[401], x[398]}), .y(y[271]));
  Fx272 Fx272_inst(.x({x[407], x[401], x[399]}), .y(y[272]));
endmodule

module R1ind0(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[1] & ~x[3] & x[4] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[0] & x[1] & ~x[2] & x[5] & ~x[6]) | (x[0] & ~x[3] & x[4] & x[5] & ~x[6]) | (x[0] & ~x[2] & x[3] & x[4]) | (x[1] & x[2] & ~x[3] & x[5]) | (x[1] & ~x[3] & x[4] & x[5]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[0] & x[2] & ~x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[3] & ~x[5] & x[6]) | (x[0] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[1] & x[2] & ~x[3] & x[6]) | (x[1] & x[4] & ~x[5] & x[6]) | (x[2] & x[4] & x[6]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [7:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[1] = (x[1] & ~x[2] & x[3] & ~x[4] & x[5]) | (x[1] & ~x[2] & x[3] & ~x[4] & x[6]) | (x[1] & ~x[2] & ~x[4] & x[5] & x[6]) | (x[0] & x[2] & x[3] & x[4] & x[5]) | (x[0] & ~x[2] & x[3] & x[6]) | (x[0] & ~x[4] & x[5] & x[6]) | (x[3] & x[5] & x[6]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [47:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[16] ^ x[47];
  assign t[11] = (x[0] & x[1] & x[2] & ~x[5] & ~x[6]) | (x[0] & x[1] & x[3] & ~x[4] & ~x[6]) | (x[0] & x[2] & x[3] & ~x[5] & ~x[6]) | (~x[1] & x[2] & x[3] & x[4] & ~x[6]) | (x[1] & x[2] & x[3] & ~x[5]) | (x[1] & x[3] & x[4] & ~x[5]) | (x[0] & x[2] & ~x[4] & x[5]);
  assign t[12] = (x[8] & x[9] & x[10] & ~x[13] & ~x[14]) | (x[8] & x[9] & x[11] & ~x[12] & ~x[14]) | (x[8] & x[10] & x[11] & ~x[13] & ~x[14]) | (~x[9] & x[10] & x[11] & x[12] & ~x[14]) | (x[9] & x[10] & x[11] & ~x[13]) | (x[9] & x[11] & x[12] & ~x[13]) | (x[8] & x[10] & ~x[12] & x[13]);
  assign t[13] = (x[16] & x[17] & x[18] & ~x[21] & ~x[22]) | (x[16] & x[17] & x[19] & ~x[20] & ~x[22]) | (x[16] & x[18] & x[19] & ~x[21] & ~x[22]) | (~x[17] & x[18] & x[19] & x[20] & ~x[22]) | (x[17] & x[18] & x[19] & ~x[21]) | (x[17] & x[19] & x[20] & ~x[21]) | (x[16] & x[18] & ~x[20] & x[21]);
  assign t[14] = (x[24] & x[25] & x[26] & ~x[29] & ~x[30]) | (x[24] & x[25] & x[27] & ~x[28] & ~x[30]) | (x[24] & x[26] & x[27] & ~x[29] & ~x[30]) | (~x[25] & x[26] & x[27] & x[28] & ~x[30]) | (x[25] & x[26] & x[27] & ~x[29]) | (x[25] & x[27] & x[28] & ~x[29]) | (x[24] & x[26] & ~x[28] & x[29]);
  assign t[15] = (x[32] & x[33] & x[34] & ~x[37] & ~x[38]) | (x[32] & x[33] & x[35] & ~x[36] & ~x[38]) | (x[32] & x[34] & x[35] & ~x[37] & ~x[38]) | (~x[33] & x[34] & x[35] & x[36] & ~x[38]) | (x[33] & x[34] & x[35] & ~x[37]) | (x[33] & x[35] & x[36] & ~x[37]) | (x[32] & x[34] & ~x[36] & x[37]);
  assign t[16] = (x[40] & x[41] & x[42] & ~x[45] & ~x[46]) | (x[40] & x[41] & x[43] & ~x[44] & ~x[46]) | (x[40] & x[42] & x[43] & ~x[45] & ~x[46]) | (~x[41] & x[42] & x[43] & x[44] & ~x[46]) | (x[41] & x[42] & x[43] & ~x[45]) | (x[41] & x[43] & x[44] & ~x[45]) | (x[40] & x[42] & ~x[44] & x[45]);
  assign t[1] = ~(t[5] & t[6]);
  assign t[2] = ~(t[7] | t[8]);
  assign t[3] = ~(t[9] | t[4]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[15];
  assign t[7] = t[13] ^ x[23];
  assign t[8] = t[14] ^ x[31];
  assign t[9] = t[15] ^ x[39];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind66(x, y);
 input [48:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] ? t[6] : t[1];
  assign t[10] = t[16] ^ x[48];
  assign t[11] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[12] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign t[13] = (x[17] & x[18] & x[19] & ~x[22] & ~x[23]) | (x[17] & x[18] & x[20] & ~x[21] & ~x[23]) | (x[17] & x[19] & x[20] & ~x[22] & ~x[23]) | (~x[18] & x[19] & x[20] & x[21] & ~x[23]) | (x[18] & x[19] & x[20] & ~x[22]) | (x[18] & x[20] & x[21] & ~x[22]) | (x[17] & x[19] & ~x[21] & x[22]);
  assign t[14] = (x[25] & x[26] & x[27] & ~x[30] & ~x[31]) | (x[25] & x[26] & x[28] & ~x[29] & ~x[31]) | (x[25] & x[27] & x[28] & ~x[30] & ~x[31]) | (~x[26] & x[27] & x[28] & x[29] & ~x[31]) | (x[26] & x[27] & x[28] & ~x[30]) | (x[26] & x[28] & x[29] & ~x[30]) | (x[25] & x[27] & ~x[29] & x[30]);
  assign t[15] = (x[33] & x[34] & x[35] & ~x[38] & ~x[39]) | (x[33] & x[34] & x[36] & ~x[37] & ~x[39]) | (x[33] & x[35] & x[36] & ~x[38] & ~x[39]) | (~x[34] & x[35] & x[36] & x[37] & ~x[39]) | (x[34] & x[35] & x[36] & ~x[38]) | (x[34] & x[36] & x[37] & ~x[38]) | (x[33] & x[35] & ~x[37] & x[38]);
  assign t[16] = (x[41] & x[42] & x[43] & ~x[46] & ~x[47]) | (x[41] & x[42] & x[44] & ~x[45] & ~x[47]) | (x[41] & x[43] & x[44] & ~x[46] & ~x[47]) | (~x[42] & x[43] & x[44] & x[45] & ~x[47]) | (x[42] & x[43] & x[44] & ~x[46]) | (x[42] & x[44] & x[45] & ~x[46]) | (x[41] & x[43] & ~x[45] & x[46]);
  assign t[1] = ~(t[6] & t[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = t[7] & t[8];
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[8];
  assign t[6] = t[12] ^ x[16];
  assign t[7] = t[13] ^ x[24];
  assign t[8] = t[14] ^ x[32];
  assign t[9] = t[15] ^ x[40];
  assign y = ~(~x[0] & ~t[0]);
endmodule

module R1ind67(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind68(x, y);
 input [48:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[1] & t[5];
  assign t[10] = t[16] ^ x[48];
  assign t[11] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[12] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign t[13] = (x[17] & x[18] & x[19] & ~x[22] & ~x[23]) | (x[17] & x[18] & x[20] & ~x[21] & ~x[23]) | (x[17] & x[19] & x[20] & ~x[22] & ~x[23]) | (~x[18] & x[19] & x[20] & x[21] & ~x[23]) | (x[18] & x[19] & x[20] & ~x[22]) | (x[18] & x[20] & x[21] & ~x[22]) | (x[17] & x[19] & ~x[21] & x[22]);
  assign t[14] = (x[25] & x[26] & x[27] & ~x[30] & ~x[31]) | (x[25] & x[26] & x[28] & ~x[29] & ~x[31]) | (x[25] & x[27] & x[28] & ~x[30] & ~x[31]) | (~x[26] & x[27] & x[28] & x[29] & ~x[31]) | (x[26] & x[27] & x[28] & ~x[30]) | (x[26] & x[28] & x[29] & ~x[30]) | (x[25] & x[27] & ~x[29] & x[30]);
  assign t[15] = (x[33] & x[34] & x[35] & ~x[38] & ~x[39]) | (x[33] & x[34] & x[36] & ~x[37] & ~x[39]) | (x[33] & x[35] & x[36] & ~x[38] & ~x[39]) | (~x[34] & x[35] & x[36] & x[37] & ~x[39]) | (x[34] & x[35] & x[36] & ~x[38]) | (x[34] & x[36] & x[37] & ~x[38]) | (x[33] & x[35] & ~x[37] & x[38]);
  assign t[16] = (x[41] & x[42] & x[43] & ~x[46] & ~x[47]) | (x[41] & x[42] & x[44] & ~x[45] & ~x[47]) | (x[41] & x[43] & x[44] & ~x[46] & ~x[47]) | (~x[42] & x[43] & x[44] & x[45] & ~x[47]) | (x[42] & x[43] & x[44] & ~x[46]) | (x[42] & x[44] & x[45] & ~x[46]) | (x[41] & x[43] & ~x[45] & x[46]);
  assign t[1] = ~(t[2] & t[6]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[3] = ~(t[8] & t[4]);
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[8];
  assign t[6] = t[12] ^ x[16];
  assign t[7] = t[13] ^ x[24];
  assign t[8] = t[14] ^ x[32];
  assign t[9] = t[15] ^ x[40];
  assign y = ~x[0] & t[0];
endmodule

module R1ind69(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind70(x, y);
 input [8:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = ~x[0] & t[0];
endmodule

module R1ind71(x, y);
 input [48:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[5] | t[1];
  assign t[10] = t[16] ^ x[48];
  assign t[11] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign t[12] = (x[9] & x[10] & x[11] & ~x[14] & ~x[15]) | (x[9] & x[10] & x[12] & ~x[13] & ~x[15]) | (x[9] & x[11] & x[12] & ~x[14] & ~x[15]) | (~x[10] & x[11] & x[12] & x[13] & ~x[15]) | (x[10] & x[11] & x[12] & ~x[14]) | (x[10] & x[12] & x[13] & ~x[14]) | (x[9] & x[11] & ~x[13] & x[14]);
  assign t[13] = (x[17] & x[18] & x[19] & ~x[22] & ~x[23]) | (x[17] & x[18] & x[20] & ~x[21] & ~x[23]) | (x[17] & x[19] & x[20] & ~x[22] & ~x[23]) | (~x[18] & x[19] & x[20] & x[21] & ~x[23]) | (x[18] & x[19] & x[20] & ~x[22]) | (x[18] & x[20] & x[21] & ~x[22]) | (x[17] & x[19] & ~x[21] & x[22]);
  assign t[14] = (x[25] & x[26] & x[27] & ~x[30] & ~x[31]) | (x[25] & x[26] & x[28] & ~x[29] & ~x[31]) | (x[25] & x[27] & x[28] & ~x[30] & ~x[31]) | (~x[26] & x[27] & x[28] & x[29] & ~x[31]) | (x[26] & x[27] & x[28] & ~x[30]) | (x[26] & x[28] & x[29] & ~x[30]) | (x[25] & x[27] & ~x[29] & x[30]);
  assign t[15] = (x[33] & x[34] & x[35] & ~x[38] & ~x[39]) | (x[33] & x[34] & x[36] & ~x[37] & ~x[39]) | (x[33] & x[35] & x[36] & ~x[38] & ~x[39]) | (~x[34] & x[35] & x[36] & x[37] & ~x[39]) | (x[34] & x[35] & x[36] & ~x[38]) | (x[34] & x[36] & x[37] & ~x[38]) | (x[33] & x[35] & ~x[37] & x[38]);
  assign t[16] = (x[41] & x[42] & x[43] & ~x[46] & ~x[47]) | (x[41] & x[42] & x[44] & ~x[45] & ~x[47]) | (x[41] & x[43] & x[44] & ~x[46] & ~x[47]) | (~x[42] & x[43] & x[44] & x[45] & ~x[47]) | (x[42] & x[43] & x[44] & ~x[46]) | (x[42] & x[44] & x[45] & ~x[46]) | (x[41] & x[43] & ~x[45] & x[46]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[3] = ~(t[8] | t[4]);
  assign t[4] = ~(t[9] & t[10]);
  assign t[5] = t[11] ^ x[8];
  assign t[6] = t[12] ^ x[16];
  assign t[7] = t[13] ^ x[24];
  assign t[8] = t[14] ^ x[32];
  assign t[9] = t[15] ^ x[40];
  assign y = ~x[0] & t[0];
endmodule

module R1ind72(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind73(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind74(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind75(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind76(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind77(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind78(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind79(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind80(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind81(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind82(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind83(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind84(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind85(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind86(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind87(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind88(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind89(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind90(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind91(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind92(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind93(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind94(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind95(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind96(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind97(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind98(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind99(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind100(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind101(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind102(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind103(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind104(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind105(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind106(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind107(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind108(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind109(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind110(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind111(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind112(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind113(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind114(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind115(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind116(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind117(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind118(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind119(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind120(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind121(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind122(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind123(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind124(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind125(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind126(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind127(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind128(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind129(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind130(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind131(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind132(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & x[3] & ~x[6] & ~x[7]) | (x[1] & x[2] & x[4] & ~x[5] & ~x[7]) | (x[1] & x[3] & x[4] & ~x[6] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[2] & x[3] & x[4] & ~x[6]) | (x[2] & x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind133(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[2] & ~x[4] & x[5] & ~x[7]) | (~x[2] & x[3] & x[4] & x[5] & ~x[7]) | (x[1] & x[2] & ~x[3] & x[6] & ~x[7]) | (x[1] & ~x[4] & x[5] & x[6] & ~x[7]) | (x[1] & ~x[3] & x[4] & x[5]) | (x[2] & x[3] & ~x[4] & x[6]) | (x[2] & ~x[4] & x[5] & x[6]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind134(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[1] & x[3] & ~x[4] & x[5] & ~x[6]) | (x[1] & x[3] & ~x[4] & ~x[6] & x[7]) | (x[1] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[2] & x[3] & ~x[4] & x[7]) | (x[2] & x[5] & ~x[6] & x[7]) | (x[3] & x[5] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind135(x, y);
 input [9:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[8];
  assign t[1] = (x[2] & ~x[3] & x[4] & ~x[5] & x[6]) | (x[2] & ~x[3] & x[4] & ~x[5] & x[7]) | (x[2] & ~x[3] & ~x[5] & x[6] & x[7]) | (x[1] & x[3] & x[4] & x[5] & x[6]) | (x[1] & ~x[3] & x[4] & x[7]) | (x[1] & ~x[5] & x[6] & x[7]) | (x[4] & x[6] & x[7]);
  assign y = x[0] ? x[9] : t[0];
endmodule

module R1ind136(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[52] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind137(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[48] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind138(x, y);
 input [29:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[18];
  assign t[19] = t[26] ^ x[19];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[27];
  assign t[21] = t[28] ^ x[28];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[24] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[25] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[26] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[27] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[28] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[29] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind139(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[18];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[20];
  assign t[29] = t[38] ^ x[28];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[29];
  assign t[31] = t[40] ^ x[30];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[34] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[35] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[36] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[37] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[41] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind140(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[52] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind141(x, y);
 input [31:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[17] & t[18];
  assign t[11] = t[19] ^ t[10];
  assign t[12] = t[38] ^ t[17];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[39] ^ t[40];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[40]);
  assign t[18] = ~(t[38] ^ t[17]);
  assign t[19] = t[38] & t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[27];
  assign t[21] = t[28] & t[29];
  assign t[22] = t[30] ^ t[21];
  assign t[23] = t[41] ^ t[28];
  assign t[24] = t[38] ^ t[31];
  assign t[25] = t[32] ^ t[16];
  assign t[26] = t[42] ^ t[43];
  assign t[27] = t[28] & t[33];
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[41] ^ t[28]);
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] & t[34];
  assign t[31] = t[40] ^ t[44];
  assign t[32] = t[38] ^ t[15];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[27];
  assign t[35] = t[43] ^ t[45];
  assign t[36] = t[41] ^ t[26];
  assign t[37] = t[46] ^ x[9];
  assign t[38] = t[47] ^ x[17];
  assign t[39] = t[48] ^ x[18];
  assign t[3] = ~(t[5] ^ t[37]);
  assign t[40] = t[49] ^ x[19];
  assign t[41] = t[50] ^ x[27];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[29];
  assign t[44] = t[53] ^ x[30];
  assign t[45] = t[54] ^ x[31];
  assign t[46] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[47] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[4] = ~(t[6] ^ t[7]);
  assign t[50] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[54] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[9] = t[15] ^ t[16];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind142(x, y);
 input [29:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[18];
  assign t[19] = t[26] ^ x[19];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[27];
  assign t[21] = t[28] ^ x[28];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[24] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[25] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[26] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[27] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[28] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[29] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind143(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[18];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[20];
  assign t[29] = t[38] ^ x[28];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[29];
  assign t[31] = t[40] ^ x[30];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[34] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[35] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[36] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[37] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[41] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind144(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[52] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind145(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[48] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind146(x, y);
 input [29:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[18];
  assign t[19] = t[26] ^ x[19];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[27];
  assign t[21] = t[28] ^ x[28];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[24] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[25] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[26] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[27] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[28] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[29] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind147(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[18];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[20];
  assign t[29] = t[38] ^ x[28];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[29];
  assign t[31] = t[40] ^ x[30];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[34] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[35] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[36] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[37] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[41] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind148(x, y);
 input [39:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[18] ^ t[19];
  assign t[13] = ~(t[41]);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[20] ^ t[9]);
  assign t[17] = ~t[21];
  assign t[18] = t[39] ^ t[15];
  assign t[19] = t[13] & t[20];
  assign t[1] = ~t[3];
  assign t[20] = t[39] ^ t[22];
  assign t[21] = t[23] ^ t[24];
  assign t[22] = t[41] ^ t[43];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] & t[28];
  assign t[25] = t[44] & t[29];
  assign t[26] = t[30] & t[31];
  assign t[27] = t[32] ^ t[30];
  assign t[28] = t[33] ^ t[26];
  assign t[29] = t[34] ^ t[35];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[44] ^ t[30]);
  assign t[32] = t[46] ^ t[45];
  assign t[33] = ~(t[36] ^ t[27]);
  assign t[34] = t[44] ^ t[32];
  assign t[35] = t[30] & t[36];
  assign t[36] = t[44] ^ t[37];
  assign t[37] = t[45] ^ t[47];
  assign t[38] = t[48] ^ x[9];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[25];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[27];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[37];
  assign t[46] = t[56] ^ x[38];
  assign t[47] = t[57] ^ x[39];
  assign t[48] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[49] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[51] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[52] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[53] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[54] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[55] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[56] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[57] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[39] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind149(x, y);
 input [39:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[39] ^ t[14];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[41] ^ t[42];
  assign t[13] = t[14] & t[18];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[39] ^ t[14]);
  assign t[16] = t[39] & t[19];
  assign t[17] = ~t[20];
  assign t[18] = t[39] ^ t[21];
  assign t[19] = t[22] ^ t[13];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] ^ t[24]);
  assign t[21] = t[42] ^ t[43];
  assign t[22] = t[39] ^ t[12];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[29] ^ t[30];
  assign t[26] = t[31] & t[32];
  assign t[27] = t[33] ^ t[26];
  assign t[28] = t[44] ^ t[31];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[31] & t[34];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[44] ^ t[31]);
  assign t[33] = t[44] & t[35];
  assign t[34] = t[44] ^ t[36];
  assign t[35] = t[37] ^ t[30];
  assign t[36] = t[46] ^ t[47];
  assign t[37] = t[44] ^ t[29];
  assign t[38] = t[48] ^ x[9];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[25];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[27];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[37];
  assign t[46] = t[56] ^ x[38];
  assign t[47] = t[57] ^ x[39];
  assign t[48] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[49] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[51] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[52] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[53] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[54] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[55] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[56] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[57] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind150(x, y);
 input [37:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[22] ^ t[9]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[15];
  assign t[14] = t[23] ^ t[24];
  assign t[15] = t[16] & t[17];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[25] ^ t[16]);
  assign t[18] = t[26] ^ x[9];
  assign t[19] = t[27] ^ x[17];
  assign t[1] = ~t[3];
  assign t[20] = t[28] ^ x[18];
  assign t[21] = t[29] ^ x[26];
  assign t[22] = t[30] ^ x[27];
  assign t[23] = t[31] ^ x[35];
  assign t[24] = t[32] ^ x[36];
  assign t[25] = t[33] ^ x[37];
  assign t[26] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[27] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[28] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[29] = (x[19] & x[20] & x[21] & ~x[24] & ~x[25]) | (x[19] & x[20] & x[22] & ~x[23] & ~x[25]) | (x[19] & x[21] & x[22] & ~x[24] & ~x[25]) | (~x[20] & x[21] & x[22] & x[23] & ~x[25]) | (x[20] & x[21] & x[22] & ~x[24]) | (x[20] & x[22] & x[23] & ~x[24]) | (x[19] & x[21] & ~x[23] & x[24]);
  assign t[2] = ~(t[4]);
  assign t[30] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[31] = (x[28] & x[30] & ~x[31] & x[32] & ~x[33]) | (x[28] & x[30] & ~x[31] & ~x[33] & x[34]) | (x[28] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[29] & x[30] & ~x[31] & x[34]) | (x[29] & x[32] & ~x[33] & x[34]) | (x[30] & x[32] & x[34]);
  assign t[32] = (x[29] & ~x[30] & x[31] & ~x[32] & x[33]) | (x[29] & ~x[30] & x[31] & ~x[32] & x[34]) | (x[29] & ~x[30] & ~x[32] & x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[28] & ~x[30] & x[31] & x[34]) | (x[28] & ~x[32] & x[33] & x[34]) | (x[31] & x[33] & x[34]);
  assign t[33] = (x[28] & x[29] & ~x[31] & x[32] & ~x[34]) | (~x[29] & x[30] & x[31] & x[32] & ~x[34]) | (x[28] & x[29] & ~x[30] & x[33] & ~x[34]) | (x[28] & ~x[31] & x[32] & x[33] & ~x[34]) | (x[28] & ~x[30] & x[31] & x[32]) | (x[29] & x[30] & ~x[31] & x[33]) | (x[29] & ~x[31] & x[32] & x[33]);
  assign t[3] = ~(t[5] ^ t[18]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[19] ^ t[20];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11] ^ t[21]);
  assign t[9] = ~(t[19]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind151(x, y);
 input [39:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[29]);
  assign t[12] = ~(t[30] ^ t[11]);
  assign t[13] = ~t[15];
  assign t[14] = t[30] ^ t[16];
  assign t[15] = ~(t[17]);
  assign t[16] = t[29] ^ t[31];
  assign t[17] = t[18] ^ t[19];
  assign t[18] = t[20] ^ t[21];
  assign t[19] = t[22] & t[23];
  assign t[1] = ~t[3];
  assign t[20] = t[32] ^ t[33];
  assign t[21] = t[22] & t[24];
  assign t[22] = ~(t[33]);
  assign t[23] = ~(t[34] ^ t[22]);
  assign t[24] = t[34] ^ t[25];
  assign t[25] = t[33] ^ t[35];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[17];
  assign t[28] = t[38] ^ x[25];
  assign t[29] = t[39] ^ x[26];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[27];
  assign t[31] = t[41] ^ x[28];
  assign t[32] = t[42] ^ x[36];
  assign t[33] = t[43] ^ x[37];
  assign t[34] = t[44] ^ x[38];
  assign t[35] = t[45] ^ x[39];
  assign t[36] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[37] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[38] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[39] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[3] = ~(t[5] ^ t[26]);
  assign t[40] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[41] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[42] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[43] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[44] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[45] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13] ^ t[27]);
  assign t[9] = t[28] ^ t[29];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind152(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[52] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind153(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[48] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind154(x, y);
 input [29:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[18];
  assign t[19] = t[26] ^ x[19];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[27];
  assign t[21] = t[28] ^ x[28];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[24] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[25] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[26] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[27] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[28] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[29] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind155(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[18];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[20];
  assign t[29] = t[38] ^ x[28];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[29];
  assign t[31] = t[40] ^ x[30];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[34] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[35] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[36] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[37] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[41] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind156(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[52] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind157(x, y);
 input [31:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[17] & t[18];
  assign t[11] = t[19] ^ t[10];
  assign t[12] = t[38] ^ t[17];
  assign t[13] = t[20] ^ t[21];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[39] ^ t[40];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[40]);
  assign t[18] = ~(t[38] ^ t[17]);
  assign t[19] = t[38] & t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[27];
  assign t[21] = t[28] & t[29];
  assign t[22] = t[30] ^ t[21];
  assign t[23] = t[41] ^ t[28];
  assign t[24] = t[38] ^ t[31];
  assign t[25] = t[32] ^ t[16];
  assign t[26] = t[42] ^ t[43];
  assign t[27] = t[28] & t[33];
  assign t[28] = ~(t[43]);
  assign t[29] = ~(t[41] ^ t[28]);
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] & t[34];
  assign t[31] = t[40] ^ t[44];
  assign t[32] = t[38] ^ t[15];
  assign t[33] = t[41] ^ t[35];
  assign t[34] = t[36] ^ t[27];
  assign t[35] = t[43] ^ t[45];
  assign t[36] = t[41] ^ t[26];
  assign t[37] = t[46] ^ x[9];
  assign t[38] = t[47] ^ x[17];
  assign t[39] = t[48] ^ x[18];
  assign t[3] = ~(t[5] ^ t[37]);
  assign t[40] = t[49] ^ x[19];
  assign t[41] = t[50] ^ x[27];
  assign t[42] = t[51] ^ x[28];
  assign t[43] = t[52] ^ x[29];
  assign t[44] = t[53] ^ x[30];
  assign t[45] = t[54] ^ x[31];
  assign t[46] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[47] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[4] = ~(t[6] ^ t[7]);
  assign t[50] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[54] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[9] = t[15] ^ t[16];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind158(x, y);
 input [29:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[18];
  assign t[19] = t[26] ^ x[19];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[27];
  assign t[21] = t[28] ^ x[28];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[24] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[25] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[26] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[27] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[28] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[29] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind159(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[18];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[20];
  assign t[29] = t[38] ^ x[28];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[29];
  assign t[31] = t[40] ^ x[30];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[34] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[35] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[36] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[37] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[41] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind160(x, y);
 input [39:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[18] ^ t[19];
  assign t[13] = ~(t[41]);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[20] ^ t[9]);
  assign t[17] = ~t[21];
  assign t[18] = t[39] ^ t[15];
  assign t[19] = t[13] & t[20];
  assign t[1] = ~t[3];
  assign t[20] = t[39] ^ t[22];
  assign t[21] = t[23] ^ t[24];
  assign t[22] = t[41] ^ t[43];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] & t[28];
  assign t[25] = t[44] & t[29];
  assign t[26] = t[30] & t[31];
  assign t[27] = t[32] ^ t[30];
  assign t[28] = t[33] ^ t[26];
  assign t[29] = t[34] ^ t[35];
  assign t[2] = t[4] ^ t[5];
  assign t[30] = ~(t[45]);
  assign t[31] = ~(t[44] ^ t[30]);
  assign t[32] = t[46] ^ t[45];
  assign t[33] = ~(t[36] ^ t[27]);
  assign t[34] = t[44] ^ t[32];
  assign t[35] = t[30] & t[36];
  assign t[36] = t[44] ^ t[37];
  assign t[37] = t[45] ^ t[47];
  assign t[38] = t[48] ^ x[9];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[25];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[27];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[37];
  assign t[46] = t[56] ^ x[38];
  assign t[47] = t[57] ^ x[39];
  assign t[48] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[49] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[51] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[52] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[53] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[54] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[55] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[56] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[57] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[39] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind161(x, y);
 input [39:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[39] ^ t[14];
  assign t[11] = ~(t[17] ^ t[40]);
  assign t[12] = t[41] ^ t[42];
  assign t[13] = t[14] & t[18];
  assign t[14] = ~(t[42]);
  assign t[15] = ~(t[39] ^ t[14]);
  assign t[16] = t[39] & t[19];
  assign t[17] = ~t[20];
  assign t[18] = t[39] ^ t[21];
  assign t[19] = t[22] ^ t[13];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[23] ^ t[24]);
  assign t[21] = t[42] ^ t[43];
  assign t[22] = t[39] ^ t[12];
  assign t[23] = t[25] ^ t[26];
  assign t[24] = t[27] ^ t[28];
  assign t[25] = t[29] ^ t[30];
  assign t[26] = t[31] & t[32];
  assign t[27] = t[33] ^ t[26];
  assign t[28] = t[44] ^ t[31];
  assign t[29] = t[45] ^ t[46];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[31] & t[34];
  assign t[31] = ~(t[46]);
  assign t[32] = ~(t[44] ^ t[31]);
  assign t[33] = t[44] & t[35];
  assign t[34] = t[44] ^ t[36];
  assign t[35] = t[37] ^ t[30];
  assign t[36] = t[46] ^ t[47];
  assign t[37] = t[44] ^ t[29];
  assign t[38] = t[48] ^ x[9];
  assign t[39] = t[49] ^ x[17];
  assign t[3] = ~(t[6] ^ t[38]);
  assign t[40] = t[50] ^ x[25];
  assign t[41] = t[51] ^ x[26];
  assign t[42] = t[52] ^ x[27];
  assign t[43] = t[53] ^ x[28];
  assign t[44] = t[54] ^ x[36];
  assign t[45] = t[55] ^ x[37];
  assign t[46] = t[56] ^ x[38];
  assign t[47] = t[57] ^ x[39];
  assign t[48] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[49] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[51] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[52] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[53] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[54] = (x[29] & x[30] & ~x[32] & x[33] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[29] & x[30] & ~x[31] & x[34] & ~x[35]) | (x[29] & ~x[32] & x[33] & x[34] & ~x[35]) | (x[29] & ~x[31] & x[32] & x[33]) | (x[30] & x[31] & ~x[32] & x[34]) | (x[30] & ~x[32] & x[33] & x[34]);
  assign t[55] = (x[29] & x[30] & x[31] & ~x[34] & ~x[35]) | (x[29] & x[30] & x[32] & ~x[33] & ~x[35]) | (x[29] & x[31] & x[32] & ~x[34] & ~x[35]) | (~x[30] & x[31] & x[32] & x[33] & ~x[35]) | (x[30] & x[31] & x[32] & ~x[34]) | (x[30] & x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[33] & x[34]);
  assign t[56] = (x[29] & x[31] & ~x[32] & x[33] & ~x[34]) | (x[29] & x[31] & ~x[32] & ~x[34] & x[35]) | (x[29] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[30] & x[31] & ~x[32] & x[35]) | (x[30] & x[33] & ~x[34] & x[35]) | (x[31] & x[33] & x[35]);
  assign t[57] = (x[30] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[30] & ~x[31] & x[32] & ~x[33] & x[35]) | (x[30] & ~x[31] & ~x[33] & x[34] & x[35]) | (x[29] & x[31] & x[32] & x[33] & x[34]) | (x[29] & ~x[31] & x[32] & x[35]) | (x[29] & ~x[33] & x[34] & x[35]) | (x[32] & x[34] & x[35]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind162(x, y);
 input [29:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[21] ^ t[9]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[15];
  assign t[14] = t[22] ^ t[23];
  assign t[15] = t[16] & t[17];
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[24] ^ t[16]);
  assign t[18] = t[25] ^ x[9];
  assign t[19] = t[26] ^ x[17];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[18];
  assign t[21] = t[28] ^ x[19];
  assign t[22] = t[29] ^ x[27];
  assign t[23] = t[30] ^ x[28];
  assign t[24] = t[31] ^ x[29];
  assign t[25] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[26] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[28] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[29] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[2] = ~(t[4]);
  assign t[30] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[31] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[3] = ~(t[5] ^ t[18]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[19] ^ t[20];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~t[11];
  assign t[9] = ~(t[19]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind163(x, y);
 input [31:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[28]);
  assign t[12] = ~(t[29] ^ t[11]);
  assign t[13] = ~t[15];
  assign t[14] = t[29] ^ t[16];
  assign t[15] = ~(t[17]);
  assign t[16] = t[28] ^ t[30];
  assign t[17] = t[18] ^ t[19];
  assign t[18] = t[20] ^ t[21];
  assign t[19] = t[22] & t[23];
  assign t[1] = ~t[3];
  assign t[20] = t[31] ^ t[32];
  assign t[21] = t[22] & t[24];
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[33] ^ t[22]);
  assign t[24] = t[33] ^ t[25];
  assign t[25] = t[32] ^ t[34];
  assign t[26] = t[35] ^ x[9];
  assign t[27] = t[36] ^ x[17];
  assign t[28] = t[37] ^ x[18];
  assign t[29] = t[38] ^ x[19];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[20];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[29];
  assign t[33] = t[42] ^ x[30];
  assign t[34] = t[43] ^ x[31];
  assign t[35] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[36] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[37] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[38] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[39] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[3] = ~(t[5] ^ t[26]);
  assign t[40] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[41] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[42] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[43] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~t[13];
  assign t[9] = t[27] ^ t[28];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind164(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[8];
  assign t[11] = t[17] ^ t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = ~(t[38]);
  assign t[14] = ~(t[37] ^ t[13]);
  assign t[15] = t[39] ^ t[38];
  assign t[16] = ~(t[21] ^ t[9]);
  assign t[17] = t[22] ^ t[23];
  assign t[18] = t[24] & t[25];
  assign t[19] = t[37] ^ t[15];
  assign t[1] = ~t[3];
  assign t[20] = t[13] & t[21];
  assign t[21] = t[37] ^ t[26];
  assign t[22] = t[40] & t[27];
  assign t[23] = t[28] & t[29];
  assign t[24] = t[30] ^ t[28];
  assign t[25] = t[31] ^ t[23];
  assign t[26] = t[38] ^ t[41];
  assign t[27] = t[32] ^ t[33];
  assign t[28] = ~(t[42]);
  assign t[29] = ~(t[40] ^ t[28]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = t[43] ^ t[42];
  assign t[31] = ~(t[34] ^ t[24]);
  assign t[32] = t[40] ^ t[30];
  assign t[33] = t[28] & t[34];
  assign t[34] = t[40] ^ t[35];
  assign t[35] = t[42] ^ t[44];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[52] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] & t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[37] & t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[13];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind165(x, y);
 input [31:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[37] ^ t[14];
  assign t[11] = ~(t[17] ^ t[18]);
  assign t[12] = t[38] ^ t[39];
  assign t[13] = t[14] & t[19];
  assign t[14] = ~(t[39]);
  assign t[15] = ~(t[37] ^ t[14]);
  assign t[16] = t[37] & t[20];
  assign t[17] = t[21] ^ t[22];
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[37] ^ t[25];
  assign t[1] = ~t[3];
  assign t[20] = t[26] ^ t[13];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[40] ^ t[29];
  assign t[25] = t[39] ^ t[41];
  assign t[26] = t[37] ^ t[12];
  assign t[27] = t[42] ^ t[43];
  assign t[28] = t[29] & t[32];
  assign t[29] = ~(t[43]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[40] ^ t[29]);
  assign t[31] = t[40] & t[33];
  assign t[32] = t[40] ^ t[34];
  assign t[33] = t[35] ^ t[28];
  assign t[34] = t[43] ^ t[44];
  assign t[35] = t[40] ^ t[27];
  assign t[36] = t[45] ^ x[9];
  assign t[37] = t[46] ^ x[17];
  assign t[38] = t[47] ^ x[18];
  assign t[39] = t[48] ^ x[19];
  assign t[3] = ~(t[6] ^ t[36]);
  assign t[40] = t[49] ^ x[27];
  assign t[41] = t[50] ^ x[28];
  assign t[42] = t[51] ^ x[29];
  assign t[43] = t[52] ^ x[30];
  assign t[44] = t[53] ^ x[31];
  assign t[45] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[46] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[47] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[48] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[49] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[5] = t[9] ^ t[10];
  assign t[6] = ~t[11];
  assign t[7] = t[12] ^ t[13];
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind166(x, y);
 input [29:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[19] ^ t[9]);
  assign t[11] = t[12] ^ t[13];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[14] & t[15];
  assign t[14] = ~(t[20]);
  assign t[15] = ~(t[22] ^ t[14]);
  assign t[16] = t[23] ^ x[9];
  assign t[17] = t[24] ^ x[17];
  assign t[18] = t[25] ^ x[18];
  assign t[19] = t[26] ^ x[19];
  assign t[1] = ~t[3];
  assign t[20] = t[27] ^ x[27];
  assign t[21] = t[28] ^ x[28];
  assign t[22] = t[29] ^ x[29];
  assign t[23] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[24] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[25] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[26] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[27] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[28] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[29] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[2] = ~(t[4]);
  assign t[3] = ~(t[5] ^ t[16]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[17] ^ t[18];
  assign t[7] = t[9] & t[10];
  assign t[8] = ~(t[11]);
  assign t[9] = ~(t[17]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind167(x, y);
 input [31:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[27] ^ t[11]);
  assign t[13] = t[15] ^ t[16];
  assign t[14] = t[27] ^ t[17];
  assign t[15] = t[18] ^ t[19];
  assign t[16] = t[20] & t[21];
  assign t[17] = t[26] ^ t[28];
  assign t[18] = t[29] ^ t[30];
  assign t[19] = t[20] & t[22];
  assign t[1] = ~t[3];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[31] ^ t[23];
  assign t[23] = t[30] ^ t[32];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[17];
  assign t[26] = t[35] ^ x[18];
  assign t[27] = t[36] ^ x[19];
  assign t[28] = t[37] ^ x[20];
  assign t[29] = t[38] ^ x[28];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[29];
  assign t[31] = t[40] ^ x[30];
  assign t[32] = t[41] ^ x[31];
  assign t[33] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[34] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[35] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[36] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[37] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[38] = (x[21] & x[22] & x[23] & ~x[26] & ~x[27]) | (x[21] & x[22] & x[24] & ~x[25] & ~x[27]) | (x[21] & x[23] & x[24] & ~x[26] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[22] & x[23] & x[24] & ~x[26]) | (x[22] & x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[25] & x[26]);
  assign t[39] = (x[21] & x[23] & ~x[24] & x[25] & ~x[26]) | (x[21] & x[23] & ~x[24] & ~x[26] & x[27]) | (x[21] & ~x[24] & x[25] & ~x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[22] & x[23] & ~x[24] & x[27]) | (x[22] & x[25] & ~x[26] & x[27]) | (x[23] & x[25] & x[27]);
  assign t[3] = ~(t[5] ^ t[24]);
  assign t[40] = (x[21] & x[22] & ~x[24] & x[25] & ~x[27]) | (~x[22] & x[23] & x[24] & x[25] & ~x[27]) | (x[21] & x[22] & ~x[23] & x[26] & ~x[27]) | (x[21] & ~x[24] & x[25] & x[26] & ~x[27]) | (x[21] & ~x[23] & x[24] & x[25]) | (x[22] & x[23] & ~x[24] & x[26]) | (x[22] & ~x[24] & x[25] & x[26]);
  assign t[41] = (x[22] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[22] & ~x[23] & x[24] & ~x[25] & x[27]) | (x[22] & ~x[23] & ~x[25] & x[26] & x[27]) | (x[21] & x[23] & x[24] & x[25] & x[26]) | (x[21] & ~x[23] & x[24] & x[27]) | (x[21] & ~x[25] & x[26] & x[27]) | (x[24] & x[26] & x[27]);
  assign t[4] = t[6] ^ t[7];
  assign t[5] = ~t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] & t[12];
  assign t[8] = ~(t[13]);
  assign t[9] = t[25] ^ t[26];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind168(x, y);
 input [20:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = t[26] ^ x[19];
  assign t[22] = t[27] ^ x[20];
  assign t[23] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[24] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[25] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[26] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind169(x, y);
 input [20:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = t[26] ^ x[19];
  assign t[22] = t[27] ^ x[20];
  assign t[23] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[24] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[25] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[26] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind170(x, y);
 input [19:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[18];
  assign t[11] = t[15] ^ x[19];
  assign t[12] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[13] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[14] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[15] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[9];
  assign t[9] = t[13] ^ x[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind171(x, y);
 input [20:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[17];
  assign t[14] = t[19] ^ x[18];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[18] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[19] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[1] = ~t[2];
  assign t[20] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[21] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind172(x, y);
 input [20:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = t[26] ^ x[19];
  assign t[22] = t[27] ^ x[20];
  assign t[23] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[24] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[25] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[26] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind173(x, y);
 input [20:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = t[26] ^ x[19];
  assign t[22] = t[27] ^ x[20];
  assign t[23] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[24] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[25] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[26] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind174(x, y);
 input [19:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[18];
  assign t[11] = t[15] ^ x[19];
  assign t[12] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[13] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[14] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[15] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[9];
  assign t[9] = t[13] ^ x[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind175(x, y);
 input [20:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[17];
  assign t[14] = t[19] ^ x[18];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[18] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[19] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[1] = ~t[2];
  assign t[20] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[21] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind176(x, y);
 input [20:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = ~(t[20]);
  assign t[11] = ~(t[19] ^ t[10]);
  assign t[12] = t[21] ^ t[20];
  assign t[13] = ~(t[16] ^ t[7]);
  assign t[14] = t[19] ^ t[12];
  assign t[15] = t[10] & t[16];
  assign t[16] = t[19] ^ t[17];
  assign t[17] = t[20] ^ t[22];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = t[26] ^ x[19];
  assign t[22] = t[27] ^ x[20];
  assign t[23] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[24] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[25] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[26] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = t[3] ^ t[4];
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] & t[8];
  assign t[5] = t[19] & t[9];
  assign t[6] = t[10] & t[11];
  assign t[7] = t[12] ^ t[10];
  assign t[8] = t[13] ^ t[6];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind177(x, y);
 input [20:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(t[1] ^ t[18]);
  assign t[10] = t[11] & t[14];
  assign t[11] = ~(t[21]);
  assign t[12] = ~(t[19] ^ t[11]);
  assign t[13] = t[19] & t[15];
  assign t[14] = t[19] ^ t[16];
  assign t[15] = t[17] ^ t[10];
  assign t[16] = t[21] ^ t[22];
  assign t[17] = t[19] ^ t[9];
  assign t[18] = t[23] ^ x[9];
  assign t[19] = t[24] ^ x[17];
  assign t[1] = ~t[2];
  assign t[20] = t[25] ^ x[18];
  assign t[21] = t[26] ^ x[19];
  assign t[22] = t[27] ^ x[20];
  assign t[23] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[24] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[25] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[26] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[27] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = ~(t[3] ^ t[4]);
  assign t[3] = t[5] ^ t[6];
  assign t[4] = t[7] ^ t[8];
  assign t[5] = t[9] ^ t[10];
  assign t[6] = t[11] & t[12];
  assign t[7] = t[13] ^ t[6];
  assign t[8] = t[19] ^ t[11];
  assign t[9] = t[20] ^ t[21];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind178(x, y);
 input [19:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[1] ^ t[8]);
  assign t[10] = t[14] ^ x[18];
  assign t[11] = t[15] ^ x[19];
  assign t[12] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[13] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[14] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[15] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[9] ^ t[10];
  assign t[5] = t[6] & t[7];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[11] ^ t[6]);
  assign t[8] = t[12] ^ x[9];
  assign t[9] = t[13] ^ x[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind179(x, y);
 input [20:0] x;
 output y;

 wire [21:0] t;
  assign t[0] = ~(t[1] ^ t[12]);
  assign t[10] = t[15] ^ t[11];
  assign t[11] = t[14] ^ t[16];
  assign t[12] = t[17] ^ x[9];
  assign t[13] = t[18] ^ x[17];
  assign t[14] = t[19] ^ x[18];
  assign t[15] = t[20] ^ x[19];
  assign t[16] = t[21] ^ x[20];
  assign t[17] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[18] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[19] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[1] = ~t[2];
  assign t[20] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[21] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[2] = ~(t[3]);
  assign t[3] = t[4] ^ t[5];
  assign t[4] = t[6] ^ t[7];
  assign t[5] = t[8] & t[9];
  assign t[6] = t[13] ^ t[14];
  assign t[7] = t[8] & t[10];
  assign t[8] = ~(t[14]);
  assign t[9] = ~(t[15] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind180(x, y);
 input [28:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[15] ^ t[8];
  assign t[11] = t[16] ^ t[17];
  assign t[12] = ~(t[23]);
  assign t[13] = ~(t[22] ^ t[12]);
  assign t[14] = t[24] ^ t[23];
  assign t[15] = ~(t[18] ^ t[9]);
  assign t[16] = t[22] ^ t[14];
  assign t[17] = t[12] & t[18];
  assign t[18] = t[22] ^ t[19];
  assign t[19] = t[23] ^ t[25];
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[9];
  assign t[21] = t[27] ^ x[17];
  assign t[22] = t[28] ^ x[25];
  assign t[23] = t[29] ^ x[26];
  assign t[24] = t[30] ^ x[27];
  assign t[25] = t[31] ^ x[28];
  assign t[26] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[27] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[28] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[29] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[31] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[3] = ~t[4];
  assign t[4] = t[5] ^ t[6];
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] & t[10];
  assign t[7] = t[22] & t[11];
  assign t[8] = t[12] & t[13];
  assign t[9] = t[14] ^ t[12];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind181(x, y);
 input [28:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[1] ^ t[20]);
  assign t[10] = t[22] ^ t[13];
  assign t[11] = t[23] ^ t[24];
  assign t[12] = t[13] & t[16];
  assign t[13] = ~(t[24]);
  assign t[14] = ~(t[22] ^ t[13]);
  assign t[15] = t[22] & t[17];
  assign t[16] = t[22] ^ t[18];
  assign t[17] = t[19] ^ t[12];
  assign t[18] = t[24] ^ t[25];
  assign t[19] = t[22] ^ t[11];
  assign t[1] = ~t[2];
  assign t[20] = t[26] ^ x[9];
  assign t[21] = t[27] ^ x[17];
  assign t[22] = t[28] ^ x[25];
  assign t[23] = t[29] ^ x[26];
  assign t[24] = t[30] ^ x[27];
  assign t[25] = t[31] ^ x[28];
  assign t[26] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[27] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[28] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[29] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[2] = ~(t[3] ^ t[21]);
  assign t[30] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[31] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5] ^ t[6]);
  assign t[5] = t[7] ^ t[8];
  assign t[6] = t[9] ^ t[10];
  assign t[7] = t[11] ^ t[12];
  assign t[8] = t[13] & t[14];
  assign t[9] = t[15] ^ t[8];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind182(x, y);
 input [27:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~(t[1] ^ t[10]);
  assign t[10] = t[15] ^ x[9];
  assign t[11] = t[16] ^ x[17];
  assign t[12] = t[17] ^ x[25];
  assign t[13] = t[18] ^ x[26];
  assign t[14] = t[19] ^ x[27];
  assign t[15] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[16] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[17] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[18] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[19] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[1] = ~t[2];
  assign t[2] = ~(t[3] ^ t[11]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[12] ^ t[13];
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[14] ^ t[8]);
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind183(x, y);
 input [28:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[1] ^ t[14]);
  assign t[10] = ~(t[17]);
  assign t[11] = ~(t[18] ^ t[10]);
  assign t[12] = t[18] ^ t[13];
  assign t[13] = t[17] ^ t[19];
  assign t[14] = t[20] ^ x[9];
  assign t[15] = t[21] ^ x[17];
  assign t[16] = t[22] ^ x[25];
  assign t[17] = t[23] ^ x[26];
  assign t[18] = t[24] ^ x[27];
  assign t[19] = t[25] ^ x[28];
  assign t[1] = ~t[2];
  assign t[20] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[21] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[22] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[23] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[24] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[25] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[2] = ~(t[3] ^ t[15]);
  assign t[3] = ~t[4];
  assign t[4] = ~(t[5]);
  assign t[5] = t[6] ^ t[7];
  assign t[6] = t[8] ^ t[9];
  assign t[7] = t[10] & t[11];
  assign t[8] = t[16] ^ t[17];
  assign t[9] = t[10] & t[12];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind184(x, y);
 input [42:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[9];
  assign t[53] = t[66] ^ x[17];
  assign t[54] = t[67] ^ x[25];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[34];
  assign t[57] = t[70] ^ x[35];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[37];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[38];
  assign t[61] = t[74] ^ x[39];
  assign t[62] = t[75] ^ x[40];
  assign t[63] = t[76] ^ x[41];
  assign t[64] = t[77] ^ x[42];
  assign t[65] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[66] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[67] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[68] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[69] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[71] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[72] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[73] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[74] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[75] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[76] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[77] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind185(x, y);
 input [42:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] ^ t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] ^ t[24];
  assign t[13] = t[25] ^ t[26];
  assign t[14] = t[27] & t[28];
  assign t[15] = t[29] ^ t[14];
  assign t[16] = t[53] ^ t[27];
  assign t[17] = t[30] ^ t[31];
  assign t[18] = t[32] & t[33];
  assign t[19] = t[34] ^ t[18];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[54] ^ t[32];
  assign t[21] = t[35] ^ t[36];
  assign t[22] = t[37] & t[38];
  assign t[23] = t[39] ^ t[22];
  assign t[24] = t[55] ^ t[37];
  assign t[25] = t[56] ^ t[57];
  assign t[26] = t[27] & t[40];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[53] ^ t[27]);
  assign t[29] = t[53] & t[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[58] ^ t[59];
  assign t[31] = t[32] & t[42];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[43];
  assign t[35] = t[60] ^ t[61];
  assign t[36] = t[37] & t[44];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[55] ^ t[37]);
  assign t[39] = t[55] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[46];
  assign t[41] = t[47] ^ t[26];
  assign t[42] = t[54] ^ t[48];
  assign t[43] = t[49] ^ t[31];
  assign t[44] = t[55] ^ t[50];
  assign t[45] = t[51] ^ t[36];
  assign t[46] = t[57] ^ t[62];
  assign t[47] = t[53] ^ t[25];
  assign t[48] = t[59] ^ t[63];
  assign t[49] = t[54] ^ t[30];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[61] ^ t[64];
  assign t[51] = t[55] ^ t[35];
  assign t[52] = t[65] ^ x[9];
  assign t[53] = t[66] ^ x[17];
  assign t[54] = t[67] ^ x[25];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[34];
  assign t[57] = t[70] ^ x[35];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[37];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[73] ^ x[38];
  assign t[61] = t[74] ^ x[39];
  assign t[62] = t[75] ^ x[40];
  assign t[63] = t[76] ^ x[41];
  assign t[64] = t[77] ^ x[42];
  assign t[65] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[66] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[67] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[68] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[69] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[71] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[72] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[73] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[74] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[75] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[76] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[77] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind186(x, y);
 input [39:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[9];
  assign t[23] = t[33] ^ x[17];
  assign t[24] = t[34] ^ x[18];
  assign t[25] = t[35] ^ x[26];
  assign t[26] = t[36] ^ x[27];
  assign t[27] = t[37] ^ x[35];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[37];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[38];
  assign t[31] = t[41] ^ x[39];
  assign t[32] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[33] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[34] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[35] = (x[19] & x[21] & ~x[22] & x[23] & ~x[24]) | (x[19] & x[21] & ~x[22] & ~x[24] & x[25]) | (x[19] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[19] & x[21] & x[22] & x[23] & x[24]) | (x[20] & x[21] & ~x[22] & x[25]) | (x[20] & x[23] & ~x[24] & x[25]) | (x[21] & x[23] & x[25]);
  assign t[36] = (x[20] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[20] & ~x[21] & x[22] & ~x[23] & x[25]) | (x[20] & ~x[21] & ~x[23] & x[24] & x[25]) | (x[19] & x[21] & x[22] & x[23] & x[24]) | (x[19] & ~x[21] & x[22] & x[25]) | (x[19] & ~x[23] & x[24] & x[25]) | (x[22] & x[24] & x[25]);
  assign t[37] = (x[28] & x[30] & ~x[31] & x[32] & ~x[33]) | (x[28] & x[30] & ~x[31] & ~x[33] & x[34]) | (x[28] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[29] & x[30] & ~x[31] & x[34]) | (x[29] & x[32] & ~x[33] & x[34]) | (x[30] & x[32] & x[34]);
  assign t[38] = (x[29] & ~x[30] & x[31] & ~x[32] & x[33]) | (x[29] & ~x[30] & x[31] & ~x[32] & x[34]) | (x[29] & ~x[30] & ~x[32] & x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[28] & ~x[30] & x[31] & x[34]) | (x[28] & ~x[32] & x[33] & x[34]) | (x[31] & x[33] & x[34]);
  assign t[39] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[3] = ~t[6];
  assign t[40] = (x[19] & x[20] & ~x[22] & x[23] & ~x[25]) | (~x[20] & x[21] & x[22] & x[23] & ~x[25]) | (x[19] & x[20] & ~x[21] & x[24] & ~x[25]) | (x[19] & ~x[22] & x[23] & x[24] & ~x[25]) | (x[19] & ~x[21] & x[22] & x[23]) | (x[20] & x[21] & ~x[22] & x[24]) | (x[20] & ~x[22] & x[23] & x[24]);
  assign t[41] = (x[28] & x[29] & ~x[31] & x[32] & ~x[34]) | (~x[29] & x[30] & x[31] & x[32] & ~x[34]) | (x[28] & x[29] & ~x[30] & x[33] & ~x[34]) | (x[28] & ~x[31] & x[32] & x[33] & ~x[34]) | (x[28] & ~x[30] & x[31] & x[32]) | (x[29] & x[30] & ~x[31] & x[33]) | (x[29] & ~x[31] & x[32] & x[33]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind187(x, y);
 input [42:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[9];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[18];
  assign t[37] = t[50] ^ x[19];
  assign t[38] = t[51] ^ x[27];
  assign t[39] = t[52] ^ x[28];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[29];
  assign t[41] = t[54] ^ x[37];
  assign t[42] = t[55] ^ x[38];
  assign t[43] = t[56] ^ x[39];
  assign t[44] = t[57] ^ x[40];
  assign t[45] = t[58] ^ x[41];
  assign t[46] = t[59] ^ x[42];
  assign t[47] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[54] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[55] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[56] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[57] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[58] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[59] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind188(x, y);
 input [42:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[9];
  assign t[53] = t[66] ^ x[17];
  assign t[54] = t[67] ^ x[25];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[34];
  assign t[57] = t[70] ^ x[35];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[37];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[38];
  assign t[61] = t[74] ^ x[39];
  assign t[62] = t[75] ^ x[40];
  assign t[63] = t[76] ^ x[41];
  assign t[64] = t[77] ^ x[42];
  assign t[65] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[66] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[67] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[68] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[69] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[71] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[72] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[73] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[74] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[75] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[76] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[77] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind189(x, y);
 input [42:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = t[20] ^ t[21];
  assign t[12] = t[22] ^ t[23];
  assign t[13] = t[24] ^ t[25];
  assign t[14] = t[26] ^ t[27];
  assign t[15] = t[28] & t[29];
  assign t[16] = t[30] ^ t[15];
  assign t[17] = t[54] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[3] ^ t[53]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[55] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[56] ^ t[38];
  assign t[26] = t[57] ^ t[58];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[58]);
  assign t[29] = ~(t[54] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[54] & t[42];
  assign t[31] = t[59] ^ t[60];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[60]);
  assign t[34] = ~(t[55] ^ t[33]);
  assign t[35] = t[55] & t[44];
  assign t[36] = t[61] ^ t[62];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[62]);
  assign t[39] = ~(t[56] ^ t[38]);
  assign t[3] = ~t[6];
  assign t[40] = t[56] & t[46];
  assign t[41] = t[54] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[55] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[56] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[58] ^ t[63];
  assign t[48] = t[54] ^ t[26];
  assign t[49] = t[60] ^ t[64];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] ^ t[31];
  assign t[51] = t[62] ^ t[65];
  assign t[52] = t[56] ^ t[36];
  assign t[53] = t[66] ^ x[9];
  assign t[54] = t[67] ^ x[17];
  assign t[55] = t[68] ^ x[25];
  assign t[56] = t[69] ^ x[33];
  assign t[57] = t[70] ^ x[34];
  assign t[58] = t[71] ^ x[35];
  assign t[59] = t[72] ^ x[36];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = t[73] ^ x[37];
  assign t[61] = t[74] ^ x[38];
  assign t[62] = t[75] ^ x[39];
  assign t[63] = t[76] ^ x[40];
  assign t[64] = t[77] ^ x[41];
  assign t[65] = t[78] ^ x[42];
  assign t[66] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[67] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[68] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[69] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[71] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[72] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[73] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[74] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[75] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[76] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[77] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[78] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[8] = t[14] ^ t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind190(x, y);
 input [39:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[9];
  assign t[23] = t[33] ^ x[17];
  assign t[24] = t[34] ^ x[18];
  assign t[25] = t[35] ^ x[26];
  assign t[26] = t[36] ^ x[27];
  assign t[27] = t[37] ^ x[35];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[37];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[38];
  assign t[31] = t[41] ^ x[39];
  assign t[32] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[33] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[34] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[35] = (x[19] & x[21] & ~x[22] & x[23] & ~x[24]) | (x[19] & x[21] & ~x[22] & ~x[24] & x[25]) | (x[19] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[19] & x[21] & x[22] & x[23] & x[24]) | (x[20] & x[21] & ~x[22] & x[25]) | (x[20] & x[23] & ~x[24] & x[25]) | (x[21] & x[23] & x[25]);
  assign t[36] = (x[20] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[20] & ~x[21] & x[22] & ~x[23] & x[25]) | (x[20] & ~x[21] & ~x[23] & x[24] & x[25]) | (x[19] & x[21] & x[22] & x[23] & x[24]) | (x[19] & ~x[21] & x[22] & x[25]) | (x[19] & ~x[23] & x[24] & x[25]) | (x[22] & x[24] & x[25]);
  assign t[37] = (x[28] & x[30] & ~x[31] & x[32] & ~x[33]) | (x[28] & x[30] & ~x[31] & ~x[33] & x[34]) | (x[28] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[29] & x[30] & ~x[31] & x[34]) | (x[29] & x[32] & ~x[33] & x[34]) | (x[30] & x[32] & x[34]);
  assign t[38] = (x[29] & ~x[30] & x[31] & ~x[32] & x[33]) | (x[29] & ~x[30] & x[31] & ~x[32] & x[34]) | (x[29] & ~x[30] & ~x[32] & x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[28] & ~x[30] & x[31] & x[34]) | (x[28] & ~x[32] & x[33] & x[34]) | (x[31] & x[33] & x[34]);
  assign t[39] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[3] = ~t[6];
  assign t[40] = (x[19] & x[20] & ~x[22] & x[23] & ~x[25]) | (~x[20] & x[21] & x[22] & x[23] & ~x[25]) | (x[19] & x[20] & ~x[21] & x[24] & ~x[25]) | (x[19] & ~x[22] & x[23] & x[24] & ~x[25]) | (x[19] & ~x[21] & x[22] & x[23]) | (x[20] & x[21] & ~x[22] & x[24]) | (x[20] & ~x[22] & x[23] & x[24]);
  assign t[41] = (x[28] & x[29] & ~x[31] & x[32] & ~x[34]) | (~x[29] & x[30] & x[31] & x[32] & ~x[34]) | (x[28] & x[29] & ~x[30] & x[33] & ~x[34]) | (x[28] & ~x[31] & x[32] & x[33] & ~x[34]) | (x[28] & ~x[30] & x[31] & x[32]) | (x[29] & x[30] & ~x[31] & x[33]) | (x[29] & ~x[31] & x[32] & x[33]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind191(x, y);
 input [42:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[9];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[18];
  assign t[37] = t[50] ^ x[19];
  assign t[38] = t[51] ^ x[27];
  assign t[39] = t[52] ^ x[28];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[29];
  assign t[41] = t[54] ^ x[37];
  assign t[42] = t[55] ^ x[38];
  assign t[43] = t[56] ^ x[39];
  assign t[44] = t[57] ^ x[40];
  assign t[45] = t[58] ^ x[41];
  assign t[46] = t[59] ^ x[42];
  assign t[47] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[54] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[55] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[56] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[57] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[58] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[59] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind192(x, y);
 input [42:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] & t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] & t[24];
  assign t[13] = t[53] & t[25];
  assign t[14] = t[26] & t[27];
  assign t[15] = t[28] ^ t[26];
  assign t[16] = t[29] ^ t[14];
  assign t[17] = t[54] & t[30];
  assign t[18] = t[31] & t[32];
  assign t[19] = t[33] ^ t[31];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[34] ^ t[18];
  assign t[21] = t[55] & t[35];
  assign t[22] = t[36] & t[37];
  assign t[23] = t[38] ^ t[36];
  assign t[24] = t[39] ^ t[22];
  assign t[25] = t[40] ^ t[41];
  assign t[26] = ~(t[56]);
  assign t[27] = ~(t[53] ^ t[26]);
  assign t[28] = t[57] ^ t[56];
  assign t[29] = ~(t[42] ^ t[15]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[44];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[54] ^ t[31]);
  assign t[33] = t[59] ^ t[58];
  assign t[34] = ~(t[45] ^ t[19]);
  assign t[35] = t[46] ^ t[47];
  assign t[36] = ~(t[60]);
  assign t[37] = ~(t[55] ^ t[36]);
  assign t[38] = t[61] ^ t[60];
  assign t[39] = ~(t[48] ^ t[23]);
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[28];
  assign t[41] = t[26] & t[42];
  assign t[42] = t[53] ^ t[49];
  assign t[43] = t[54] ^ t[33];
  assign t[44] = t[31] & t[45];
  assign t[45] = t[54] ^ t[50];
  assign t[46] = t[55] ^ t[38];
  assign t[47] = t[36] & t[48];
  assign t[48] = t[55] ^ t[51];
  assign t[49] = t[56] ^ t[62];
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[58] ^ t[63];
  assign t[51] = t[60] ^ t[64];
  assign t[52] = t[65] ^ x[9];
  assign t[53] = t[66] ^ x[17];
  assign t[54] = t[67] ^ x[25];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[34];
  assign t[57] = t[70] ^ x[35];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[37];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[73] ^ x[38];
  assign t[61] = t[74] ^ x[39];
  assign t[62] = t[75] ^ x[40];
  assign t[63] = t[76] ^ x[41];
  assign t[64] = t[77] ^ x[42];
  assign t[65] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[66] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[67] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[68] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[69] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[6] = t[11] ^ t[12];
  assign t[70] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[71] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[72] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[73] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[74] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[75] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[76] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[77] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] & t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind193(x, y);
 input [42:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[19] ^ t[20];
  assign t[11] = t[21] ^ t[22];
  assign t[12] = t[23] ^ t[24];
  assign t[13] = t[25] ^ t[26];
  assign t[14] = t[27] & t[28];
  assign t[15] = t[29] ^ t[14];
  assign t[16] = t[53] ^ t[27];
  assign t[17] = t[30] ^ t[31];
  assign t[18] = t[32] & t[33];
  assign t[19] = t[34] ^ t[18];
  assign t[1] = ~(t[3] ^ t[52]);
  assign t[20] = t[54] ^ t[32];
  assign t[21] = t[35] ^ t[36];
  assign t[22] = t[37] & t[38];
  assign t[23] = t[39] ^ t[22];
  assign t[24] = t[55] ^ t[37];
  assign t[25] = t[56] ^ t[57];
  assign t[26] = t[27] & t[40];
  assign t[27] = ~(t[57]);
  assign t[28] = ~(t[53] ^ t[27]);
  assign t[29] = t[53] & t[41];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[58] ^ t[59];
  assign t[31] = t[32] & t[42];
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[43];
  assign t[35] = t[60] ^ t[61];
  assign t[36] = t[37] & t[44];
  assign t[37] = ~(t[61]);
  assign t[38] = ~(t[55] ^ t[37]);
  assign t[39] = t[55] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ t[46];
  assign t[41] = t[47] ^ t[26];
  assign t[42] = t[54] ^ t[48];
  assign t[43] = t[49] ^ t[31];
  assign t[44] = t[55] ^ t[50];
  assign t[45] = t[51] ^ t[36];
  assign t[46] = t[57] ^ t[62];
  assign t[47] = t[53] ^ t[25];
  assign t[48] = t[59] ^ t[63];
  assign t[49] = t[54] ^ t[30];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[61] ^ t[64];
  assign t[51] = t[55] ^ t[35];
  assign t[52] = t[65] ^ x[9];
  assign t[53] = t[66] ^ x[17];
  assign t[54] = t[67] ^ x[25];
  assign t[55] = t[68] ^ x[33];
  assign t[56] = t[69] ^ x[34];
  assign t[57] = t[70] ^ x[35];
  assign t[58] = t[71] ^ x[36];
  assign t[59] = t[72] ^ x[37];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[73] ^ x[38];
  assign t[61] = t[74] ^ x[39];
  assign t[62] = t[75] ^ x[40];
  assign t[63] = t[76] ^ x[41];
  assign t[64] = t[77] ^ x[42];
  assign t[65] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[66] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[67] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[68] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[69] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[71] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[72] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[73] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[74] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[75] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[76] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[77] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[7] = t[13] ^ t[14];
  assign t[8] = t[15] ^ t[16];
  assign t[9] = t[17] ^ t[18];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind194(x, y);
 input [39:0] x;
 output y;

 wire [41:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[23] ^ t[24];
  assign t[11] = t[16] & t[17];
  assign t[12] = t[25] ^ t[26];
  assign t[13] = t[18] & t[19];
  assign t[14] = t[27] ^ t[28];
  assign t[15] = t[20] & t[21];
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[29] ^ t[16]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[30] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[22]);
  assign t[20] = ~(t[27]);
  assign t[21] = ~(t[31] ^ t[20]);
  assign t[22] = t[32] ^ x[9];
  assign t[23] = t[33] ^ x[17];
  assign t[24] = t[34] ^ x[18];
  assign t[25] = t[35] ^ x[26];
  assign t[26] = t[36] ^ x[27];
  assign t[27] = t[37] ^ x[35];
  assign t[28] = t[38] ^ x[36];
  assign t[29] = t[39] ^ x[37];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[40] ^ x[38];
  assign t[31] = t[41] ^ x[39];
  assign t[32] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[33] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[34] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[35] = (x[19] & x[21] & ~x[22] & x[23] & ~x[24]) | (x[19] & x[21] & ~x[22] & ~x[24] & x[25]) | (x[19] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[19] & x[21] & x[22] & x[23] & x[24]) | (x[20] & x[21] & ~x[22] & x[25]) | (x[20] & x[23] & ~x[24] & x[25]) | (x[21] & x[23] & x[25]);
  assign t[36] = (x[20] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[20] & ~x[21] & x[22] & ~x[23] & x[25]) | (x[20] & ~x[21] & ~x[23] & x[24] & x[25]) | (x[19] & x[21] & x[22] & x[23] & x[24]) | (x[19] & ~x[21] & x[22] & x[25]) | (x[19] & ~x[23] & x[24] & x[25]) | (x[22] & x[24] & x[25]);
  assign t[37] = (x[28] & x[30] & ~x[31] & x[32] & ~x[33]) | (x[28] & x[30] & ~x[31] & ~x[33] & x[34]) | (x[28] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[29] & x[30] & ~x[31] & x[34]) | (x[29] & x[32] & ~x[33] & x[34]) | (x[30] & x[32] & x[34]);
  assign t[38] = (x[29] & ~x[30] & x[31] & ~x[32] & x[33]) | (x[29] & ~x[30] & x[31] & ~x[32] & x[34]) | (x[29] & ~x[30] & ~x[32] & x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[28] & ~x[30] & x[31] & x[34]) | (x[28] & ~x[32] & x[33] & x[34]) | (x[31] & x[33] & x[34]);
  assign t[39] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[3] = ~t[6];
  assign t[40] = (x[19] & x[20] & ~x[22] & x[23] & ~x[25]) | (~x[20] & x[21] & x[22] & x[23] & ~x[25]) | (x[19] & x[20] & ~x[21] & x[24] & ~x[25]) | (x[19] & ~x[22] & x[23] & x[24] & ~x[25]) | (x[19] & ~x[21] & x[22] & x[23]) | (x[20] & x[21] & ~x[22] & x[24]) | (x[20] & ~x[22] & x[23] & x[24]);
  assign t[41] = (x[28] & x[29] & ~x[31] & x[32] & ~x[34]) | (~x[29] & x[30] & x[31] & x[32] & ~x[34]) | (x[28] & x[29] & ~x[30] & x[33] & ~x[34]) | (x[28] & ~x[31] & x[32] & x[33] & ~x[34]) | (x[28] & ~x[30] & x[31] & x[32]) | (x[29] & x[30] & ~x[31] & x[33]) | (x[29] & ~x[31] & x[32] & x[33]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind195(x, y);
 input [42:0] x;
 output y;

 wire [59:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] ^ t[17];
  assign t[11] = t[18] & t[19];
  assign t[12] = t[20] ^ t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[25];
  assign t[15] = t[26] & t[27];
  assign t[16] = t[35] ^ t[36];
  assign t[17] = t[18] & t[28];
  assign t[18] = ~(t[36]);
  assign t[19] = ~(t[37] ^ t[18]);
  assign t[1] = ~(t[3] ^ t[34]);
  assign t[20] = t[38] ^ t[39];
  assign t[21] = t[22] & t[29];
  assign t[22] = ~(t[39]);
  assign t[23] = ~(t[40] ^ t[22]);
  assign t[24] = t[41] ^ t[42];
  assign t[25] = t[26] & t[30];
  assign t[26] = ~(t[42]);
  assign t[27] = ~(t[43] ^ t[26]);
  assign t[28] = t[37] ^ t[31];
  assign t[29] = t[40] ^ t[32];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[43] ^ t[33];
  assign t[31] = t[36] ^ t[44];
  assign t[32] = t[39] ^ t[45];
  assign t[33] = t[42] ^ t[46];
  assign t[34] = t[47] ^ x[9];
  assign t[35] = t[48] ^ x[17];
  assign t[36] = t[49] ^ x[18];
  assign t[37] = t[50] ^ x[19];
  assign t[38] = t[51] ^ x[27];
  assign t[39] = t[52] ^ x[28];
  assign t[3] = ~t[6];
  assign t[40] = t[53] ^ x[29];
  assign t[41] = t[54] ^ x[37];
  assign t[42] = t[55] ^ x[38];
  assign t[43] = t[56] ^ x[39];
  assign t[44] = t[57] ^ x[40];
  assign t[45] = t[58] ^ x[41];
  assign t[46] = t[59] ^ x[42];
  assign t[47] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[48] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[49] = (x[10] & x[12] & ~x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[13] & ~x[15] & x[16]) | (x[10] & ~x[13] & x[14] & ~x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[11] & x[12] & ~x[13] & x[16]) | (x[11] & x[14] & ~x[15] & x[16]) | (x[12] & x[14] & x[16]);
  assign t[4] = ~(t[7]);
  assign t[50] = (x[10] & x[11] & ~x[13] & x[14] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[10] & x[11] & ~x[12] & x[15] & ~x[16]) | (x[10] & ~x[13] & x[14] & x[15] & ~x[16]) | (x[10] & ~x[12] & x[13] & x[14]) | (x[11] & x[12] & ~x[13] & x[15]) | (x[11] & ~x[13] & x[14] & x[15]);
  assign t[51] = (x[20] & x[21] & x[22] & ~x[25] & ~x[26]) | (x[20] & x[21] & x[23] & ~x[24] & ~x[26]) | (x[20] & x[22] & x[23] & ~x[25] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[21] & x[22] & x[23] & ~x[25]) | (x[21] & x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[24] & x[25]);
  assign t[52] = (x[20] & x[22] & ~x[23] & x[24] & ~x[25]) | (x[20] & x[22] & ~x[23] & ~x[25] & x[26]) | (x[20] & ~x[23] & x[24] & ~x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[21] & x[22] & ~x[23] & x[26]) | (x[21] & x[24] & ~x[25] & x[26]) | (x[22] & x[24] & x[26]);
  assign t[53] = (x[20] & x[21] & ~x[23] & x[24] & ~x[26]) | (~x[21] & x[22] & x[23] & x[24] & ~x[26]) | (x[20] & x[21] & ~x[22] & x[25] & ~x[26]) | (x[20] & ~x[23] & x[24] & x[25] & ~x[26]) | (x[20] & ~x[22] & x[23] & x[24]) | (x[21] & x[22] & ~x[23] & x[25]) | (x[21] & ~x[23] & x[24] & x[25]);
  assign t[54] = (x[30] & x[31] & x[32] & ~x[35] & ~x[36]) | (x[30] & x[31] & x[33] & ~x[34] & ~x[36]) | (x[30] & x[32] & x[33] & ~x[35] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[31] & x[32] & x[33] & ~x[35]) | (x[31] & x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[34] & x[35]);
  assign t[55] = (x[30] & x[32] & ~x[33] & x[34] & ~x[35]) | (x[30] & x[32] & ~x[33] & ~x[35] & x[36]) | (x[30] & ~x[33] & x[34] & ~x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[31] & x[32] & ~x[33] & x[36]) | (x[31] & x[34] & ~x[35] & x[36]) | (x[32] & x[34] & x[36]);
  assign t[56] = (x[30] & x[31] & ~x[33] & x[34] & ~x[36]) | (~x[31] & x[32] & x[33] & x[34] & ~x[36]) | (x[30] & x[31] & ~x[32] & x[35] & ~x[36]) | (x[30] & ~x[33] & x[34] & x[35] & ~x[36]) | (x[30] & ~x[32] & x[33] & x[34]) | (x[31] & x[32] & ~x[33] & x[35]) | (x[31] & ~x[33] & x[34] & x[35]);
  assign t[57] = (x[11] & ~x[12] & x[13] & ~x[14] & x[15]) | (x[11] & ~x[12] & x[13] & ~x[14] & x[16]) | (x[11] & ~x[12] & ~x[14] & x[15] & x[16]) | (x[10] & x[12] & x[13] & x[14] & x[15]) | (x[10] & ~x[12] & x[13] & x[16]) | (x[10] & ~x[14] & x[15] & x[16]) | (x[13] & x[15] & x[16]);
  assign t[58] = (x[21] & ~x[22] & x[23] & ~x[24] & x[25]) | (x[21] & ~x[22] & x[23] & ~x[24] & x[26]) | (x[21] & ~x[22] & ~x[24] & x[25] & x[26]) | (x[20] & x[22] & x[23] & x[24] & x[25]) | (x[20] & ~x[22] & x[23] & x[26]) | (x[20] & ~x[24] & x[25] & x[26]) | (x[23] & x[25] & x[26]);
  assign t[59] = (x[31] & ~x[32] & x[33] & ~x[34] & x[35]) | (x[31] & ~x[32] & x[33] & ~x[34] & x[36]) | (x[31] & ~x[32] & ~x[34] & x[35] & x[36]) | (x[30] & x[32] & x[33] & x[34] & x[35]) | (x[30] & ~x[32] & x[33] & x[36]) | (x[30] & ~x[34] & x[35] & x[36]) | (x[33] & x[35] & x[36]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = t[14] ^ t[15];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind196(x, y);
 input [50:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] & t[19];
  assign t[11] = ~t[20];
  assign t[12] = t[56] & t[21];
  assign t[13] = t[22] & t[23];
  assign t[14] = t[24] ^ t[22];
  assign t[15] = t[25] ^ t[13];
  assign t[16] = t[57] & t[26];
  assign t[17] = t[27] & t[28];
  assign t[18] = t[29] ^ t[27];
  assign t[19] = t[30] ^ t[17];
  assign t[1] = ~(t[3] ^ t[54]);
  assign t[20] = t[31] ^ t[32];
  assign t[21] = t[33] ^ t[34];
  assign t[22] = ~(t[58]);
  assign t[23] = ~(t[56] ^ t[22]);
  assign t[24] = t[59] ^ t[58];
  assign t[25] = ~(t[35] ^ t[14]);
  assign t[26] = t[36] ^ t[37];
  assign t[27] = ~(t[60]);
  assign t[28] = ~(t[57] ^ t[27]);
  assign t[29] = t[61] ^ t[60];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = ~(t[38] ^ t[18]);
  assign t[31] = t[39] ^ t[40];
  assign t[32] = t[41] & t[42];
  assign t[33] = t[56] ^ t[24];
  assign t[34] = t[22] & t[35];
  assign t[35] = t[56] ^ t[43];
  assign t[36] = t[57] ^ t[29];
  assign t[37] = t[27] & t[38];
  assign t[38] = t[57] ^ t[44];
  assign t[39] = t[62] & t[45];
  assign t[3] = ~t[6];
  assign t[40] = t[46] & t[47];
  assign t[41] = t[48] ^ t[46];
  assign t[42] = t[49] ^ t[40];
  assign t[43] = t[58] ^ t[63];
  assign t[44] = t[60] ^ t[64];
  assign t[45] = t[50] ^ t[51];
  assign t[46] = ~(t[65]);
  assign t[47] = ~(t[62] ^ t[46]);
  assign t[48] = t[66] ^ t[65];
  assign t[49] = ~(t[52] ^ t[41]);
  assign t[4] = t[7] ^ t[8];
  assign t[50] = t[62] ^ t[48];
  assign t[51] = t[46] & t[52];
  assign t[52] = t[62] ^ t[53];
  assign t[53] = t[65] ^ t[67];
  assign t[54] = t[68] ^ x[9];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[25];
  assign t[57] = t[71] ^ x[33];
  assign t[58] = t[72] ^ x[34];
  assign t[59] = t[73] ^ x[35];
  assign t[5] = t[9] ^ t[10];
  assign t[60] = t[74] ^ x[36];
  assign t[61] = t[75] ^ x[37];
  assign t[62] = t[76] ^ x[45];
  assign t[63] = t[77] ^ x[46];
  assign t[64] = t[78] ^ x[47];
  assign t[65] = t[79] ^ x[48];
  assign t[66] = t[80] ^ x[49];
  assign t[67] = t[81] ^ x[50];
  assign t[68] = (x[2] & x[3] & x[4] & ~x[7] & ~x[8]) | (x[2] & x[3] & x[5] & ~x[6] & ~x[8]) | (x[2] & x[4] & x[5] & ~x[7] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[3] & x[4] & x[5] & ~x[7]) | (x[3] & x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[6] & x[7]);
  assign t[69] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[6] = ~(t[11] ^ t[55]);
  assign t[70] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[71] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[72] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[73] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[74] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[75] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[76] = (x[38] & x[39] & ~x[41] & x[42] & ~x[44]) | (~x[39] & x[40] & x[41] & x[42] & ~x[44]) | (x[38] & x[39] & ~x[40] & x[43] & ~x[44]) | (x[38] & ~x[41] & x[42] & x[43] & ~x[44]) | (x[38] & ~x[40] & x[41] & x[42]) | (x[39] & x[40] & ~x[41] & x[43]) | (x[39] & ~x[41] & x[42] & x[43]);
  assign t[77] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[78] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[79] = (x[38] & x[40] & ~x[41] & x[42] & ~x[43]) | (x[38] & x[40] & ~x[41] & ~x[43] & x[44]) | (x[38] & ~x[41] & x[42] & ~x[43] & x[44]) | (x[38] & x[40] & x[41] & x[42] & x[43]) | (x[39] & x[40] & ~x[41] & x[44]) | (x[39] & x[42] & ~x[43] & x[44]) | (x[40] & x[42] & x[44]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[38] & x[39] & x[40] & ~x[43] & ~x[44]) | (x[38] & x[39] & x[41] & ~x[42] & ~x[44]) | (x[38] & x[40] & x[41] & ~x[43] & ~x[44]) | (~x[39] & x[40] & x[41] & x[42] & ~x[44]) | (x[39] & x[40] & x[41] & ~x[43]) | (x[39] & x[41] & x[42] & ~x[43]) | (x[38] & x[40] & ~x[42] & x[43]);
  assign t[81] = (x[39] & ~x[40] & x[41] & ~x[42] & x[43]) | (x[39] & ~x[40] & x[41] & ~x[42] & x[44]) | (x[39] & ~x[40] & ~x[42] & x[43] & x[44]) | (x[38] & x[40] & x[41] & x[42] & x[43]) | (x[38] & ~x[40] & x[41] & x[44]) | (x[38] & ~x[42] & x[43] & x[44]) | (x[41] & x[43] & x[44]);
  assign t[8] = t[14] & t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind197(x, y);
 input [50:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[18] ^ t[19];
  assign t[11] = ~t[20];
  assign t[12] = t[21] ^ t[22];
  assign t[13] = t[23] & t[24];
  assign t[14] = t[25] ^ t[13];
  assign t[15] = t[56] ^ t[23];
  assign t[16] = t[26] ^ t[27];
  assign t[17] = t[28] & t[29];
  assign t[18] = t[30] ^ t[17];
  assign t[19] = t[57] ^ t[28];
  assign t[1] = ~(t[3] ^ t[54]);
  assign t[20] = ~(t[31] ^ t[32]);
  assign t[21] = t[58] ^ t[59];
  assign t[22] = t[23] & t[33];
  assign t[23] = ~(t[59]);
  assign t[24] = ~(t[56] ^ t[23]);
  assign t[25] = t[56] & t[34];
  assign t[26] = t[60] ^ t[61];
  assign t[27] = t[28] & t[35];
  assign t[28] = ~(t[61]);
  assign t[29] = ~(t[57] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[57] & t[36];
  assign t[31] = t[37] ^ t[38];
  assign t[32] = t[39] ^ t[40];
  assign t[33] = t[56] ^ t[41];
  assign t[34] = t[42] ^ t[22];
  assign t[35] = t[57] ^ t[43];
  assign t[36] = t[44] ^ t[27];
  assign t[37] = t[45] ^ t[46];
  assign t[38] = t[47] & t[48];
  assign t[39] = t[49] ^ t[38];
  assign t[3] = ~t[6];
  assign t[40] = t[62] ^ t[47];
  assign t[41] = t[59] ^ t[63];
  assign t[42] = t[56] ^ t[21];
  assign t[43] = t[61] ^ t[64];
  assign t[44] = t[57] ^ t[26];
  assign t[45] = t[65] ^ t[66];
  assign t[46] = t[47] & t[50];
  assign t[47] = ~(t[66]);
  assign t[48] = ~(t[62] ^ t[47]);
  assign t[49] = t[62] & t[51];
  assign t[4] = ~(t[7] ^ t[8]);
  assign t[50] = t[62] ^ t[52];
  assign t[51] = t[53] ^ t[46];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[62] ^ t[45];
  assign t[54] = t[68] ^ x[9];
  assign t[55] = t[69] ^ x[17];
  assign t[56] = t[70] ^ x[25];
  assign t[57] = t[71] ^ x[33];
  assign t[58] = t[72] ^ x[34];
  assign t[59] = t[73] ^ x[35];
  assign t[5] = ~(t[9] ^ t[10]);
  assign t[60] = t[74] ^ x[36];
  assign t[61] = t[75] ^ x[37];
  assign t[62] = t[76] ^ x[45];
  assign t[63] = t[77] ^ x[46];
  assign t[64] = t[78] ^ x[47];
  assign t[65] = t[79] ^ x[48];
  assign t[66] = t[80] ^ x[49];
  assign t[67] = t[81] ^ x[50];
  assign t[68] = (x[2] & x[3] & ~x[5] & x[6] & ~x[8]) | (~x[3] & x[4] & x[5] & x[6] & ~x[8]) | (x[2] & x[3] & ~x[4] & x[7] & ~x[8]) | (x[2] & ~x[5] & x[6] & x[7] & ~x[8]) | (x[2] & ~x[4] & x[5] & x[6]) | (x[3] & x[4] & ~x[5] & x[7]) | (x[3] & ~x[5] & x[6] & x[7]);
  assign t[69] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[6] = ~(t[11] ^ t[55]);
  assign t[70] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[71] = (x[26] & x[27] & ~x[29] & x[30] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[26] & x[27] & ~x[28] & x[31] & ~x[32]) | (x[26] & ~x[29] & x[30] & x[31] & ~x[32]) | (x[26] & ~x[28] & x[29] & x[30]) | (x[27] & x[28] & ~x[29] & x[31]) | (x[27] & ~x[29] & x[30] & x[31]);
  assign t[72] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[73] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[74] = (x[26] & x[27] & x[28] & ~x[31] & ~x[32]) | (x[26] & x[27] & x[29] & ~x[30] & ~x[32]) | (x[26] & x[28] & x[29] & ~x[31] & ~x[32]) | (~x[27] & x[28] & x[29] & x[30] & ~x[32]) | (x[27] & x[28] & x[29] & ~x[31]) | (x[27] & x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[30] & x[31]);
  assign t[75] = (x[26] & x[28] & ~x[29] & x[30] & ~x[31]) | (x[26] & x[28] & ~x[29] & ~x[31] & x[32]) | (x[26] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[27] & x[28] & ~x[29] & x[32]) | (x[27] & x[30] & ~x[31] & x[32]) | (x[28] & x[30] & x[32]);
  assign t[76] = (x[38] & x[39] & ~x[41] & x[42] & ~x[44]) | (~x[39] & x[40] & x[41] & x[42] & ~x[44]) | (x[38] & x[39] & ~x[40] & x[43] & ~x[44]) | (x[38] & ~x[41] & x[42] & x[43] & ~x[44]) | (x[38] & ~x[40] & x[41] & x[42]) | (x[39] & x[40] & ~x[41] & x[43]) | (x[39] & ~x[41] & x[42] & x[43]);
  assign t[77] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[78] = (x[27] & ~x[28] & x[29] & ~x[30] & x[31]) | (x[27] & ~x[28] & x[29] & ~x[30] & x[32]) | (x[27] & ~x[28] & ~x[30] & x[31] & x[32]) | (x[26] & x[28] & x[29] & x[30] & x[31]) | (x[26] & ~x[28] & x[29] & x[32]) | (x[26] & ~x[30] & x[31] & x[32]) | (x[29] & x[31] & x[32]);
  assign t[79] = (x[38] & x[39] & x[40] & ~x[43] & ~x[44]) | (x[38] & x[39] & x[41] & ~x[42] & ~x[44]) | (x[38] & x[40] & x[41] & ~x[43] & ~x[44]) | (~x[39] & x[40] & x[41] & x[42] & ~x[44]) | (x[39] & x[40] & x[41] & ~x[43]) | (x[39] & x[41] & x[42] & ~x[43]) | (x[38] & x[40] & ~x[42] & x[43]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[38] & x[40] & ~x[41] & x[42] & ~x[43]) | (x[38] & x[40] & ~x[41] & ~x[43] & x[44]) | (x[38] & ~x[41] & x[42] & ~x[43] & x[44]) | (x[38] & x[40] & x[41] & x[42] & x[43]) | (x[39] & x[40] & ~x[41] & x[44]) | (x[39] & x[42] & ~x[43] & x[44]) | (x[40] & x[42] & x[44]);
  assign t[81] = (x[39] & ~x[40] & x[41] & ~x[42] & x[43]) | (x[39] & ~x[40] & x[41] & ~x[42] & x[44]) | (x[39] & ~x[40] & ~x[42] & x[43] & x[44]) | (x[38] & x[40] & x[41] & x[42] & x[43]) | (x[38] & ~x[40] & x[41] & x[44]) | (x[38] & ~x[42] & x[43] & x[44]) | (x[41] & x[43] & x[44]);
  assign t[8] = t[14] ^ t[15];
  assign t[9] = t[16] ^ t[17];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind198(x, y);
 input [47:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[15] & t[16];
  assign t[12] = t[28] ^ t[29];
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[19]);
  assign t[15] = ~(t[26]);
  assign t[16] = ~(t[30] ^ t[15]);
  assign t[17] = ~(t[28]);
  assign t[18] = ~(t[31] ^ t[17]);
  assign t[19] = t[20] ^ t[21];
  assign t[1] = ~(t[3] ^ t[24]);
  assign t[20] = t[32] ^ t[33];
  assign t[21] = t[22] & t[23];
  assign t[22] = ~(t[32]);
  assign t[23] = ~(t[34] ^ t[22]);
  assign t[24] = t[35] ^ x[9];
  assign t[25] = t[36] ^ x[17];
  assign t[26] = t[37] ^ x[25];
  assign t[27] = t[38] ^ x[26];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[35];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[41] ^ x[36];
  assign t[31] = t[42] ^ x[37];
  assign t[32] = t[43] ^ x[45];
  assign t[33] = t[44] ^ x[46];
  assign t[34] = t[45] ^ x[47];
  assign t[35] = (x[2] & x[4] & ~x[5] & x[6] & ~x[7]) | (x[2] & x[4] & ~x[5] & ~x[7] & x[8]) | (x[2] & ~x[5] & x[6] & ~x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[3] & x[4] & ~x[5] & x[8]) | (x[3] & x[6] & ~x[7] & x[8]) | (x[4] & x[6] & x[8]);
  assign t[36] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[37] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[38] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[39] = (x[27] & x[29] & ~x[30] & x[31] & ~x[32]) | (x[27] & x[29] & ~x[30] & ~x[32] & x[33]) | (x[27] & ~x[30] & x[31] & ~x[32] & x[33]) | (x[27] & x[29] & x[30] & x[31] & x[32]) | (x[28] & x[29] & ~x[30] & x[33]) | (x[28] & x[31] & ~x[32] & x[33]) | (x[29] & x[31] & x[33]);
  assign t[3] = ~t[6];
  assign t[40] = (x[28] & ~x[29] & x[30] & ~x[31] & x[32]) | (x[28] & ~x[29] & x[30] & ~x[31] & x[33]) | (x[28] & ~x[29] & ~x[31] & x[32] & x[33]) | (x[27] & x[29] & x[30] & x[31] & x[32]) | (x[27] & ~x[29] & x[30] & x[33]) | (x[27] & ~x[31] & x[32] & x[33]) | (x[30] & x[32] & x[33]);
  assign t[41] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[42] = (x[27] & x[28] & ~x[30] & x[31] & ~x[33]) | (~x[28] & x[29] & x[30] & x[31] & ~x[33]) | (x[27] & x[28] & ~x[29] & x[32] & ~x[33]) | (x[27] & ~x[30] & x[31] & x[32] & ~x[33]) | (x[27] & ~x[29] & x[30] & x[31]) | (x[28] & x[29] & ~x[30] & x[32]) | (x[28] & ~x[30] & x[31] & x[32]);
  assign t[43] = (x[38] & x[40] & ~x[41] & x[42] & ~x[43]) | (x[38] & x[40] & ~x[41] & ~x[43] & x[44]) | (x[38] & ~x[41] & x[42] & ~x[43] & x[44]) | (x[38] & x[40] & x[41] & x[42] & x[43]) | (x[39] & x[40] & ~x[41] & x[44]) | (x[39] & x[42] & ~x[43] & x[44]) | (x[40] & x[42] & x[44]);
  assign t[44] = (x[39] & ~x[40] & x[41] & ~x[42] & x[43]) | (x[39] & ~x[40] & x[41] & ~x[42] & x[44]) | (x[39] & ~x[40] & ~x[42] & x[43] & x[44]) | (x[38] & x[40] & x[41] & x[42] & x[43]) | (x[38] & ~x[40] & x[41] & x[44]) | (x[38] & ~x[42] & x[43] & x[44]) | (x[41] & x[43] & x[44]);
  assign t[45] = (x[38] & x[39] & ~x[41] & x[42] & ~x[44]) | (~x[39] & x[40] & x[41] & x[42] & ~x[44]) | (x[38] & x[39] & ~x[40] & x[43] & ~x[44]) | (x[38] & ~x[41] & x[42] & x[43] & ~x[44]) | (x[38] & ~x[40] & x[41] & x[42]) | (x[39] & x[40] & ~x[41] & x[43]) | (x[39] & ~x[41] & x[42] & x[43]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9] ^ t[25]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~t[14];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1ind199(x, y);
 input [50:0] x;
 output y;

 wire [63:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[15] ^ t[16];
  assign t[11] = t[17] & t[18];
  assign t[12] = t[19] ^ t[20];
  assign t[13] = t[21] & t[22];
  assign t[14] = ~(t[23]);
  assign t[15] = t[38] ^ t[39];
  assign t[16] = t[17] & t[24];
  assign t[17] = ~(t[39]);
  assign t[18] = ~(t[40] ^ t[17]);
  assign t[19] = t[41] ^ t[42];
  assign t[1] = ~(t[3] ^ t[36]);
  assign t[20] = t[21] & t[25];
  assign t[21] = ~(t[42]);
  assign t[22] = ~(t[43] ^ t[21]);
  assign t[23] = t[26] ^ t[27];
  assign t[24] = t[40] ^ t[28];
  assign t[25] = t[43] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[39] ^ t[44];
  assign t[29] = t[42] ^ t[45];
  assign t[2] = ~(t[4] ^ t[5]);
  assign t[30] = t[46] ^ t[47];
  assign t[31] = t[32] & t[34];
  assign t[32] = ~(t[47]);
  assign t[33] = ~(t[48] ^ t[32]);
  assign t[34] = t[48] ^ t[35];
  assign t[35] = t[47] ^ t[49];
  assign t[36] = t[50] ^ x[9];
  assign t[37] = t[51] ^ x[17];
  assign t[38] = t[52] ^ x[25];
  assign t[39] = t[53] ^ x[26];
  assign t[3] = ~t[6];
  assign t[40] = t[54] ^ x[27];
  assign t[41] = t[55] ^ x[35];
  assign t[42] = t[56] ^ x[36];
  assign t[43] = t[57] ^ x[37];
  assign t[44] = t[58] ^ x[38];
  assign t[45] = t[59] ^ x[39];
  assign t[46] = t[60] ^ x[47];
  assign t[47] = t[61] ^ x[48];
  assign t[48] = t[62] ^ x[49];
  assign t[49] = t[63] ^ x[50];
  assign t[4] = ~(t[7]);
  assign t[50] = (x[3] & ~x[4] & x[5] & ~x[6] & x[7]) | (x[3] & ~x[4] & x[5] & ~x[6] & x[8]) | (x[3] & ~x[4] & ~x[6] & x[7] & x[8]) | (x[2] & x[4] & x[5] & x[6] & x[7]) | (x[2] & ~x[4] & x[5] & x[8]) | (x[2] & ~x[6] & x[7] & x[8]) | (x[5] & x[7] & x[8]);
  assign t[51] = (x[10] & x[11] & x[12] & ~x[15] & ~x[16]) | (x[10] & x[11] & x[13] & ~x[14] & ~x[16]) | (x[10] & x[12] & x[13] & ~x[15] & ~x[16]) | (~x[11] & x[12] & x[13] & x[14] & ~x[16]) | (x[11] & x[12] & x[13] & ~x[15]) | (x[11] & x[13] & x[14] & ~x[15]) | (x[10] & x[12] & ~x[14] & x[15]);
  assign t[52] = (x[18] & x[19] & x[20] & ~x[23] & ~x[24]) | (x[18] & x[19] & x[21] & ~x[22] & ~x[24]) | (x[18] & x[20] & x[21] & ~x[23] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[19] & x[20] & x[21] & ~x[23]) | (x[19] & x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[22] & x[23]);
  assign t[53] = (x[18] & x[20] & ~x[21] & x[22] & ~x[23]) | (x[18] & x[20] & ~x[21] & ~x[23] & x[24]) | (x[18] & ~x[21] & x[22] & ~x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[19] & x[20] & ~x[21] & x[24]) | (x[19] & x[22] & ~x[23] & x[24]) | (x[20] & x[22] & x[24]);
  assign t[54] = (x[18] & x[19] & ~x[21] & x[22] & ~x[24]) | (~x[19] & x[20] & x[21] & x[22] & ~x[24]) | (x[18] & x[19] & ~x[20] & x[23] & ~x[24]) | (x[18] & ~x[21] & x[22] & x[23] & ~x[24]) | (x[18] & ~x[20] & x[21] & x[22]) | (x[19] & x[20] & ~x[21] & x[23]) | (x[19] & ~x[21] & x[22] & x[23]);
  assign t[55] = (x[28] & x[29] & x[30] & ~x[33] & ~x[34]) | (x[28] & x[29] & x[31] & ~x[32] & ~x[34]) | (x[28] & x[30] & x[31] & ~x[33] & ~x[34]) | (~x[29] & x[30] & x[31] & x[32] & ~x[34]) | (x[29] & x[30] & x[31] & ~x[33]) | (x[29] & x[31] & x[32] & ~x[33]) | (x[28] & x[30] & ~x[32] & x[33]);
  assign t[56] = (x[28] & x[30] & ~x[31] & x[32] & ~x[33]) | (x[28] & x[30] & ~x[31] & ~x[33] & x[34]) | (x[28] & ~x[31] & x[32] & ~x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[29] & x[30] & ~x[31] & x[34]) | (x[29] & x[32] & ~x[33] & x[34]) | (x[30] & x[32] & x[34]);
  assign t[57] = (x[28] & x[29] & ~x[31] & x[32] & ~x[34]) | (~x[29] & x[30] & x[31] & x[32] & ~x[34]) | (x[28] & x[29] & ~x[30] & x[33] & ~x[34]) | (x[28] & ~x[31] & x[32] & x[33] & ~x[34]) | (x[28] & ~x[30] & x[31] & x[32]) | (x[29] & x[30] & ~x[31] & x[33]) | (x[29] & ~x[31] & x[32] & x[33]);
  assign t[58] = (x[19] & ~x[20] & x[21] & ~x[22] & x[23]) | (x[19] & ~x[20] & x[21] & ~x[22] & x[24]) | (x[19] & ~x[20] & ~x[22] & x[23] & x[24]) | (x[18] & x[20] & x[21] & x[22] & x[23]) | (x[18] & ~x[20] & x[21] & x[24]) | (x[18] & ~x[22] & x[23] & x[24]) | (x[21] & x[23] & x[24]);
  assign t[59] = (x[29] & ~x[30] & x[31] & ~x[32] & x[33]) | (x[29] & ~x[30] & x[31] & ~x[32] & x[34]) | (x[29] & ~x[30] & ~x[32] & x[33] & x[34]) | (x[28] & x[30] & x[31] & x[32] & x[33]) | (x[28] & ~x[30] & x[31] & x[34]) | (x[28] & ~x[32] & x[33] & x[34]) | (x[31] & x[33] & x[34]);
  assign t[5] = ~(t[8]);
  assign t[60] = (x[40] & x[41] & x[42] & ~x[45] & ~x[46]) | (x[40] & x[41] & x[43] & ~x[44] & ~x[46]) | (x[40] & x[42] & x[43] & ~x[45] & ~x[46]) | (~x[41] & x[42] & x[43] & x[44] & ~x[46]) | (x[41] & x[42] & x[43] & ~x[45]) | (x[41] & x[43] & x[44] & ~x[45]) | (x[40] & x[42] & ~x[44] & x[45]);
  assign t[61] = (x[40] & x[42] & ~x[43] & x[44] & ~x[45]) | (x[40] & x[42] & ~x[43] & ~x[45] & x[46]) | (x[40] & ~x[43] & x[44] & ~x[45] & x[46]) | (x[40] & x[42] & x[43] & x[44] & x[45]) | (x[41] & x[42] & ~x[43] & x[46]) | (x[41] & x[44] & ~x[45] & x[46]) | (x[42] & x[44] & x[46]);
  assign t[62] = (x[40] & x[41] & ~x[43] & x[44] & ~x[46]) | (~x[41] & x[42] & x[43] & x[44] & ~x[46]) | (x[40] & x[41] & ~x[42] & x[45] & ~x[46]) | (x[40] & ~x[43] & x[44] & x[45] & ~x[46]) | (x[40] & ~x[42] & x[43] & x[44]) | (x[41] & x[42] & ~x[43] & x[45]) | (x[41] & ~x[43] & x[44] & x[45]);
  assign t[63] = (x[41] & ~x[42] & x[43] & ~x[44] & x[45]) | (x[41] & ~x[42] & x[43] & ~x[44] & x[46]) | (x[41] & ~x[42] & ~x[44] & x[45] & x[46]) | (x[40] & x[42] & x[43] & x[44] & x[45]) | (x[40] & ~x[42] & x[43] & x[46]) | (x[40] & ~x[44] & x[45] & x[46]) | (x[43] & x[45] & x[46]);
  assign t[6] = ~(t[9] ^ t[37]);
  assign t[7] = t[10] ^ t[11];
  assign t[8] = t[12] ^ t[13];
  assign t[9] = ~t[14];
  assign y = x[0] ? x[1] : t[0];
endmodule

module R1_ind(x, y);
 input [536:0] x;
 output [199:0] y;

  R1ind0 R1ind0_inst(.x({x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[17], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[28], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[29], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[39], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[40], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[50], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[51], x[47], x[46], x[45], x[44], x[43], x[42], x[41]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[61], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[58], x[57], x[56], x[55], x[54], x[53], x[52]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[72], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[73], x[69], x[68], x[67], x[66], x[65], x[64], x[63]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[84], x[80], x[79], x[78], x[77], x[76], x[75], x[74]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[94], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[95], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[105], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[106], x[102], x[101], x[100], x[99], x[98], x[97], x[96]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[116], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[117], x[113], x[112], x[111], x[110], x[109], x[108], x[107]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[127], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[128], x[124], x[123], x[122], x[121], x[120], x[119], x[118]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[138], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[139], x[135], x[134], x[133], x[132], x[131], x[130], x[129]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[150], x[146], x[145], x[144], x[143], x[142], x[141], x[140]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[161], x[157], x[156], x[155], x[154], x[153], x[152], x[151]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[172], x[168], x[167], x[166], x[165], x[164], x[163], x[162]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[183], x[179], x[178], x[177], x[176], x[175], x[174], x[173]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[232]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[232]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[232]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[232]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[232]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[232]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[243], x[242], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[245], x[244], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[247], x[246], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[232]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[258], x[257], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[232]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[260], x[259], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[232]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[262], x[261], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[232]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[232]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[273], x[272], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[232]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[275], x[274], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[232]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[277], x[276], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[232]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[232]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[288], x[287], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[232]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[290], x[289], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[232]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[292], x[291], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[232]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[232]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[303], x[302], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[232]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[305], x[304], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[232]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[307], x[306], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[232]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[232]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[318], x[317], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[232]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[320], x[319], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[232]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[322], x[321], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[232]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[232]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[333], x[332], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[232]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[335], x[334], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[232]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[337], x[336], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[232]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[346], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[232]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[348], x[347], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[232]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[350], x[349], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[232]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[352], x[351], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[232]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[361], x[360], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[232]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[363], x[362], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[232]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[365], x[364], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[232]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[367], x[366], x[359], x[358], x[357], x[356], x[355], x[354], x[353], x[232]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[376], x[375], x[374], x[373], x[372], x[371], x[370], x[369], x[368], x[232]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[378], x[377], x[374], x[373], x[372], x[371], x[370], x[369], x[368], x[232]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[380], x[379], x[374], x[373], x[372], x[371], x[370], x[369], x[368], x[232]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[382], x[381], x[374], x[373], x[372], x[371], x[370], x[369], x[368], x[232]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[391], x[390], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[232]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[393], x[392], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[232]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[395], x[394], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[232]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[397], x[396], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[232]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[232]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[408], x[407], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[232]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[410], x[409], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[232]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[232]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[232]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[423], x[422], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[232]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[425], x[424], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[232]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[427], x[426], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[232]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[436], x[435], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[232]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[438], x[437], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[232]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[440], x[439], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[232]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[442], x[441], x[434], x[433], x[432], x[431], x[430], x[429], x[428], x[232]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[451], x[450], x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[232]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[453], x[452], x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[232]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[455], x[454], x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[232]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[457], x[456], x[449], x[448], x[447], x[446], x[445], x[444], x[443], x[232]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[232]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[468], x[467], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[232]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[470], x[469], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[232]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[472], x[471], x[464], x[463], x[462], x[461], x[460], x[459], x[458], x[232]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[150], x[147], x[149], x[84], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[81], x[83], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[473], x[232]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[150], x[149], x[147], x[84], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[83], x[81], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[302], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[474], x[232]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[148], x[150], x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[82], x[84], x[83], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[304], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[475], x[232]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[150], x[148], x[149], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[84], x[82], x[83], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[306], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[476], x[232]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[161], x[158], x[160], x[95], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[92], x[94], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[477], x[232]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[161], x[95], x[160], x[158], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[94], x[92], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[317], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[478], x[232]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[159], x[161], x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[93], x[95], x[94], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[319], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[479], x[232]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[161], x[159], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[95], x[93], x[94], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[321], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[480], x[232]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[172], x[169], x[171], x[62], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[59], x[61], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[481], x[232]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[172], x[171], x[169], x[62], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[61], x[59], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[332], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[482], x[232]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[170], x[172], x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[60], x[62], x[61], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[334], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[483], x[232]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[172], x[170], x[171], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[62], x[60], x[61], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[336], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[484], x[232]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[183], x[180], x[182], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[73], x[70], x[72], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[485], x[232]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[183], x[182], x[180], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[73], x[72], x[70], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[347], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[486], x[232]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[181], x[183], x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[71], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[73], x[72], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[349], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[487], x[232]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[183], x[181], x[182], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[73], x[71], x[72], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[351], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[488], x[232]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[117], x[114], x[116], x[84], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[81], x[83], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[489], x[232]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[117], x[116], x[114], x[84], x[115], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[83], x[81], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[257], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[490], x[232]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[115], x[117], x[116], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[82], x[84], x[83], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[259], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[491], x[232]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[117], x[115], x[116], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[84], x[82], x[83], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[261], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[492], x[232]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[128], x[125], x[127], x[95], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[92], x[94], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[493], x[232]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[128], x[95], x[127], x[125], x[126], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[94], x[92], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[272], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[494], x[232]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[126], x[128], x[127], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[93], x[95], x[94], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[274], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[495], x[232]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[128], x[126], x[127], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[95], x[93], x[94], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[276], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[496], x[232]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[139], x[136], x[138], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[62], x[59], x[61], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[497], x[232]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[139], x[138], x[136], x[137], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[62], x[61], x[59], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[287], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[498], x[232]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[137], x[139], x[138], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[60], x[62], x[61], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[289], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[499], x[232]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[139], x[137], x[138], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[62], x[60], x[61], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[291], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[500], x[232]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[106], x[103], x[105], x[73], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[70], x[72], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[501], x[232]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[106], x[105], x[103], x[73], x[104], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[72], x[70], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[242], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[502], x[232]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[104], x[106], x[105], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[71], x[73], x[72], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[244], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[503], x[232]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[106], x[104], x[105], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[73], x[71], x[72], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[246], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[504], x[232]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[150], x[147], x[149], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[505], x[232]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[150], x[149], x[147], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[302], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[506], x[232]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[148], x[150], x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[304], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[507], x[232]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[150], x[148], x[149], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[306], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[508], x[232]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[161], x[158], x[160], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[509], x[232]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[161], x[160], x[158], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[317], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[510], x[232]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[159], x[161], x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[319], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[511], x[232]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[161], x[159], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[321], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[512], x[232]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[172], x[169], x[171], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[513], x[232]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[172], x[171], x[169], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[332], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[514], x[232]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[170], x[172], x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[334], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[515], x[232]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[172], x[170], x[171], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[336], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[516], x[232]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[183], x[180], x[182], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[517], x[232]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[183], x[182], x[180], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[347], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[518], x[232]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[181], x[183], x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[349], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[519], x[232]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[183], x[181], x[182], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[351], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[520], x[232]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[150], x[51], x[84], x[147], x[149], x[48], x[50], x[81], x[83], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[521], x[232]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[150], x[51], x[84], x[149], x[147], x[50], x[48], x[83], x[81], x[148], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[49], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[82], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[302], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[522], x[232]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[148], x[49], x[82], x[150], x[149], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[51], x[50], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[84], x[83], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[304], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[523], x[232]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[150], x[51], x[84], x[148], x[149], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[49], x[50], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[82], x[83], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[306], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[524], x[232]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[161], x[18], x[95], x[158], x[160], x[15], x[17], x[92], x[94], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[525], x[232]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[95], x[161], x[18], x[94], x[92], x[160], x[158], x[17], x[15], x[93], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[159], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[16], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[317], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[526], x[232]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[159], x[16], x[93], x[161], x[160], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[18], x[17], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[95], x[94], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[319], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[527], x[232]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[161], x[18], x[95], x[159], x[160], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[16], x[17], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[93], x[94], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[321], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[528], x[232]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[172], x[29], x[62], x[169], x[171], x[26], x[28], x[59], x[61], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[529], x[232]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[172], x[29], x[62], x[171], x[169], x[28], x[26], x[61], x[59], x[170], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[27], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[60], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[332], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[530], x[232]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[170], x[27], x[60], x[172], x[171], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[29], x[28], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[62], x[61], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[334], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[531], x[232]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[172], x[29], x[62], x[170], x[171], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[27], x[28], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[60], x[61], x[59], x[58], x[57], x[56], x[55], x[54], x[53], x[52], x[336], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[532], x[232]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[183], x[180], x[182], x[40], x[73], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[37], x[39], x[70], x[72], x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[533], x[232]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[183], x[182], x[180], x[40], x[73], x[181], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[39], x[37], x[72], x[70], x[38], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[71], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[347], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[534], x[232]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[181], x[183], x[182], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[38], x[71], x[40], x[39], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[73], x[72], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[349], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[535], x[232]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[183], x[181], x[182], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[40], x[73], x[38], x[39], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[71], x[72], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[351], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[536], x[232]}), .y(y[199]));
endmodule

module R2ind0(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[4] & ~t[5] & ~t[6] & ~t[7]) | (t[2] & ~t[3] & ~t[5] & ~t[6] & ~t[8]) | (t[2] & ~t[3] & ~t[4] & ~t[7] & ~t[8]) | (~t[2] & t[3] & t[4] & t[5] & ~t[8]) | (~t[2] & t[3] & t[6] & t[7] & ~t[8]) | (t[2] & ~t[4] & ~t[6] & t[8]) | (~t[2] & t[4] & t[6] & t[8]);
  assign t[2] = t[9] ^ x[7];
  assign t[3] = t[10] ^ x[1];
  assign t[4] = t[11] ^ x[2];
  assign t[5] = t[12] ^ x[3];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[3] & ~t[4] & ~t[5] & ~t[6] & ~t[7]) | (~t[2] & t[3] & ~t[5] & ~t[6] & ~t[8]) | (~t[2] & t[3] & ~t[4] & ~t[7] & ~t[8]) | (t[2] & ~t[3] & t[4] & t[5] & ~t[8]) | (t[2] & ~t[3] & t[6] & t[7] & ~t[8]) | (t[3] & ~t[5] & ~t[7] & t[8]) | (~t[3] & t[5] & t[7] & t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[7];
  assign t[4] = t[11] ^ x[2];
  assign t[5] = t[12] ^ x[3];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & ~t[4] & t[5] & ~t[6] & ~t[8]) | (t[2] & ~t[4] & ~t[5] & t[6] & ~t[7] & t[8]) | (~t[3] & t[4] & ~t[5] & ~t[6] & ~t[8]) | (~t[2] & t[4] & ~t[5] & ~t[6] & ~t[7]) | (~t[2] & ~t[3] & t[4] & ~t[7] & ~t[8]) | (~t[2] & t[4] & t[5] & ~t[6] & t[7]) | (t[4] & ~t[5] & t[7] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[7];
  assign t[5] = t[12] ^ x[3];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & t[4] & ~t[5] & ~t[7] & ~t[8]) | (t[3] & ~t[4] & ~t[5] & ~t[6] & t[7] & t[8]) | (~t[3] & ~t[4] & t[5] & ~t[6] & ~t[7]) | (~t[2] & ~t[4] & t[5] & ~t[7] & ~t[8]) | (~t[2] & ~t[3] & t[5] & ~t[6] & ~t[8]) | (~t[3] & t[4] & t[5] & t[6] & ~t[7]) | (~t[4] & t[5] & t[6] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[7];
  assign t[6] = t[13] ^ x[4];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & ~t[4] & ~t[6] & t[7] & ~t[8]) | (t[2] & t[4] & ~t[5] & ~t[6] & ~t[7] & t[8]) | (~t[3] & ~t[4] & t[6] & ~t[7] & ~t[8]) | (~t[2] & ~t[4] & ~t[5] & t[6] & ~t[7]) | (~t[2] & ~t[3] & ~t[5] & t[6] & ~t[8]) | (~t[2] & ~t[4] & t[5] & t[6] & t[7]) | (t[5] & t[6] & ~t[7] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[4];
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[5];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[3] & ~t[5] & t[6] & ~t[7] & ~t[8]) | (t[3] & ~t[4] & t[5] & ~t[6] & ~t[7] & t[8]) | (~t[3] & ~t[4] & ~t[5] & ~t[6] & t[7]) | (~t[2] & ~t[5] & ~t[6] & t[7] & ~t[8]) | (~t[2] & ~t[3] & ~t[4] & t[7] & ~t[8]) | (~t[3] & t[4] & ~t[5] & t[6] & t[7]) | (t[4] & ~t[6] & t[7] & ~t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[4];
  assign t[6] = t[13] ^ x[5];
  assign t[7] = t[14] ^ x[7];
  assign t[8] = t[15] ^ x[6];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind6(x, y);
 input [7:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ x[7];
  assign t[10] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[11] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[12] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[13] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & t[4] & ~t[5] & t[6] & ~t[7] & ~t[8]) | (t[3] & ~t[4] & t[5] & ~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[5] & ~t[6] & ~t[7] & t[8]) | (~t[2] & ~t[3] & ~t[6] & ~t[7] & t[8]) | (~t[2] & ~t[3] & ~t[4] & ~t[5] & t[8]) | (t[2] & t[3] & ~t[6] & ~t[7] & t[8]) | (t[2] & t[3] & ~t[4] & ~t[5] & t[8]);
  assign t[2] = t[9] ^ x[1];
  assign t[3] = t[10] ^ x[2];
  assign t[4] = t[11] ^ x[3];
  assign t[5] = t[12] ^ x[4];
  assign t[6] = t[13] ^ x[5];
  assign t[7] = t[14] ^ x[6];
  assign t[8] = t[15] ^ x[7];
  assign t[9] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign y = t[0];
endmodule

module R2ind7(x, y);
 input [47:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[101] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[102] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[107] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[108] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[109] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[114] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[115] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[116] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[6];
  assign t[13] = t[25] ^ x[7];
  assign t[14] = t[26] ^ x[14];
  assign t[15] = t[27] ^ x[15];
  assign t[16] = t[28] ^ x[22];
  assign t[17] = t[29] ^ x[23];
  assign t[18] = t[30] ^ x[30];
  assign t[19] = t[31] ^ x[31];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[32] ^ x[38];
  assign t[21] = t[33] ^ x[39];
  assign t[22] = t[34] ^ x[46];
  assign t[23] = t[35] ^ x[47];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[6];
  assign t[37] = t[79] ^ x[1];
  assign t[38] = t[80] ^ x[2];
  assign t[39] = t[81] ^ x[3];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[82] ^ x[7];
  assign t[41] = t[83] ^ x[4];
  assign t[42] = t[84] ^ x[5];
  assign t[43] = t[85] ^ x[14];
  assign t[44] = t[86] ^ x[9];
  assign t[45] = t[87] ^ x[10];
  assign t[46] = t[88] ^ x[11];
  assign t[47] = t[89] ^ x[15];
  assign t[48] = t[90] ^ x[12];
  assign t[49] = t[91] ^ x[13];
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = t[92] ^ x[22];
  assign t[51] = t[93] ^ x[17];
  assign t[52] = t[94] ^ x[18];
  assign t[53] = t[95] ^ x[19];
  assign t[54] = t[96] ^ x[23];
  assign t[55] = t[97] ^ x[20];
  assign t[56] = t[98] ^ x[21];
  assign t[57] = t[99] ^ x[30];
  assign t[58] = t[100] ^ x[25];
  assign t[59] = t[101] ^ x[26];
  assign t[5] = ~(t[11]);
  assign t[60] = t[102] ^ x[27];
  assign t[61] = t[103] ^ x[31];
  assign t[62] = t[104] ^ x[28];
  assign t[63] = t[105] ^ x[29];
  assign t[64] = t[106] ^ x[38];
  assign t[65] = t[107] ^ x[33];
  assign t[66] = t[108] ^ x[34];
  assign t[67] = t[109] ^ x[35];
  assign t[68] = t[110] ^ x[39];
  assign t[69] = t[111] ^ x[36];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[37];
  assign t[71] = t[113] ^ x[46];
  assign t[72] = t[114] ^ x[41];
  assign t[73] = t[115] ^ x[42];
  assign t[74] = t[116] ^ x[43];
  assign t[75] = t[117] ^ x[47];
  assign t[76] = t[118] ^ x[44];
  assign t[77] = t[119] ^ x[45];
  assign t[78] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[79] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[81] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[86] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[87] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[88] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[93] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[94] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[95] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind8(x, y);
 input [47:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[101] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[102] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[107] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[108] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[109] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[114] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[115] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[116] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[6];
  assign t[13] = t[25] ^ x[7];
  assign t[14] = t[26] ^ x[14];
  assign t[15] = t[27] ^ x[15];
  assign t[16] = t[28] ^ x[22];
  assign t[17] = t[29] ^ x[23];
  assign t[18] = t[30] ^ x[30];
  assign t[19] = t[31] ^ x[31];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[32] ^ x[38];
  assign t[21] = t[33] ^ x[39];
  assign t[22] = t[34] ^ x[46];
  assign t[23] = t[35] ^ x[47];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[6];
  assign t[37] = t[79] ^ x[1];
  assign t[38] = t[80] ^ x[2];
  assign t[39] = t[81] ^ x[3];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[82] ^ x[7];
  assign t[41] = t[83] ^ x[4];
  assign t[42] = t[84] ^ x[5];
  assign t[43] = t[85] ^ x[14];
  assign t[44] = t[86] ^ x[9];
  assign t[45] = t[87] ^ x[10];
  assign t[46] = t[88] ^ x[11];
  assign t[47] = t[89] ^ x[15];
  assign t[48] = t[90] ^ x[12];
  assign t[49] = t[91] ^ x[13];
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = t[92] ^ x[22];
  assign t[51] = t[93] ^ x[17];
  assign t[52] = t[94] ^ x[18];
  assign t[53] = t[95] ^ x[19];
  assign t[54] = t[96] ^ x[23];
  assign t[55] = t[97] ^ x[20];
  assign t[56] = t[98] ^ x[21];
  assign t[57] = t[99] ^ x[30];
  assign t[58] = t[100] ^ x[25];
  assign t[59] = t[101] ^ x[26];
  assign t[5] = ~(t[11]);
  assign t[60] = t[102] ^ x[27];
  assign t[61] = t[103] ^ x[31];
  assign t[62] = t[104] ^ x[28];
  assign t[63] = t[105] ^ x[29];
  assign t[64] = t[106] ^ x[38];
  assign t[65] = t[107] ^ x[33];
  assign t[66] = t[108] ^ x[34];
  assign t[67] = t[109] ^ x[35];
  assign t[68] = t[110] ^ x[39];
  assign t[69] = t[111] ^ x[36];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[37];
  assign t[71] = t[113] ^ x[46];
  assign t[72] = t[114] ^ x[41];
  assign t[73] = t[115] ^ x[42];
  assign t[74] = t[116] ^ x[43];
  assign t[75] = t[117] ^ x[47];
  assign t[76] = t[118] ^ x[44];
  assign t[77] = t[119] ^ x[45];
  assign t[78] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[79] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[81] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[86] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[87] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[88] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[93] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[94] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[95] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind9(x, y);
 input [47:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[101] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[102] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[107] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[108] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[109] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[114] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[115] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[116] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[6];
  assign t[13] = t[25] ^ x[7];
  assign t[14] = t[26] ^ x[14];
  assign t[15] = t[27] ^ x[15];
  assign t[16] = t[28] ^ x[22];
  assign t[17] = t[29] ^ x[23];
  assign t[18] = t[30] ^ x[30];
  assign t[19] = t[31] ^ x[31];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[32] ^ x[38];
  assign t[21] = t[33] ^ x[39];
  assign t[22] = t[34] ^ x[46];
  assign t[23] = t[35] ^ x[47];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[6];
  assign t[37] = t[79] ^ x[1];
  assign t[38] = t[80] ^ x[2];
  assign t[39] = t[81] ^ x[3];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[82] ^ x[7];
  assign t[41] = t[83] ^ x[4];
  assign t[42] = t[84] ^ x[5];
  assign t[43] = t[85] ^ x[14];
  assign t[44] = t[86] ^ x[9];
  assign t[45] = t[87] ^ x[10];
  assign t[46] = t[88] ^ x[11];
  assign t[47] = t[89] ^ x[15];
  assign t[48] = t[90] ^ x[12];
  assign t[49] = t[91] ^ x[13];
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = t[92] ^ x[22];
  assign t[51] = t[93] ^ x[17];
  assign t[52] = t[94] ^ x[18];
  assign t[53] = t[95] ^ x[19];
  assign t[54] = t[96] ^ x[23];
  assign t[55] = t[97] ^ x[20];
  assign t[56] = t[98] ^ x[21];
  assign t[57] = t[99] ^ x[30];
  assign t[58] = t[100] ^ x[25];
  assign t[59] = t[101] ^ x[26];
  assign t[5] = ~(t[11]);
  assign t[60] = t[102] ^ x[27];
  assign t[61] = t[103] ^ x[31];
  assign t[62] = t[104] ^ x[28];
  assign t[63] = t[105] ^ x[29];
  assign t[64] = t[106] ^ x[38];
  assign t[65] = t[107] ^ x[33];
  assign t[66] = t[108] ^ x[34];
  assign t[67] = t[109] ^ x[35];
  assign t[68] = t[110] ^ x[39];
  assign t[69] = t[111] ^ x[36];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[37];
  assign t[71] = t[113] ^ x[46];
  assign t[72] = t[114] ^ x[41];
  assign t[73] = t[115] ^ x[42];
  assign t[74] = t[116] ^ x[43];
  assign t[75] = t[117] ^ x[47];
  assign t[76] = t[118] ^ x[44];
  assign t[77] = t[119] ^ x[45];
  assign t[78] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[79] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[81] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[86] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[87] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[88] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[93] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[94] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[95] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind10(x, y);
 input [47:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[101] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[102] = (x[24] & ~1'b0) | (~x[24] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[107] = (x[32] & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0);
  assign t[108] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[109] = (x[32] & ~1'b0) | (~x[32] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[114] = (x[40] & ~1'b0 & ~1'b0) | (~x[40] & 1'b0 & ~1'b0) | (~x[40] & ~1'b0 & 1'b0) | (x[40] & 1'b0 & 1'b0);
  assign t[115] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[116] = (x[40] & ~1'b0) | (~x[40] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[6];
  assign t[13] = t[25] ^ x[7];
  assign t[14] = t[26] ^ x[14];
  assign t[15] = t[27] ^ x[15];
  assign t[16] = t[28] ^ x[22];
  assign t[17] = t[29] ^ x[23];
  assign t[18] = t[30] ^ x[30];
  assign t[19] = t[31] ^ x[31];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[32] ^ x[38];
  assign t[21] = t[33] ^ x[39];
  assign t[22] = t[34] ^ x[46];
  assign t[23] = t[35] ^ x[47];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[6];
  assign t[37] = t[79] ^ x[1];
  assign t[38] = t[80] ^ x[2];
  assign t[39] = t[81] ^ x[3];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[82] ^ x[7];
  assign t[41] = t[83] ^ x[4];
  assign t[42] = t[84] ^ x[5];
  assign t[43] = t[85] ^ x[14];
  assign t[44] = t[86] ^ x[9];
  assign t[45] = t[87] ^ x[10];
  assign t[46] = t[88] ^ x[11];
  assign t[47] = t[89] ^ x[15];
  assign t[48] = t[90] ^ x[12];
  assign t[49] = t[91] ^ x[13];
  assign t[4] = ~(t[10] | t[5]);
  assign t[50] = t[92] ^ x[22];
  assign t[51] = t[93] ^ x[17];
  assign t[52] = t[94] ^ x[18];
  assign t[53] = t[95] ^ x[19];
  assign t[54] = t[96] ^ x[23];
  assign t[55] = t[97] ^ x[20];
  assign t[56] = t[98] ^ x[21];
  assign t[57] = t[99] ^ x[30];
  assign t[58] = t[100] ^ x[25];
  assign t[59] = t[101] ^ x[26];
  assign t[5] = ~(t[11]);
  assign t[60] = t[102] ^ x[27];
  assign t[61] = t[103] ^ x[31];
  assign t[62] = t[104] ^ x[28];
  assign t[63] = t[105] ^ x[29];
  assign t[64] = t[106] ^ x[38];
  assign t[65] = t[107] ^ x[33];
  assign t[66] = t[108] ^ x[34];
  assign t[67] = t[109] ^ x[35];
  assign t[68] = t[110] ^ x[39];
  assign t[69] = t[111] ^ x[36];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[37];
  assign t[71] = t[113] ^ x[46];
  assign t[72] = t[114] ^ x[41];
  assign t[73] = t[115] ^ x[42];
  assign t[74] = t[116] ^ x[43];
  assign t[75] = t[117] ^ x[47];
  assign t[76] = t[118] ^ x[44];
  assign t[77] = t[119] ^ x[45];
  assign t[78] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[79] = (x[0] & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[81] = (x[0] & ~1'b0) | (~x[0] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[86] = (x[8] & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0);
  assign t[87] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[88] = (x[8] & ~1'b0) | (~x[8] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[93] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[94] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[95] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[24] & ~1'b0 & ~1'b0) | (~x[24] & 1'b0 & ~1'b0) | (~x[24] & ~1'b0 & 1'b0) | (x[24] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind14(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = t[8] & t[9];
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind15(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = t[8] & t[9];
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind16(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = t[8] & t[9];
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind17(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(~x[0] & ~t[1]);
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] ? t[7] : t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] & t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = t[8] & t[9];
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind19(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind20(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind21(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind22(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind23(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind24(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind25(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind28(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[2] & t[6];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind29(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[2] & t[6];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind30(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[2] & t[6];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind31(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[2] & t[6];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[3] & t[7]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] | t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] & t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] | t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind32(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind33(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind34(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind35(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind36(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind37(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind38(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind39(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind40(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind41(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind42(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind43(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind44(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind45(x, y);
 input [8:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[10] = t[17] ^ x[8];
  assign t[11] = t[18] ^ x[5];
  assign t[12] = t[19] ^ x[6];
  assign t[13] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[14] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[15] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[16] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[17] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[1] = (t[2] & ~t[3]) | (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[7];
  assign t[3] = t[5] ^ x[8];
  assign t[4] = (t[6] & ~t[8] & ~t[9] & ~t[10] & ~t[11]) | (t[6] & ~t[7] & ~t[9] & ~t[10] & ~t[12]) | (t[6] & ~t[7] & ~t[8] & ~t[11] & ~t[12]) | (~t[6] & t[7] & t[8] & t[9] & ~t[12]) | (~t[6] & t[7] & t[10] & t[11] & ~t[12]) | (t[6] & ~t[8] & ~t[10] & t[12]) | (~t[6] & t[8] & t[10] & t[12]);
  assign t[5] = (t[6] & t[7] & ~t[8] & ~t[10] & t[11] & ~t[12]) | (t[6] & t[8] & ~t[9] & ~t[10] & ~t[11] & t[12]) | (~t[7] & ~t[8] & t[10] & ~t[11] & ~t[12]) | (~t[6] & ~t[8] & ~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[7] & ~t[9] & t[10] & ~t[12]) | (~t[6] & ~t[8] & t[9] & t[10] & t[11]) | (t[9] & t[10] & ~t[11] & ~t[12]);
  assign t[6] = t[13] ^ x[7];
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[3];
  assign t[9] = t[16] ^ x[4];
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind46(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind47(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind48(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind49(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] | t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind50(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] | t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0);
endmodule

module R2ind51(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] | t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind52(x, y);
 input [48:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~x[0] & t[1];
  assign t[100] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[101] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[102] = (x[25] & ~1'b0) | (~x[25] & 1'b0);
  assign t[103] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[104] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[107] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[108] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[109] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[10] = (t[20] & ~t[21]) | (~t[20] & t[21]);
  assign t[110] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[111] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[112] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[113] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[114] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[115] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[116] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[117] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[118] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = (t[22] & ~t[23]) | (~t[22] & t[23]);
  assign t[12] = t[24] ^ x[7];
  assign t[13] = t[25] ^ x[8];
  assign t[14] = t[26] ^ x[15];
  assign t[15] = t[27] ^ x[16];
  assign t[16] = t[28] ^ x[23];
  assign t[17] = t[29] ^ x[24];
  assign t[18] = t[30] ^ x[31];
  assign t[19] = t[31] ^ x[32];
  assign t[1] = t[6] | t[2];
  assign t[20] = t[32] ^ x[39];
  assign t[21] = t[33] ^ x[40];
  assign t[22] = t[34] ^ x[47];
  assign t[23] = t[35] ^ x[48];
  assign t[24] = (t[36] & ~t[38] & ~t[39] & ~t[40] & ~t[41]) | (t[36] & ~t[37] & ~t[39] & ~t[40] & ~t[42]) | (t[36] & ~t[37] & ~t[38] & ~t[41] & ~t[42]) | (~t[36] & t[37] & t[38] & t[39] & ~t[42]) | (~t[36] & t[37] & t[40] & t[41] & ~t[42]) | (t[36] & ~t[38] & ~t[40] & t[42]) | (~t[36] & t[38] & t[40] & t[42]);
  assign t[25] = (t[36] & t[37] & ~t[38] & ~t[40] & t[41] & ~t[42]) | (t[36] & t[38] & ~t[39] & ~t[40] & ~t[41] & t[42]) | (~t[37] & ~t[38] & t[40] & ~t[41] & ~t[42]) | (~t[36] & ~t[38] & ~t[39] & t[40] & ~t[41]) | (~t[36] & ~t[37] & ~t[39] & t[40] & ~t[42]) | (~t[36] & ~t[38] & t[39] & t[40] & t[41]) | (t[39] & t[40] & ~t[41] & ~t[42]);
  assign t[26] = (t[43] & ~t[45] & ~t[46] & ~t[47] & ~t[48]) | (t[43] & ~t[44] & ~t[46] & ~t[47] & ~t[49]) | (t[43] & ~t[44] & ~t[45] & ~t[48] & ~t[49]) | (~t[43] & t[44] & t[45] & t[46] & ~t[49]) | (~t[43] & t[44] & t[47] & t[48] & ~t[49]) | (t[43] & ~t[45] & ~t[47] & t[49]) | (~t[43] & t[45] & t[47] & t[49]);
  assign t[27] = (t[43] & t[44] & ~t[45] & ~t[47] & t[48] & ~t[49]) | (t[43] & t[45] & ~t[46] & ~t[47] & ~t[48] & t[49]) | (~t[44] & ~t[45] & t[47] & ~t[48] & ~t[49]) | (~t[43] & ~t[45] & ~t[46] & t[47] & ~t[48]) | (~t[43] & ~t[44] & ~t[46] & t[47] & ~t[49]) | (~t[43] & ~t[45] & t[46] & t[47] & t[48]) | (t[46] & t[47] & ~t[48] & ~t[49]);
  assign t[28] = (t[50] & ~t[52] & ~t[53] & ~t[54] & ~t[55]) | (t[50] & ~t[51] & ~t[53] & ~t[54] & ~t[56]) | (t[50] & ~t[51] & ~t[52] & ~t[55] & ~t[56]) | (~t[50] & t[51] & t[52] & t[53] & ~t[56]) | (~t[50] & t[51] & t[54] & t[55] & ~t[56]) | (t[50] & ~t[52] & ~t[54] & t[56]) | (~t[50] & t[52] & t[54] & t[56]);
  assign t[29] = (t[50] & t[51] & ~t[52] & ~t[54] & t[55] & ~t[56]) | (t[50] & t[52] & ~t[53] & ~t[54] & ~t[55] & t[56]) | (~t[51] & ~t[52] & t[54] & ~t[55] & ~t[56]) | (~t[50] & ~t[52] & ~t[53] & t[54] & ~t[55]) | (~t[50] & ~t[51] & ~t[53] & t[54] & ~t[56]) | (~t[50] & ~t[52] & t[53] & t[54] & t[55]) | (t[53] & t[54] & ~t[55] & ~t[56]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (t[57] & ~t[59] & ~t[60] & ~t[61] & ~t[62]) | (t[57] & ~t[58] & ~t[60] & ~t[61] & ~t[63]) | (t[57] & ~t[58] & ~t[59] & ~t[62] & ~t[63]) | (~t[57] & t[58] & t[59] & t[60] & ~t[63]) | (~t[57] & t[58] & t[61] & t[62] & ~t[63]) | (t[57] & ~t[59] & ~t[61] & t[63]) | (~t[57] & t[59] & t[61] & t[63]);
  assign t[31] = (t[57] & t[58] & ~t[59] & ~t[61] & t[62] & ~t[63]) | (t[57] & t[59] & ~t[60] & ~t[61] & ~t[62] & t[63]) | (~t[58] & ~t[59] & t[61] & ~t[62] & ~t[63]) | (~t[57] & ~t[59] & ~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[58] & ~t[60] & t[61] & ~t[63]) | (~t[57] & ~t[59] & t[60] & t[61] & t[62]) | (t[60] & t[61] & ~t[62] & ~t[63]);
  assign t[32] = (t[64] & ~t[66] & ~t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[67] & ~t[68] & ~t[70]) | (t[64] & ~t[65] & ~t[66] & ~t[69] & ~t[70]) | (~t[64] & t[65] & t[66] & t[67] & ~t[70]) | (~t[64] & t[65] & t[68] & t[69] & ~t[70]) | (t[64] & ~t[66] & ~t[68] & t[70]) | (~t[64] & t[66] & t[68] & t[70]);
  assign t[33] = (t[64] & t[65] & ~t[66] & ~t[68] & t[69] & ~t[70]) | (t[64] & t[66] & ~t[67] & ~t[68] & ~t[69] & t[70]) | (~t[65] & ~t[66] & t[68] & ~t[69] & ~t[70]) | (~t[64] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[65] & ~t[67] & t[68] & ~t[70]) | (~t[64] & ~t[66] & t[67] & t[68] & t[69]) | (t[67] & t[68] & ~t[69] & ~t[70]);
  assign t[34] = (t[71] & ~t[73] & ~t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[74] & ~t[75] & ~t[77]) | (t[71] & ~t[72] & ~t[73] & ~t[76] & ~t[77]) | (~t[71] & t[72] & t[73] & t[74] & ~t[77]) | (~t[71] & t[72] & t[75] & t[76] & ~t[77]) | (t[71] & ~t[73] & ~t[75] & t[77]) | (~t[71] & t[73] & t[75] & t[77]);
  assign t[35] = (t[71] & t[72] & ~t[73] & ~t[75] & t[76] & ~t[77]) | (t[71] & t[73] & ~t[74] & ~t[75] & ~t[76] & t[77]) | (~t[72] & ~t[73] & t[75] & ~t[76] & ~t[77]) | (~t[71] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[72] & ~t[74] & t[75] & ~t[77]) | (~t[71] & ~t[73] & t[74] & t[75] & t[76]) | (t[74] & t[75] & ~t[76] & ~t[77]);
  assign t[36] = t[78] ^ x[7];
  assign t[37] = t[79] ^ x[2];
  assign t[38] = t[80] ^ x[3];
  assign t[39] = t[81] ^ x[4];
  assign t[3] = ~(t[8] & t[4]);
  assign t[40] = t[82] ^ x[8];
  assign t[41] = t[83] ^ x[5];
  assign t[42] = t[84] ^ x[6];
  assign t[43] = t[85] ^ x[15];
  assign t[44] = t[86] ^ x[10];
  assign t[45] = t[87] ^ x[11];
  assign t[46] = t[88] ^ x[12];
  assign t[47] = t[89] ^ x[16];
  assign t[48] = t[90] ^ x[13];
  assign t[49] = t[91] ^ x[14];
  assign t[4] = ~(t[9] | t[5]);
  assign t[50] = t[92] ^ x[23];
  assign t[51] = t[93] ^ x[18];
  assign t[52] = t[94] ^ x[19];
  assign t[53] = t[95] ^ x[20];
  assign t[54] = t[96] ^ x[24];
  assign t[55] = t[97] ^ x[21];
  assign t[56] = t[98] ^ x[22];
  assign t[57] = t[99] ^ x[31];
  assign t[58] = t[100] ^ x[26];
  assign t[59] = t[101] ^ x[27];
  assign t[5] = ~(t[10] & t[11]);
  assign t[60] = t[102] ^ x[28];
  assign t[61] = t[103] ^ x[32];
  assign t[62] = t[104] ^ x[29];
  assign t[63] = t[105] ^ x[30];
  assign t[64] = t[106] ^ x[39];
  assign t[65] = t[107] ^ x[34];
  assign t[66] = t[108] ^ x[35];
  assign t[67] = t[109] ^ x[36];
  assign t[68] = t[110] ^ x[40];
  assign t[69] = t[111] ^ x[37];
  assign t[6] = (t[12] & ~t[13]) | (~t[12] & t[13]);
  assign t[70] = t[112] ^ x[38];
  assign t[71] = t[113] ^ x[47];
  assign t[72] = t[114] ^ x[42];
  assign t[73] = t[115] ^ x[43];
  assign t[74] = t[116] ^ x[44];
  assign t[75] = t[117] ^ x[48];
  assign t[76] = t[118] ^ x[45];
  assign t[77] = t[119] ^ x[46];
  assign t[78] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[79] = (x[1] & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0);
  assign t[7] = (t[14] & ~t[15]) | (~t[14] & t[15]);
  assign t[80] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[81] = (x[1] & ~1'b0) | (~x[1] & 1'b0);
  assign t[82] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[83] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[84] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[85] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[86] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[87] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[88] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[89] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[8] = (t[16] & ~t[17]) | (~t[16] & t[17]);
  assign t[90] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[91] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[92] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[93] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[94] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[95] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[96] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[97] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[98] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[99] = (x[25] & ~1'b0 & ~1'b0) | (~x[25] & 1'b0 & ~1'b0) | (~x[25] & ~1'b0 & 1'b0) | (x[25] & 1'b0 & 1'b0);
  assign t[9] = (t[18] & ~t[19]) | (~t[18] & t[19]);
  assign y = (t[0] & ~1'b0) | (~t[0] & 1'b0);
endmodule

module R2ind53(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind54(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind55(y);
 output y;

  assign y = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
endmodule

module R2ind56(x, y);
 input [36:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[101] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[102] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[103] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[104] = (t[108] & t[109] & ~t[110] & t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[110] & ~t[111] & t[112] & ~t[113] & t[114]) | (~t[109] & t[110] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[109] & t[110] & ~t[113] & ~t[114]) | (~t[108] & t[110] & t[111] & ~t[112] & t[113]) | (t[110] & ~t[111] & t[113] & ~t[114]);
  assign t[105] = (t[109] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & t[109] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[109] & ~t[110] & ~t[113] & ~t[114]) | (t[108] & ~t[109] & t[110] & t[111] & ~t[114]) | (t[108] & ~t[109] & t[112] & t[113] & ~t[114]) | (t[109] & ~t[111] & ~t[113] & t[114]) | (~t[109] & t[111] & t[113] & t[114]);
  assign t[106] = (t[108] & t[109] & t[110] & ~t[111] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[111] & ~t[112] & t[113] & t[114]) | (~t[109] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[110] & t[111] & ~t[113] & ~t[114]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[114]) | (~t[109] & t[110] & t[111] & t[112] & ~t[113]) | (~t[110] & t[111] & t[112] & ~t[114]);
  assign t[107] = (t[108] & t[109] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[108] & ~t[109] & ~t[110] & t[113] & ~t[114]) | (~t[109] & t[110] & ~t[111] & t[112] & t[113]) | (t[110] & ~t[112] & t[113] & ~t[114]);
  assign t[108] = t[129] ^ x[7];
  assign t[109] = t[130] ^ x[34];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[32];
  assign t[111] = t[132] ^ x[35];
  assign t[112] = t[133] ^ x[8];
  assign t[113] = t[134] ^ x[36];
  assign t[114] = t[135] ^ x[6];
  assign t[115] = t[136] ^ x[14];
  assign t[116] = t[137] ^ x[16];
  assign t[117] = t[138] ^ x[15];
  assign t[118] = t[139] ^ x[17];
  assign t[119] = t[140] ^ x[18];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[19];
  assign t[121] = t[142] ^ x[13];
  assign t[122] = t[143] ^ x[25];
  assign t[123] = t[144] ^ x[27];
  assign t[124] = t[145] ^ x[26];
  assign t[125] = t[146] ^ x[28];
  assign t[126] = t[147] ^ x[29];
  assign t[127] = t[148] ^ x[30];
  assign t[128] = t[149] ^ x[24];
  assign t[129] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[131] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[132] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[133] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[134] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[135] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[136] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[137] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[138] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[139] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[141] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[142] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[143] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[144] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[145] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[146] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[147] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[148] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[149] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[63]);
  assign t[15] = ~(t[62] ^ t[14]);
  assign t[16] = t[64] ^ t[63];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[62] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[62] ^ t[27];
  assign t[23] = t[65] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[63] ^ t[66];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[67]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[65] ^ t[29]);
  assign t[31] = t[68] ^ t[67];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[65] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[65] ^ t[36];
  assign t[36] = t[67] ^ t[69];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[70]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[62] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[61]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[65] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[71]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[62] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[63] = (t[74] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[74] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[64] = (t[74] & ~t[78]) | (~t[74] & t[78]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[74] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[74] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[67] = (t[80] & ~t[83] & ~t[85]) | (~t[82] & t[83] & ~t[84]) | (~t[80] & ~t[83] & t[85]) | (t[82] & t[83] & t[84]);
  assign t[68] = (t[80] & ~t[84]) | (~t[80] & t[84]);
  assign t[69] = (t[80] & ~t[83] & ~t[84]) | (~t[82] & t[83] & ~t[85]) | (~t[80] & ~t[83] & t[84]) | (t[82] & t[83] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[72] & ~t[86]) | (~t[72] & t[86]);
  assign t[71] = (t[72] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[73]) | (~t[72] & ~t[88] & t[89]) | (t[87] & t[88] & t[73]);
  assign t[72] = t[90] ^ x[7];
  assign t[73] = t[91] ^ x[8];
  assign t[74] = t[92] ^ x[14];
  assign t[75] = t[93] ^ x[15];
  assign t[76] = t[94] ^ x[16];
  assign t[77] = t[95] ^ x[17];
  assign t[78] = t[96] ^ x[18];
  assign t[79] = t[97] ^ x[19];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[25];
  assign t[81] = t[99] ^ x[26];
  assign t[82] = t[100] ^ x[27];
  assign t[83] = t[101] ^ x[28];
  assign t[84] = t[102] ^ x[29];
  assign t[85] = t[103] ^ x[30];
  assign t[86] = t[104] ^ x[32];
  assign t[87] = t[105] ^ x[34];
  assign t[88] = t[106] ^ x[35];
  assign t[89] = t[107] ^ x[36];
  assign t[8] = t[62] & t[13];
  assign t[90] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[91] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[92] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[93] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[94] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[95] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[96] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[97] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[98] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[99] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind57(x, y);
 input [36:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[101] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[102] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[103] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[104] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[105] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[106] = t[127] ^ x[7];
  assign t[107] = t[128] ^ x[34];
  assign t[108] = t[129] ^ x[32];
  assign t[109] = t[130] ^ x[35];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[8];
  assign t[111] = t[132] ^ x[36];
  assign t[112] = t[133] ^ x[6];
  assign t[113] = t[134] ^ x[14];
  assign t[114] = t[135] ^ x[16];
  assign t[115] = t[136] ^ x[15];
  assign t[116] = t[137] ^ x[17];
  assign t[117] = t[138] ^ x[18];
  assign t[118] = t[139] ^ x[19];
  assign t[119] = t[140] ^ x[13];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[25];
  assign t[121] = t[142] ^ x[27];
  assign t[122] = t[143] ^ x[26];
  assign t[123] = t[144] ^ x[28];
  assign t[124] = t[145] ^ x[29];
  assign t[125] = t[146] ^ x[30];
  assign t[126] = t[147] ^ x[24];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[135] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[136] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[137] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[138] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[139] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[141] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[142] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[143] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[144] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[145] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[146] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[147] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[61]);
  assign t[15] = ~(t[60] ^ t[14]);
  assign t[16] = t[62] ^ t[61];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[60] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[60] ^ t[27];
  assign t[23] = t[63] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[61] ^ t[64];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[65]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[63] ^ t[29]);
  assign t[31] = t[66] ^ t[65];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[63] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[63] ^ t[36];
  assign t[36] = t[65] ^ t[67];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[68]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[60] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[59]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[63] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[42]);
  assign t[56] = ~(t[57] ^ t[69]);
  assign t[57] = ~t[58];
  assign t[58] = ~(t[48]);
  assign t[59] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[61] = (t[72] & ~t[75] & ~t[77]) | (~t[74] & t[75] & ~t[76]) | (~t[72] & ~t[75] & t[77]) | (t[74] & t[75] & t[76]);
  assign t[62] = (t[72] & ~t[76]) | (~t[72] & t[76]);
  assign t[63] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[64] = (t[72] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[77]) | (~t[72] & ~t[75] & t[76]) | (t[74] & t[75] & t[77]);
  assign t[65] = (t[78] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[78] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[66] = (t[78] & ~t[82]) | (~t[78] & t[82]);
  assign t[67] = (t[78] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[78] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[68] = (t[70] & ~t[84]) | (~t[70] & t[84]);
  assign t[69] = (t[70] & ~t[86] & ~t[71]) | (~t[85] & t[86] & ~t[87]) | (~t[70] & ~t[86] & t[71]) | (t[85] & t[86] & t[87]);
  assign t[6] = t[10] & t[11];
  assign t[70] = t[88] ^ x[7];
  assign t[71] = t[89] ^ x[8];
  assign t[72] = t[90] ^ x[14];
  assign t[73] = t[91] ^ x[15];
  assign t[74] = t[92] ^ x[16];
  assign t[75] = t[93] ^ x[17];
  assign t[76] = t[94] ^ x[18];
  assign t[77] = t[95] ^ x[19];
  assign t[78] = t[96] ^ x[25];
  assign t[79] = t[97] ^ x[26];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[27];
  assign t[81] = t[99] ^ x[28];
  assign t[82] = t[100] ^ x[29];
  assign t[83] = t[101] ^ x[30];
  assign t[84] = t[102] ^ x[32];
  assign t[85] = t[103] ^ x[34];
  assign t[86] = t[104] ^ x[35];
  assign t[87] = t[105] ^ x[36];
  assign t[88] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[89] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[8] = t[60] & t[13];
  assign t[90] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[93] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[96] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[97] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[98] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[99] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind58(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[19];
  assign t[102] = t[123] ^ x[20];
  assign t[103] = t[124] ^ x[14];
  assign t[104] = t[125] ^ x[26];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[27];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[30];
  assign t[109] = t[130] ^ x[31];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[25];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[119] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[121] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[122] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[123] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[124] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[125] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[126] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[127] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[128] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[129] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[131] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[48]);
  assign t[15] = ~(t[47] ^ t[14]);
  assign t[16] = t[49] ^ t[48];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[47] ^ t[27];
  assign t[23] = t[50] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[48] ^ t[51];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[52]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[50] ^ t[29]);
  assign t[31] = t[53] ^ t[52];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[50] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[50] ^ t[36];
  assign t[36] = t[52] ^ t[54];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[27] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[36] ^ t[24];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[58] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[49] = (t[58] & ~t[62]) | (~t[58] & t[62]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[58] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[52] = (t[64] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[64] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[64] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[57]) | (~t[56] & ~t[71] & t[72]) | (t[70] & t[71] & t[57]);
  assign t[56] = t[73] ^ x[8];
  assign t[57] = t[74] ^ x[9];
  assign t[58] = t[75] ^ x[15];
  assign t[59] = t[76] ^ x[16];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[17];
  assign t[61] = t[78] ^ x[18];
  assign t[62] = t[79] ^ x[19];
  assign t[63] = t[80] ^ x[20];
  assign t[64] = t[81] ^ x[26];
  assign t[65] = t[82] ^ x[27];
  assign t[66] = t[83] ^ x[28];
  assign t[67] = t[84] ^ x[29];
  assign t[68] = t[85] ^ x[30];
  assign t[69] = t[86] ^ x[31];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[33];
  assign t[71] = t[88] ^ x[34];
  assign t[72] = t[89] ^ x[35];
  assign t[73] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[86] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[87] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[88] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[47] & t[13];
  assign t[90] = t[111] ^ x[8];
  assign t[91] = t[112] ^ x[33];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[9];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[15];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[16];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind59(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[20];
  assign t[105] = t[126] ^ x[14];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[31];
  assign t[112] = t[133] ^ x[25];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[121] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[122] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[123] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[126] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[127] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[128] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[129] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[132] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[133] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[50]);
  assign t[15] = ~(t[49] ^ t[14]);
  assign t[16] = t[51] ^ t[50];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[49] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[49] ^ t[27];
  assign t[23] = t[52] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[50] ^ t[53];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[54]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[52] ^ t[29]);
  assign t[31] = t[55] ^ t[54];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[52] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[52] ^ t[36];
  assign t[36] = t[54] ^ t[56];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[57]);
  assign t[42] = t[44] ^ t[9];
  assign t[43] = ~t[45];
  assign t[44] = t[16] ^ t[21];
  assign t[45] = ~(t[46]);
  assign t[46] = t[47] ^ t[24];
  assign t[47] = t[31] ^ t[34];
  assign t[48] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[49] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[60] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[60] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[51] = (t[60] & ~t[64]) | (~t[60] & t[64]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[60] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[60] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[54] = (t[66] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[66] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[55] = (t[66] & ~t[70]) | (~t[66] & t[70]);
  assign t[56] = (t[66] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[66] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[57] = (t[58] & ~t[73] & ~t[59]) | (~t[72] & t[73] & ~t[74]) | (~t[58] & ~t[73] & t[59]) | (t[72] & t[73] & t[74]);
  assign t[58] = t[75] ^ x[8];
  assign t[59] = t[76] ^ x[9];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[15];
  assign t[61] = t[78] ^ x[16];
  assign t[62] = t[79] ^ x[17];
  assign t[63] = t[80] ^ x[18];
  assign t[64] = t[81] ^ x[19];
  assign t[65] = t[82] ^ x[20];
  assign t[66] = t[83] ^ x[26];
  assign t[67] = t[84] ^ x[27];
  assign t[68] = t[85] ^ x[28];
  assign t[69] = t[86] ^ x[29];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[30];
  assign t[71] = t[88] ^ x[31];
  assign t[72] = t[89] ^ x[33];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[35];
  assign t[75] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[76] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[77] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[8] = t[49] & t[13];
  assign t[90] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[7];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind60(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[15];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[16];
  assign t[104] = t[125] ^ x[19];
  assign t[105] = t[126] ^ x[13];
  assign t[106] = t[127] ^ x[25];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[26];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[27];
  assign t[111] = t[132] ^ x[30];
  assign t[112] = t[133] ^ x[24];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[47] ^ t[15];
  assign t[120] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[121] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[122] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[123] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[124] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[125] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[126] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[127] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[128] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[129] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[131] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[132] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[133] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[48] ^ t[49];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[49]);
  assign t[16] = ~(t[47] ^ t[15]);
  assign t[17] = t[47] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[50] ^ t[30];
  assign t[26] = t[49] ^ t[51];
  assign t[27] = t[47] ^ t[13];
  assign t[28] = t[52] ^ t[53];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[50] ^ t[30]);
  assign t[32] = t[50] & t[34];
  assign t[33] = t[50] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[53] ^ t[54];
  assign t[36] = t[50] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[26] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[35] ^ t[23];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[60]) | (~t[58] & t[60]);
  assign t[49] = (t[58] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[60]) | (~t[58] & ~t[62] & t[63]) | (t[61] & t[62] & t[60]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[62] & ~t[60]) | (~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[62] & t[60]) | (t[61] & t[62] & t[63]);
  assign t[52] = (t[64] & ~t[66]) | (~t[64] & t[66]);
  assign t[53] = (t[64] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[66]) | (~t[64] & ~t[68] & t[69]) | (t[67] & t[68] & t[66]);
  assign t[54] = (t[64] & ~t[68] & ~t[66]) | (~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[68] & t[66]) | (t[67] & t[68] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[56] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = t[74] ^ x[7];
  assign t[57] = t[75] ^ x[8];
  assign t[58] = t[76] ^ x[14];
  assign t[59] = t[77] ^ x[15];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[16];
  assign t[61] = t[79] ^ x[17];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[19];
  assign t[64] = t[82] ^ x[25];
  assign t[65] = t[83] ^ x[26];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[29];
  assign t[69] = t[87] ^ x[30];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[32];
  assign t[71] = t[89] ^ x[33];
  assign t[72] = t[90] ^ x[34];
  assign t[73] = t[91] ^ x[35];
  assign t[74] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[83] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[89] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[7];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[8];
  assign t[95] = t[116] ^ x[33];
  assign t[96] = t[117] ^ x[34];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[6];
  assign t[99] = t[120] ^ x[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind61(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[19];
  assign t[103] = t[124] ^ x[13];
  assign t[104] = t[125] ^ x[25];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[30];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[24];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[119] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[11] = t[45] ^ t[15];
  assign t[120] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[121] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[122] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[123] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[126] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[127] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[128] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[129] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[46] ^ t[47];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[47]);
  assign t[16] = ~(t[45] ^ t[15]);
  assign t[17] = t[45] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[45] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[48] ^ t[30];
  assign t[26] = t[47] ^ t[49];
  assign t[27] = t[45] ^ t[13];
  assign t[28] = t[50] ^ t[51];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[51]);
  assign t[31] = ~(t[48] ^ t[30]);
  assign t[32] = t[48] & t[34];
  assign t[33] = t[48] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[51] ^ t[52];
  assign t[36] = t[48] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[5]);
  assign t[41] = ~(t[42] ^ t[53]);
  assign t[42] = ~t[43];
  assign t[43] = ~(t[18]);
  assign t[44] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[56] & ~t[58]) | (~t[56] & t[58]);
  assign t[47] = (t[56] & ~t[60] & ~t[61]) | (~t[59] & t[60] & ~t[58]) | (~t[56] & ~t[60] & t[61]) | (t[59] & t[60] & t[58]);
  assign t[48] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[49] = (t[56] & ~t[60] & ~t[58]) | (~t[59] & t[60] & ~t[61]) | (~t[56] & ~t[60] & t[58]) | (t[59] & t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[44]);
  assign t[50] = (t[62] & ~t[64]) | (~t[62] & t[64]);
  assign t[51] = (t[62] & ~t[66] & ~t[67]) | (~t[65] & t[66] & ~t[64]) | (~t[62] & ~t[66] & t[67]) | (t[65] & t[66] & t[64]);
  assign t[52] = (t[62] & ~t[66] & ~t[64]) | (~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[66] & t[64]) | (t[65] & t[66] & t[67]);
  assign t[53] = (t[54] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[54] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[54] = t[72] ^ x[7];
  assign t[55] = t[73] ^ x[8];
  assign t[56] = t[74] ^ x[14];
  assign t[57] = t[75] ^ x[15];
  assign t[58] = t[76] ^ x[16];
  assign t[59] = t[77] ^ x[17];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[25];
  assign t[63] = t[81] ^ x[26];
  assign t[64] = t[82] ^ x[27];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[29];
  assign t[67] = t[85] ^ x[30];
  assign t[68] = t[86] ^ x[32];
  assign t[69] = t[87] ^ x[33];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[34];
  assign t[71] = t[89] ^ x[35];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[81] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[86] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[87] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[88] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[111] ^ x[7];
  assign t[91] = t[112] ^ x[32];
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[6];
  assign t[97] = t[118] ^ x[14];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind62(x, y);
 input [35:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[101] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[102] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[103] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[104] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[105] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[35]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[114] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[115] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[116] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[118] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[119] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[11] = ~(t[37] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[38] ^ t[39];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = x[0] ? x[35] : t[18];
  assign t[18] = ~(t[19] ^ t[20]);
  assign t[19] = ~t[21];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[23] ^ t[41]);
  assign t[22] = t[24] ^ t[8];
  assign t[23] = ~t[25];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = ~(t[28]);
  assign t[26] = t[42] ^ t[35];
  assign t[27] = t[10] & t[29];
  assign t[28] = t[30] ^ t[14];
  assign t[29] = t[37] ^ t[7];
  assign t[2] = ~t[4];
  assign t[30] = t[31] ^ t[32];
  assign t[31] = t[43] ^ t[38];
  assign t[32] = t[15] & t[33];
  assign t[33] = t[40] ^ t[13];
  assign t[34] = (t[44] & ~t[46] & ~t[48]) | (~t[45] & t[46] & ~t[47]) | (~t[44] & ~t[46] & t[48]) | (t[45] & t[46] & t[47]);
  assign t[35] = (t[49] & ~t[51] & ~t[53]) | (~t[50] & t[51] & ~t[52]) | (~t[49] & ~t[51] & t[53]) | (t[50] & t[51] & t[52]);
  assign t[36] = (t[49] & ~t[51] & ~t[52]) | (~t[50] & t[51] & ~t[53]) | (~t[49] & ~t[51] & t[52]) | (t[50] & t[51] & t[53]);
  assign t[37] = (t[49] & ~t[54]) | (~t[49] & t[54]);
  assign t[38] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[39] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[60]) | (~t[55] & t[60]);
  assign t[41] = (t[44] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[44] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[42] = (t[49] & ~t[52]) | (~t[49] & t[52]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = t[61] ^ x[8];
  assign t[45] = t[62] ^ x[9];
  assign t[46] = t[63] ^ x[10];
  assign t[47] = t[64] ^ x[11];
  assign t[48] = t[65] ^ x[12];
  assign t[49] = t[66] ^ x[18];
  assign t[4] = ~(t[6] ^ t[34]);
  assign t[50] = t[67] ^ x[19];
  assign t[51] = t[68] ^ x[20];
  assign t[52] = t[69] ^ x[21];
  assign t[53] = t[70] ^ x[22];
  assign t[54] = t[71] ^ x[23];
  assign t[55] = t[72] ^ x[29];
  assign t[56] = t[73] ^ x[30];
  assign t[57] = t[74] ^ x[31];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[34];
  assign t[61] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[62] = (t[79] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (~t[78] & t[79] & ~t[81] & ~t[82] & ~t[84]) | (~t[78] & t[79] & ~t[80] & ~t[83] & ~t[84]) | (t[78] & ~t[79] & t[80] & t[81] & ~t[84]) | (t[78] & ~t[79] & t[82] & t[83] & ~t[84]) | (t[79] & ~t[81] & ~t[83] & t[84]) | (~t[79] & t[81] & t[83] & t[84]);
  assign t[63] = (t[78] & t[79] & t[80] & ~t[81] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & ~t[81] & ~t[82] & t[83] & t[84]) | (~t[79] & ~t[80] & t[81] & ~t[82] & ~t[83]) | (~t[78] & ~t[80] & t[81] & ~t[83] & ~t[84]) | (~t[78] & ~t[79] & t[81] & ~t[82] & ~t[84]) | (~t[79] & t[80] & t[81] & t[82] & ~t[83]) | (~t[80] & t[81] & t[82] & ~t[84]);
  assign t[64] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[65] = (t[78] & t[79] & ~t[81] & t[82] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & ~t[81] & ~t[82] & t[83]) | (~t[78] & ~t[81] & ~t[82] & t[83] & ~t[84]) | (~t[78] & ~t[79] & ~t[80] & t[83] & ~t[84]) | (~t[79] & t[80] & ~t[81] & t[82] & t[83]) | (t[80] & ~t[82] & t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = ~t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[72] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[73] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[74] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[8];
  assign t[79] = t[100] ^ x[9];
  assign t[7] = t[35] ^ t[36];
  assign t[80] = t[101] ^ x[6];
  assign t[81] = t[102] ^ x[10];
  assign t[82] = t[103] ^ x[11];
  assign t[83] = t[104] ^ x[12];
  assign t[84] = t[105] ^ x[7];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[23];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[29];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[32];
  assign t[97] = t[118] ^ x[33];
  assign t[98] = t[119] ^ x[28];
  assign t[99] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~t[17]) | (~t[0] & t[17]);
endmodule

module R2ind63(x, y);
 input [36:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & t[124] & ~t[125] & t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[125] & ~t[126] & t[127] & ~t[128] & t[129]) | (~t[124] & t[125] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[124] & t[125] & ~t[128] & ~t[129]) | (~t[123] & t[125] & t[126] & ~t[127] & t[128]) | (t[125] & ~t[126] & t[128] & ~t[129]);
  assign t[101] = (t[124] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & t[124] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[124] & ~t[125] & ~t[128] & ~t[129]) | (t[123] & ~t[124] & t[125] & t[126] & ~t[129]) | (t[123] & ~t[124] & t[127] & t[128] & ~t[129]) | (t[124] & ~t[126] & ~t[128] & t[129]) | (~t[124] & t[126] & t[128] & t[129]);
  assign t[102] = (t[123] & t[124] & t[125] & ~t[126] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[126] & ~t[127] & t[128] & t[129]) | (~t[124] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[125] & t[126] & ~t[128] & ~t[129]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[129]) | (~t[124] & t[125] & t[126] & t[127] & ~t[128]) | (~t[125] & t[126] & t[127] & ~t[129]);
  assign t[103] = (t[123] & t[124] & ~t[125] & ~t[127] & t[128] & ~t[129]) | (t[123] & t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[129]) | (~t[123] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[123] & ~t[124] & ~t[126] & t[127] & ~t[129]) | (~t[123] & ~t[125] & t[126] & t[127] & t[128]) | (t[126] & t[127] & ~t[128] & ~t[129]);
  assign t[104] = (t[123] & t[124] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[123] & ~t[124] & ~t[125] & t[128] & ~t[129]) | (~t[124] & t[125] & ~t[126] & t[127] & t[128]) | (t[125] & ~t[127] & t[128] & ~t[129]);
  assign t[105] = (t[109] & t[110] & ~t[111] & t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[111] & ~t[112] & t[113] & ~t[114] & t[115]) | (~t[110] & t[111] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[110] & t[111] & ~t[114] & ~t[115]) | (~t[109] & t[111] & t[112] & ~t[113] & t[114]) | (t[111] & ~t[112] & t[114] & ~t[115]);
  assign t[106] = (t[110] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & t[110] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[110] & ~t[111] & ~t[114] & ~t[115]) | (t[109] & ~t[110] & t[111] & t[112] & ~t[115]) | (t[109] & ~t[110] & t[113] & t[114] & ~t[115]) | (t[110] & ~t[112] & ~t[114] & t[115]) | (~t[110] & t[112] & t[114] & t[115]);
  assign t[107] = (t[109] & t[110] & t[111] & ~t[112] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[112] & ~t[113] & t[114] & t[115]) | (~t[110] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[111] & t[112] & ~t[114] & ~t[115]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[115]) | (~t[110] & t[111] & t[112] & t[113] & ~t[114]) | (~t[111] & t[112] & t[113] & ~t[115]);
  assign t[108] = (t[109] & t[110] & ~t[112] & t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[109] & ~t[110] & ~t[111] & t[114] & ~t[115]) | (~t[110] & t[111] & ~t[112] & t[113] & t[114]) | (t[111] & ~t[113] & t[114] & ~t[115]);
  assign t[109] = t[130] ^ x[7];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[34];
  assign t[111] = t[132] ^ x[32];
  assign t[112] = t[133] ^ x[35];
  assign t[113] = t[134] ^ x[8];
  assign t[114] = t[135] ^ x[36];
  assign t[115] = t[136] ^ x[6];
  assign t[116] = t[137] ^ x[14];
  assign t[117] = t[138] ^ x[16];
  assign t[118] = t[139] ^ x[15];
  assign t[119] = t[140] ^ x[17];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[18];
  assign t[121] = t[142] ^ x[19];
  assign t[122] = t[143] ^ x[13];
  assign t[123] = t[144] ^ x[25];
  assign t[124] = t[145] ^ x[27];
  assign t[125] = t[146] ^ x[26];
  assign t[126] = t[147] ^ x[28];
  assign t[127] = t[148] ^ x[29];
  assign t[128] = t[149] ^ x[30];
  assign t[129] = t[150] ^ x[24];
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[131] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[132] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[133] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[134] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[135] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[136] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[137] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[138] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[139] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[141] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[142] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[143] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[144] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[145] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[146] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[147] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[148] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[149] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[14] = ~(t[64]);
  assign t[150] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[15] = ~(t[63] ^ t[14]);
  assign t[16] = t[65] ^ t[64];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[63] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[63] ^ t[27];
  assign t[23] = t[66] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[64] ^ t[67];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[68]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[66] ^ t[29]);
  assign t[31] = t[69] ^ t[68];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[66] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[66] ^ t[36];
  assign t[36] = t[68] ^ t[70];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[71]);
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~t[46];
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~(t[49] ^ t[50]);
  assign t[47] = t[16] ^ t[21];
  assign t[48] = t[63] ^ t[14];
  assign t[49] = t[51] ^ t[24];
  assign t[4] = ~(t[7] ^ t[62]);
  assign t[50] = t[18] ^ t[52];
  assign t[51] = t[31] ^ t[34];
  assign t[52] = t[66] ^ t[29];
  assign t[53] = x[0] ? x[33] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~t[57];
  assign t[56] = ~(t[58]);
  assign t[57] = ~(t[59] ^ t[72]);
  assign t[58] = t[27] ^ t[9];
  assign t[59] = ~t[60];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[61]);
  assign t[61] = t[36] ^ t[24];
  assign t[62] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[63] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[64] = (t[75] & ~t[78] & ~t[80]) | (~t[77] & t[78] & ~t[79]) | (~t[75] & ~t[78] & t[80]) | (t[77] & t[78] & t[79]);
  assign t[65] = (t[75] & ~t[79]) | (~t[75] & t[79]);
  assign t[66] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[67] = (t[75] & ~t[78] & ~t[79]) | (~t[77] & t[78] & ~t[80]) | (~t[75] & ~t[78] & t[79]) | (t[77] & t[78] & t[80]);
  assign t[68] = (t[81] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[81] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[69] = (t[81] & ~t[85]) | (~t[81] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[81] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[81] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[71] = (t[73] & ~t[87]) | (~t[73] & t[87]);
  assign t[72] = (t[73] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[74]) | (~t[73] & ~t[89] & t[90]) | (t[88] & t[89] & t[74]);
  assign t[73] = t[91] ^ x[7];
  assign t[74] = t[92] ^ x[8];
  assign t[75] = t[93] ^ x[14];
  assign t[76] = t[94] ^ x[15];
  assign t[77] = t[95] ^ x[16];
  assign t[78] = t[96] ^ x[17];
  assign t[79] = t[97] ^ x[18];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[19];
  assign t[81] = t[99] ^ x[25];
  assign t[82] = t[100] ^ x[26];
  assign t[83] = t[101] ^ x[27];
  assign t[84] = t[102] ^ x[28];
  assign t[85] = t[103] ^ x[29];
  assign t[86] = t[104] ^ x[30];
  assign t[87] = t[105] ^ x[32];
  assign t[88] = t[106] ^ x[34];
  assign t[89] = t[107] ^ x[35];
  assign t[8] = t[63] & t[13];
  assign t[90] = t[108] ^ x[36];
  assign t[91] = (t[109] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[110] & ~t[111] & ~t[114] & ~t[115]) | (~t[109] & t[110] & t[111] & t[112] & ~t[115]) | (~t[109] & t[110] & t[113] & t[114] & ~t[115]) | (t[109] & ~t[111] & ~t[113] & t[115]) | (~t[109] & t[111] & t[113] & t[115]);
  assign t[92] = (t[109] & t[110] & ~t[111] & ~t[113] & t[114] & ~t[115]) | (t[109] & t[111] & ~t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & t[113] & ~t[114] & ~t[115]) | (~t[109] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[109] & ~t[110] & ~t[112] & t[113] & ~t[115]) | (~t[109] & ~t[111] & t[112] & t[113] & t[114]) | (t[112] & t[113] & ~t[114] & ~t[115]);
  assign t[93] = (t[116] & ~t[118] & ~t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[119] & ~t[120] & ~t[122]) | (t[116] & ~t[117] & ~t[118] & ~t[121] & ~t[122]) | (~t[116] & t[117] & t[118] & t[119] & ~t[122]) | (~t[116] & t[117] & t[120] & t[121] & ~t[122]) | (t[116] & ~t[118] & ~t[120] & t[122]) | (~t[116] & t[118] & t[120] & t[122]);
  assign t[94] = (t[116] & t[117] & ~t[118] & t[119] & ~t[120] & ~t[122]) | (t[116] & ~t[118] & ~t[119] & t[120] & ~t[121] & t[122]) | (~t[117] & t[118] & ~t[119] & ~t[120] & ~t[122]) | (~t[116] & t[118] & ~t[119] & ~t[120] & ~t[121]) | (~t[116] & ~t[117] & t[118] & ~t[121] & ~t[122]) | (~t[116] & t[118] & t[119] & ~t[120] & t[121]) | (t[118] & ~t[119] & t[121] & ~t[122]);
  assign t[95] = (t[117] & ~t[118] & ~t[119] & ~t[120] & ~t[121]) | (~t[116] & t[117] & ~t[119] & ~t[120] & ~t[122]) | (~t[116] & t[117] & ~t[118] & ~t[121] & ~t[122]) | (t[116] & ~t[117] & t[118] & t[119] & ~t[122]) | (t[116] & ~t[117] & t[120] & t[121] & ~t[122]) | (t[117] & ~t[119] & ~t[121] & t[122]) | (~t[117] & t[119] & t[121] & t[122]);
  assign t[96] = (t[116] & t[117] & t[118] & ~t[119] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & ~t[119] & ~t[120] & t[121] & t[122]) | (~t[117] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (~t[116] & ~t[118] & t[119] & ~t[121] & ~t[122]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[122]) | (~t[117] & t[118] & t[119] & t[120] & ~t[121]) | (~t[118] & t[119] & t[120] & ~t[122]);
  assign t[97] = (t[116] & t[117] & ~t[118] & ~t[120] & t[121] & ~t[122]) | (t[116] & t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[122]) | (~t[116] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[116] & ~t[117] & ~t[119] & t[120] & ~t[122]) | (~t[116] & ~t[118] & t[119] & t[120] & t[121]) | (t[119] & t[120] & ~t[121] & ~t[122]);
  assign t[98] = (t[116] & t[117] & ~t[119] & t[120] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[119] & ~t[120] & t[121] & ~t[122]) | (~t[116] & ~t[117] & ~t[118] & t[121] & ~t[122]) | (~t[117] & t[118] & ~t[119] & t[120] & t[121]) | (t[118] & ~t[120] & t[121] & ~t[122]);
  assign t[99] = (t[123] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[124] & ~t[125] & ~t[128] & ~t[129]) | (~t[123] & t[124] & t[125] & t[126] & ~t[129]) | (~t[123] & t[124] & t[127] & t[128] & ~t[129]) | (t[123] & ~t[125] & ~t[127] & t[129]) | (~t[123] & t[125] & t[127] & t[129]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[53]) | (~t[0] & t[37] & ~t[53]) | (~t[0] & ~t[37] & t[53]) | (t[0] & t[37] & t[53]);
endmodule

module R2ind64(x, y);
 input [36:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[107] & t[108] & ~t[109] & t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[109] & ~t[110] & t[111] & ~t[112] & t[113]) | (~t[108] & t[109] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[108] & t[109] & ~t[112] & ~t[113]) | (~t[107] & t[109] & t[110] & ~t[111] & t[112]) | (t[109] & ~t[110] & t[112] & ~t[113]);
  assign t[104] = (t[108] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & t[108] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[108] & ~t[109] & ~t[112] & ~t[113]) | (t[107] & ~t[108] & t[109] & t[110] & ~t[113]) | (t[107] & ~t[108] & t[111] & t[112] & ~t[113]) | (t[108] & ~t[110] & ~t[112] & t[113]) | (~t[108] & t[110] & t[112] & t[113]);
  assign t[105] = (t[107] & t[108] & t[109] & ~t[110] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[110] & ~t[111] & t[112] & t[113]) | (~t[108] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[109] & t[110] & ~t[112] & ~t[113]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[113]) | (~t[108] & t[109] & t[110] & t[111] & ~t[112]) | (~t[109] & t[110] & t[111] & ~t[113]);
  assign t[106] = (t[107] & t[108] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[107] & ~t[108] & ~t[109] & t[112] & ~t[113]) | (~t[108] & t[109] & ~t[110] & t[111] & t[112]) | (t[109] & ~t[111] & t[112] & ~t[113]);
  assign t[107] = t[128] ^ x[7];
  assign t[108] = t[129] ^ x[34];
  assign t[109] = t[130] ^ x[32];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[35];
  assign t[111] = t[132] ^ x[8];
  assign t[112] = t[133] ^ x[36];
  assign t[113] = t[134] ^ x[6];
  assign t[114] = t[135] ^ x[14];
  assign t[115] = t[136] ^ x[16];
  assign t[116] = t[137] ^ x[15];
  assign t[117] = t[138] ^ x[17];
  assign t[118] = t[139] ^ x[18];
  assign t[119] = t[140] ^ x[19];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[13];
  assign t[121] = t[142] ^ x[25];
  assign t[122] = t[143] ^ x[27];
  assign t[123] = t[144] ^ x[26];
  assign t[124] = t[145] ^ x[28];
  assign t[125] = t[146] ^ x[29];
  assign t[126] = t[147] ^ x[30];
  assign t[127] = t[148] ^ x[24];
  assign t[128] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[129] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[131] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[132] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[133] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[134] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[135] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[136] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[137] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[138] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[139] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[141] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[142] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[143] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[144] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[145] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[146] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[147] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[148] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[62]);
  assign t[15] = ~(t[61] ^ t[14]);
  assign t[16] = t[63] ^ t[62];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[61] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[61] ^ t[27];
  assign t[23] = t[64] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[62] ^ t[65];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[66]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[64] ^ t[29]);
  assign t[31] = t[67] ^ t[66];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[64] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[64] ^ t[36];
  assign t[36] = t[66] ^ t[68];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[69]);
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~t[46];
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~(t[49] ^ t[50]);
  assign t[47] = t[16] ^ t[21];
  assign t[48] = t[61] ^ t[14];
  assign t[49] = t[51] ^ t[24];
  assign t[4] = ~(t[7] ^ t[60]);
  assign t[50] = t[18] ^ t[52];
  assign t[51] = t[31] ^ t[34];
  assign t[52] = t[64] ^ t[29];
  assign t[53] = x[0] ? x[33] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~t[57];
  assign t[56] = ~(t[44]);
  assign t[57] = ~(t[58] ^ t[70]);
  assign t[58] = ~t[59];
  assign t[59] = ~(t[49]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[61] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[62] = (t[73] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[73] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[63] = (t[73] & ~t[77]) | (~t[73] & t[77]);
  assign t[64] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[65] = (t[73] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[73] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[66] = (t[79] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[79] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[67] = (t[79] & ~t[83]) | (~t[79] & t[83]);
  assign t[68] = (t[79] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[79] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[69] = (t[71] & ~t[85]) | (~t[71] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[71] & ~t[87] & ~t[72]) | (~t[86] & t[87] & ~t[88]) | (~t[71] & ~t[87] & t[72]) | (t[86] & t[87] & t[88]);
  assign t[71] = t[89] ^ x[7];
  assign t[72] = t[90] ^ x[8];
  assign t[73] = t[91] ^ x[14];
  assign t[74] = t[92] ^ x[15];
  assign t[75] = t[93] ^ x[16];
  assign t[76] = t[94] ^ x[17];
  assign t[77] = t[95] ^ x[18];
  assign t[78] = t[96] ^ x[19];
  assign t[79] = t[97] ^ x[25];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[26];
  assign t[81] = t[99] ^ x[27];
  assign t[82] = t[100] ^ x[28];
  assign t[83] = t[101] ^ x[29];
  assign t[84] = t[102] ^ x[30];
  assign t[85] = t[103] ^ x[32];
  assign t[86] = t[104] ^ x[34];
  assign t[87] = t[105] ^ x[35];
  assign t[88] = t[106] ^ x[36];
  assign t[89] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[8] = t[61] & t[13];
  assign t[90] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[91] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[92] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[93] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[94] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[95] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[96] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[97] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[98] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[53]) | (~t[0] & t[37] & ~t[53]) | (~t[0] & ~t[37] & t[53]) | (t[0] & t[37] & t[53]);
endmodule

module R2ind65(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[19];
  assign t[102] = t[123] ^ x[20];
  assign t[103] = t[124] ^ x[14];
  assign t[104] = t[125] ^ x[26];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[27];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[30];
  assign t[109] = t[130] ^ x[31];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[25];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[119] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[121] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[122] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[123] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[124] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[125] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[126] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[127] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[128] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[129] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[131] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[48]);
  assign t[15] = ~(t[47] ^ t[14]);
  assign t[16] = t[49] ^ t[48];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[47] ^ t[27];
  assign t[23] = t[50] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[48] ^ t[51];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[52]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[50] ^ t[29]);
  assign t[31] = t[53] ^ t[52];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[50] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[50] ^ t[36];
  assign t[36] = t[52] ^ t[54];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[27] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[36] ^ t[24];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[58] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[49] = (t[58] & ~t[62]) | (~t[58] & t[62]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[58] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[52] = (t[64] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[64] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[64] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[57]) | (~t[56] & ~t[71] & t[72]) | (t[70] & t[71] & t[57]);
  assign t[56] = t[73] ^ x[8];
  assign t[57] = t[74] ^ x[9];
  assign t[58] = t[75] ^ x[15];
  assign t[59] = t[76] ^ x[16];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[17];
  assign t[61] = t[78] ^ x[18];
  assign t[62] = t[79] ^ x[19];
  assign t[63] = t[80] ^ x[20];
  assign t[64] = t[81] ^ x[26];
  assign t[65] = t[82] ^ x[27];
  assign t[66] = t[83] ^ x[28];
  assign t[67] = t[84] ^ x[29];
  assign t[68] = t[85] ^ x[30];
  assign t[69] = t[86] ^ x[31];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[33];
  assign t[71] = t[88] ^ x[34];
  assign t[72] = t[89] ^ x[35];
  assign t[73] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[86] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[87] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[88] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[47] & t[13];
  assign t[90] = t[111] ^ x[8];
  assign t[91] = t[112] ^ x[33];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[9];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[15];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[16];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind66(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[20];
  assign t[105] = t[126] ^ x[14];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[31];
  assign t[112] = t[133] ^ x[25];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[121] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[122] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[123] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[126] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[127] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[128] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[129] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[132] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[133] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[50]);
  assign t[15] = ~(t[49] ^ t[14]);
  assign t[16] = t[51] ^ t[50];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[49] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[49] ^ t[27];
  assign t[23] = t[52] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[50] ^ t[53];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[54]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[52] ^ t[29]);
  assign t[31] = t[55] ^ t[54];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[52] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[52] ^ t[36];
  assign t[36] = t[54] ^ t[56];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[57]);
  assign t[42] = t[44] ^ t[9];
  assign t[43] = ~t[45];
  assign t[44] = t[16] ^ t[21];
  assign t[45] = ~(t[46]);
  assign t[46] = t[47] ^ t[24];
  assign t[47] = t[31] ^ t[34];
  assign t[48] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[49] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[60] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[60] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[51] = (t[60] & ~t[64]) | (~t[60] & t[64]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[60] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[60] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[54] = (t[66] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[66] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[55] = (t[66] & ~t[70]) | (~t[66] & t[70]);
  assign t[56] = (t[66] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[66] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[57] = (t[58] & ~t[73] & ~t[59]) | (~t[72] & t[73] & ~t[74]) | (~t[58] & ~t[73] & t[59]) | (t[72] & t[73] & t[74]);
  assign t[58] = t[75] ^ x[8];
  assign t[59] = t[76] ^ x[9];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[15];
  assign t[61] = t[78] ^ x[16];
  assign t[62] = t[79] ^ x[17];
  assign t[63] = t[80] ^ x[18];
  assign t[64] = t[81] ^ x[19];
  assign t[65] = t[82] ^ x[20];
  assign t[66] = t[83] ^ x[26];
  assign t[67] = t[84] ^ x[27];
  assign t[68] = t[85] ^ x[28];
  assign t[69] = t[86] ^ x[29];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[30];
  assign t[71] = t[88] ^ x[31];
  assign t[72] = t[89] ^ x[33];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[35];
  assign t[75] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[76] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[77] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[8] = t[49] & t[13];
  assign t[90] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[7];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind67(x, y);
 input [35:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[14];
  assign t[101] = t[122] ^ x[17];
  assign t[102] = t[123] ^ x[15];
  assign t[103] = t[124] ^ x[18];
  assign t[104] = t[125] ^ x[16];
  assign t[105] = t[126] ^ x[19];
  assign t[106] = t[127] ^ x[13];
  assign t[107] = t[128] ^ x[25];
  assign t[108] = t[129] ^ x[28];
  assign t[109] = t[130] ^ x[26];
  assign t[10] = t[16] ^ t[17];
  assign t[110] = t[131] ^ x[29];
  assign t[111] = t[132] ^ x[27];
  assign t[112] = t[133] ^ x[30];
  assign t[113] = t[134] ^ x[24];
  assign t[114] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[115] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[116] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[117] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[118] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[119] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[121] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[122] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[123] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[124] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[125] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[126] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[127] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[128] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[129] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[131] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[132] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[133] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[134] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[48] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[49] ^ t[50];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[50]);
  assign t[19] = ~(t[48] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[48] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[51] ^ t[29];
  assign t[25] = t[48] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[52] ^ t[53];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[53]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[51] ^ t[29]);
  assign t[31] = t[51] & t[35];
  assign t[32] = t[50] ^ t[54];
  assign t[33] = t[48] ^ t[16];
  assign t[34] = t[51] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[53] ^ t[55];
  assign t[37] = t[51] ^ t[27];
  assign t[38] = x[0] ? x[31] : t[39];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5]);
  assign t[40] = ~t[42];
  assign t[41] = ~(t[43]);
  assign t[42] = ~(t[44] ^ t[56]);
  assign t[43] = t[32] ^ t[11];
  assign t[44] = ~t[45];
  assign t[45] = ~(t[46]);
  assign t[46] = t[36] ^ t[22];
  assign t[47] = (t[57] & ~t[58]) | (~t[57] & t[58]);
  assign t[48] = (t[59] & ~t[60]) | (~t[59] & t[60]);
  assign t[49] = (t[59] & ~t[61]) | (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[47]);
  assign t[50] = (t[59] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[61]) | (~t[59] & ~t[63] & t[64]) | (t[62] & t[63] & t[61]);
  assign t[51] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[52] = (t[65] & ~t[67]) | (~t[65] & t[67]);
  assign t[53] = (t[65] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[67]) | (~t[65] & ~t[69] & t[70]) | (t[68] & t[69] & t[67]);
  assign t[54] = (t[59] & ~t[63] & ~t[61]) | (~t[62] & t[63] & ~t[64]) | (~t[59] & ~t[63] & t[61]) | (t[62] & t[63] & t[64]);
  assign t[55] = (t[65] & ~t[69] & ~t[67]) | (~t[68] & t[69] & ~t[70]) | (~t[65] & ~t[69] & t[67]) | (t[68] & t[69] & t[70]);
  assign t[56] = (t[57] & ~t[72] & ~t[74]) | (~t[71] & t[72] & ~t[73]) | (~t[57] & ~t[72] & t[74]) | (t[71] & t[72] & t[73]);
  assign t[57] = t[75] ^ x[7];
  assign t[58] = t[76] ^ x[8];
  assign t[59] = t[77] ^ x[14];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[16];
  assign t[62] = t[80] ^ x[17];
  assign t[63] = t[81] ^ x[18];
  assign t[64] = t[82] ^ x[19];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[26];
  assign t[67] = t[85] ^ x[27];
  assign t[68] = t[86] ^ x[28];
  assign t[69] = t[87] ^ x[29];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = t[89] ^ x[32];
  assign t[72] = t[90] ^ x[33];
  assign t[73] = t[91] ^ x[34];
  assign t[74] = t[92] ^ x[35];
  assign t[75] = (t[93] & ~t[95] & ~t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[96] & ~t[97] & ~t[99]) | (t[93] & ~t[94] & ~t[95] & ~t[98] & ~t[99]) | (~t[93] & t[94] & t[95] & t[96] & ~t[99]) | (~t[93] & t[94] & t[97] & t[98] & ~t[99]) | (t[93] & ~t[95] & ~t[97] & t[99]) | (~t[93] & t[95] & t[97] & t[99]);
  assign t[76] = (t[93] & t[94] & ~t[95] & t[96] & ~t[97] & ~t[99]) | (t[93] & ~t[95] & ~t[96] & t[97] & ~t[98] & t[99]) | (~t[94] & t[95] & ~t[96] & ~t[97] & ~t[99]) | (~t[93] & t[95] & ~t[96] & ~t[97] & ~t[98]) | (~t[93] & ~t[94] & t[95] & ~t[98] & ~t[99]) | (~t[93] & t[95] & t[96] & ~t[97] & t[98]) | (t[95] & ~t[96] & t[98] & ~t[99]);
  assign t[77] = (t[100] & ~t[102] & ~t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[103] & ~t[104] & ~t[106]) | (t[100] & ~t[101] & ~t[102] & ~t[105] & ~t[106]) | (~t[100] & t[101] & t[102] & t[103] & ~t[106]) | (~t[100] & t[101] & t[104] & t[105] & ~t[106]) | (t[100] & ~t[102] & ~t[104] & t[106]) | (~t[100] & t[102] & t[104] & t[106]);
  assign t[78] = (t[100] & t[101] & ~t[102] & t[103] & ~t[104] & ~t[106]) | (t[100] & ~t[102] & ~t[103] & t[104] & ~t[105] & t[106]) | (~t[101] & t[102] & ~t[103] & ~t[104] & ~t[106]) | (~t[100] & t[102] & ~t[103] & ~t[104] & ~t[105]) | (~t[100] & ~t[101] & t[102] & ~t[105] & ~t[106]) | (~t[100] & t[102] & t[103] & ~t[104] & t[105]) | (t[102] & ~t[103] & t[105] & ~t[106]);
  assign t[79] = (t[100] & t[101] & ~t[102] & ~t[104] & t[105] & ~t[106]) | (t[100] & t[102] & ~t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[102] & t[104] & ~t[105] & ~t[106]) | (~t[100] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[100] & ~t[101] & ~t[103] & t[104] & ~t[106]) | (~t[100] & ~t[102] & t[103] & t[104] & t[105]) | (t[103] & t[104] & ~t[105] & ~t[106]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (t[101] & ~t[102] & ~t[103] & ~t[104] & ~t[105]) | (~t[100] & t[101] & ~t[103] & ~t[104] & ~t[106]) | (~t[100] & t[101] & ~t[102] & ~t[105] & ~t[106]) | (t[100] & ~t[101] & t[102] & t[103] & ~t[106]) | (t[100] & ~t[101] & t[104] & t[105] & ~t[106]) | (t[101] & ~t[103] & ~t[105] & t[106]) | (~t[101] & t[103] & t[105] & t[106]);
  assign t[81] = (t[100] & t[101] & t[102] & ~t[103] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & ~t[103] & ~t[104] & t[105] & t[106]) | (~t[101] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (~t[100] & ~t[102] & t[103] & ~t[105] & ~t[106]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[106]) | (~t[101] & t[102] & t[103] & t[104] & ~t[105]) | (~t[102] & t[103] & t[104] & ~t[106]);
  assign t[82] = (t[100] & t[101] & ~t[103] & t[104] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[103] & ~t[104] & t[105] & ~t[106]) | (~t[100] & ~t[101] & ~t[102] & t[105] & ~t[106]) | (~t[101] & t[102] & ~t[103] & t[104] & t[105]) | (t[102] & ~t[104] & t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[84] = (t[107] & t[108] & ~t[109] & t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[109] & ~t[110] & t[111] & ~t[112] & t[113]) | (~t[108] & t[109] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[108] & t[109] & ~t[112] & ~t[113]) | (~t[107] & t[109] & t[110] & ~t[111] & t[112]) | (t[109] & ~t[110] & t[112] & ~t[113]);
  assign t[85] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[86] = (t[108] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & t[108] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[108] & ~t[109] & ~t[112] & ~t[113]) | (t[107] & ~t[108] & t[109] & t[110] & ~t[113]) | (t[107] & ~t[108] & t[111] & t[112] & ~t[113]) | (t[108] & ~t[110] & ~t[112] & t[113]) | (~t[108] & t[110] & t[112] & t[113]);
  assign t[87] = (t[107] & t[108] & t[109] & ~t[110] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[110] & ~t[111] & t[112] & t[113]) | (~t[108] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[109] & t[110] & ~t[112] & ~t[113]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[113]) | (~t[108] & t[109] & t[110] & t[111] & ~t[112]) | (~t[109] & t[110] & t[111] & ~t[113]);
  assign t[88] = (t[107] & t[108] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[107] & ~t[108] & ~t[109] & t[112] & ~t[113]) | (~t[108] & t[109] & ~t[110] & t[111] & t[112]) | (t[109] & ~t[111] & t[112] & ~t[113]);
  assign t[89] = (t[94] & ~t[95] & ~t[96] & ~t[97] & ~t[98]) | (~t[93] & t[94] & ~t[96] & ~t[97] & ~t[99]) | (~t[93] & t[94] & ~t[95] & ~t[98] & ~t[99]) | (t[93] & ~t[94] & t[95] & t[96] & ~t[99]) | (t[93] & ~t[94] & t[97] & t[98] & ~t[99]) | (t[94] & ~t[96] & ~t[98] & t[99]) | (~t[94] & t[96] & t[98] & t[99]);
  assign t[8] = t[12] ^ t[13];
  assign t[90] = (t[93] & t[94] & t[95] & ~t[96] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & ~t[96] & ~t[97] & t[98] & t[99]) | (~t[94] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (~t[93] & ~t[95] & t[96] & ~t[98] & ~t[99]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[99]) | (~t[94] & t[95] & t[96] & t[97] & ~t[98]) | (~t[95] & t[96] & t[97] & ~t[99]);
  assign t[91] = (t[93] & t[94] & ~t[95] & ~t[97] & t[98] & ~t[99]) | (t[93] & t[95] & ~t[96] & ~t[97] & ~t[98] & t[99]) | (~t[94] & ~t[95] & t[97] & ~t[98] & ~t[99]) | (~t[93] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[93] & ~t[94] & ~t[96] & t[97] & ~t[99]) | (~t[93] & ~t[95] & t[96] & t[97] & t[98]) | (t[96] & t[97] & ~t[98] & ~t[99]);
  assign t[92] = (t[93] & t[94] & ~t[96] & t[97] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & t[96] & ~t[97] & ~t[98] & t[99]) | (~t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[96] & ~t[97] & t[98] & ~t[99]) | (~t[93] & ~t[94] & ~t[95] & t[98] & ~t[99]) | (~t[94] & t[95] & ~t[96] & t[97] & t[98]) | (t[95] & ~t[97] & t[98] & ~t[99]);
  assign t[93] = t[114] ^ x[7];
  assign t[94] = t[115] ^ x[32];
  assign t[95] = t[116] ^ x[8];
  assign t[96] = t[117] ^ x[33];
  assign t[97] = t[118] ^ x[34];
  assign t[98] = t[119] ^ x[35];
  assign t[99] = t[120] ^ x[6];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0] & ~t[38]) | (~t[0] & t[38]);
endmodule

module R2ind68(x, y);
 input [35:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[15];
  assign t[101] = t[122] ^ x[18];
  assign t[102] = t[123] ^ x[16];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[13];
  assign t[105] = t[126] ^ x[25];
  assign t[106] = t[127] ^ x[28];
  assign t[107] = t[128] ^ x[26];
  assign t[108] = t[129] ^ x[29];
  assign t[109] = t[130] ^ x[27];
  assign t[10] = t[16] ^ t[17];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[24];
  assign t[112] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[113] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[114] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[115] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[116] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[117] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[118] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[119] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[121] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[122] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[123] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[124] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[125] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[126] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[127] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[128] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[129] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[131] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[132] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[46] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[47] ^ t[48];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[48]);
  assign t[19] = ~(t[46] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[46] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[49] ^ t[29];
  assign t[25] = t[46] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[50] ^ t[51];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[51]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[49] ^ t[29]);
  assign t[31] = t[49] & t[35];
  assign t[32] = t[48] ^ t[52];
  assign t[33] = t[46] ^ t[16];
  assign t[34] = t[49] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[51] ^ t[53];
  assign t[37] = t[49] ^ t[27];
  assign t[38] = x[0] ? x[31] : t[39];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5]);
  assign t[40] = ~t[42];
  assign t[41] = ~(t[7]);
  assign t[42] = ~(t[43] ^ t[54]);
  assign t[43] = ~t[44];
  assign t[44] = ~(t[14]);
  assign t[45] = (t[55] & ~t[56]) | (~t[55] & t[56]);
  assign t[46] = (t[57] & ~t[58]) | (~t[57] & t[58]);
  assign t[47] = (t[57] & ~t[59]) | (~t[57] & t[59]);
  assign t[48] = (t[57] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[59]) | (~t[57] & ~t[61] & t[62]) | (t[60] & t[61] & t[59]);
  assign t[49] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[4] = ~(t[6] ^ t[45]);
  assign t[50] = (t[63] & ~t[65]) | (~t[63] & t[65]);
  assign t[51] = (t[63] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[65]) | (~t[63] & ~t[67] & t[68]) | (t[66] & t[67] & t[65]);
  assign t[52] = (t[57] & ~t[61] & ~t[59]) | (~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[61] & t[59]) | (t[60] & t[61] & t[62]);
  assign t[53] = (t[63] & ~t[67] & ~t[65]) | (~t[66] & t[67] & ~t[68]) | (~t[63] & ~t[67] & t[65]) | (t[66] & t[67] & t[68]);
  assign t[54] = (t[55] & ~t[70] & ~t[71]) | (~t[69] & t[70] & ~t[72]) | (~t[55] & ~t[70] & t[71]) | (t[69] & t[70] & t[72]);
  assign t[55] = t[73] ^ x[7];
  assign t[56] = t[74] ^ x[8];
  assign t[57] = t[75] ^ x[14];
  assign t[58] = t[76] ^ x[15];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = t[78] ^ x[17];
  assign t[61] = t[79] ^ x[18];
  assign t[62] = t[80] ^ x[19];
  assign t[63] = t[81] ^ x[25];
  assign t[64] = t[82] ^ x[26];
  assign t[65] = t[83] ^ x[27];
  assign t[66] = t[84] ^ x[28];
  assign t[67] = t[85] ^ x[29];
  assign t[68] = t[86] ^ x[30];
  assign t[69] = t[87] ^ x[32];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[33];
  assign t[71] = t[89] ^ x[34];
  assign t[72] = t[90] ^ x[35];
  assign t[73] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[74] = (t[91] & t[92] & ~t[93] & t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[93] & ~t[94] & t[95] & ~t[96] & t[97]) | (~t[92] & t[93] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[92] & t[93] & ~t[96] & ~t[97]) | (~t[91] & t[93] & t[94] & ~t[95] & t[96]) | (t[93] & ~t[94] & t[96] & ~t[97]);
  assign t[75] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[76] = (t[98] & t[99] & ~t[100] & t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[100] & ~t[101] & t[102] & ~t[103] & t[104]) | (~t[99] & t[100] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[99] & t[100] & ~t[103] & ~t[104]) | (~t[98] & t[100] & t[101] & ~t[102] & t[103]) | (t[100] & ~t[101] & t[103] & ~t[104]);
  assign t[77] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[78] = (t[99] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & t[99] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[99] & ~t[100] & ~t[103] & ~t[104]) | (t[98] & ~t[99] & t[100] & t[101] & ~t[104]) | (t[98] & ~t[99] & t[102] & t[103] & ~t[104]) | (t[99] & ~t[101] & ~t[103] & t[104]) | (~t[99] & t[101] & t[103] & t[104]);
  assign t[79] = (t[98] & t[99] & t[100] & ~t[101] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[101] & ~t[102] & t[103] & t[104]) | (~t[99] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[100] & t[101] & ~t[103] & ~t[104]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[104]) | (~t[99] & t[100] & t[101] & t[102] & ~t[103]) | (~t[100] & t[101] & t[102] & ~t[104]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (t[98] & t[99] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[98] & ~t[99] & ~t[100] & t[103] & ~t[104]) | (~t[99] & t[100] & ~t[101] & t[102] & t[103]) | (t[100] & ~t[102] & t[103] & ~t[104]);
  assign t[81] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[82] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[83] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[84] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[85] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[86] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[87] = (t[92] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & t[92] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[92] & ~t[93] & ~t[96] & ~t[97]) | (t[91] & ~t[92] & t[93] & t[94] & ~t[97]) | (t[91] & ~t[92] & t[95] & t[96] & ~t[97]) | (t[92] & ~t[94] & ~t[96] & t[97]) | (~t[92] & t[94] & t[96] & t[97]);
  assign t[88] = (t[91] & t[92] & t[93] & ~t[94] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[94] & ~t[95] & t[96] & t[97]) | (~t[92] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[93] & t[94] & ~t[96] & ~t[97]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[97]) | (~t[92] & t[93] & t[94] & t[95] & ~t[96]) | (~t[93] & t[94] & t[95] & ~t[97]);
  assign t[89] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[8] = t[12] ^ t[13];
  assign t[90] = (t[91] & t[92] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[91] & ~t[92] & ~t[93] & t[96] & ~t[97]) | (~t[92] & t[93] & ~t[94] & t[95] & t[96]) | (t[93] & ~t[95] & t[96] & ~t[97]);
  assign t[91] = t[112] ^ x[7];
  assign t[92] = t[113] ^ x[32];
  assign t[93] = t[114] ^ x[8];
  assign t[94] = t[115] ^ x[33];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[35];
  assign t[97] = t[118] ^ x[6];
  assign t[98] = t[119] ^ x[14];
  assign t[99] = t[120] ^ x[17];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0] & ~t[38]) | (~t[0] & t[38]);
endmodule

module R2ind69(x, y);
 input [35:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[101] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[102] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[103] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[104] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[105] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[35]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[114] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[115] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[116] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[118] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[119] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[11] = ~(t[37] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[38] ^ t[39];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = x[0] ? x[35] : t[18];
  assign t[18] = ~(t[19] ^ t[20]);
  assign t[19] = ~t[21];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[23] ^ t[41]);
  assign t[22] = t[24] ^ t[8];
  assign t[23] = ~t[25];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = ~(t[28]);
  assign t[26] = t[42] ^ t[35];
  assign t[27] = t[10] & t[29];
  assign t[28] = t[30] ^ t[14];
  assign t[29] = t[37] ^ t[7];
  assign t[2] = ~t[4];
  assign t[30] = t[31] ^ t[32];
  assign t[31] = t[43] ^ t[38];
  assign t[32] = t[15] & t[33];
  assign t[33] = t[40] ^ t[13];
  assign t[34] = (t[44] & ~t[46] & ~t[48]) | (~t[45] & t[46] & ~t[47]) | (~t[44] & ~t[46] & t[48]) | (t[45] & t[46] & t[47]);
  assign t[35] = (t[49] & ~t[51] & ~t[53]) | (~t[50] & t[51] & ~t[52]) | (~t[49] & ~t[51] & t[53]) | (t[50] & t[51] & t[52]);
  assign t[36] = (t[49] & ~t[51] & ~t[52]) | (~t[50] & t[51] & ~t[53]) | (~t[49] & ~t[51] & t[52]) | (t[50] & t[51] & t[53]);
  assign t[37] = (t[49] & ~t[54]) | (~t[49] & t[54]);
  assign t[38] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[39] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[60]) | (~t[55] & t[60]);
  assign t[41] = (t[44] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[44] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[42] = (t[49] & ~t[52]) | (~t[49] & t[52]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = t[61] ^ x[8];
  assign t[45] = t[62] ^ x[9];
  assign t[46] = t[63] ^ x[10];
  assign t[47] = t[64] ^ x[11];
  assign t[48] = t[65] ^ x[12];
  assign t[49] = t[66] ^ x[18];
  assign t[4] = ~(t[6] ^ t[34]);
  assign t[50] = t[67] ^ x[19];
  assign t[51] = t[68] ^ x[20];
  assign t[52] = t[69] ^ x[21];
  assign t[53] = t[70] ^ x[22];
  assign t[54] = t[71] ^ x[23];
  assign t[55] = t[72] ^ x[29];
  assign t[56] = t[73] ^ x[30];
  assign t[57] = t[74] ^ x[31];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[34];
  assign t[61] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[62] = (t[79] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (~t[78] & t[79] & ~t[81] & ~t[82] & ~t[84]) | (~t[78] & t[79] & ~t[80] & ~t[83] & ~t[84]) | (t[78] & ~t[79] & t[80] & t[81] & ~t[84]) | (t[78] & ~t[79] & t[82] & t[83] & ~t[84]) | (t[79] & ~t[81] & ~t[83] & t[84]) | (~t[79] & t[81] & t[83] & t[84]);
  assign t[63] = (t[78] & t[79] & t[80] & ~t[81] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & ~t[81] & ~t[82] & t[83] & t[84]) | (~t[79] & ~t[80] & t[81] & ~t[82] & ~t[83]) | (~t[78] & ~t[80] & t[81] & ~t[83] & ~t[84]) | (~t[78] & ~t[79] & t[81] & ~t[82] & ~t[84]) | (~t[79] & t[80] & t[81] & t[82] & ~t[83]) | (~t[80] & t[81] & t[82] & ~t[84]);
  assign t[64] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[65] = (t[78] & t[79] & ~t[81] & t[82] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & ~t[81] & ~t[82] & t[83]) | (~t[78] & ~t[81] & ~t[82] & t[83] & ~t[84]) | (~t[78] & ~t[79] & ~t[80] & t[83] & ~t[84]) | (~t[79] & t[80] & ~t[81] & t[82] & t[83]) | (t[80] & ~t[82] & t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = ~t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[72] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[73] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[74] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[8];
  assign t[79] = t[100] ^ x[9];
  assign t[7] = t[35] ^ t[36];
  assign t[80] = t[101] ^ x[6];
  assign t[81] = t[102] ^ x[10];
  assign t[82] = t[103] ^ x[11];
  assign t[83] = t[104] ^ x[12];
  assign t[84] = t[105] ^ x[7];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[23];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[29];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[32];
  assign t[97] = t[118] ^ x[33];
  assign t[98] = t[119] ^ x[28];
  assign t[99] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~t[17]) | (~t[0] & t[17]);
endmodule

module R2ind70(x, y);
 input [36:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[101] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[102] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[103] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[104] = (t[108] & t[109] & ~t[110] & t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[110] & ~t[111] & t[112] & ~t[113] & t[114]) | (~t[109] & t[110] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[109] & t[110] & ~t[113] & ~t[114]) | (~t[108] & t[110] & t[111] & ~t[112] & t[113]) | (t[110] & ~t[111] & t[113] & ~t[114]);
  assign t[105] = (t[109] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & t[109] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[109] & ~t[110] & ~t[113] & ~t[114]) | (t[108] & ~t[109] & t[110] & t[111] & ~t[114]) | (t[108] & ~t[109] & t[112] & t[113] & ~t[114]) | (t[109] & ~t[111] & ~t[113] & t[114]) | (~t[109] & t[111] & t[113] & t[114]);
  assign t[106] = (t[108] & t[109] & t[110] & ~t[111] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[111] & ~t[112] & t[113] & t[114]) | (~t[109] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[110] & t[111] & ~t[113] & ~t[114]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[114]) | (~t[109] & t[110] & t[111] & t[112] & ~t[113]) | (~t[110] & t[111] & t[112] & ~t[114]);
  assign t[107] = (t[108] & t[109] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[108] & ~t[109] & ~t[110] & t[113] & ~t[114]) | (~t[109] & t[110] & ~t[111] & t[112] & t[113]) | (t[110] & ~t[112] & t[113] & ~t[114]);
  assign t[108] = t[129] ^ x[7];
  assign t[109] = t[130] ^ x[34];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[32];
  assign t[111] = t[132] ^ x[35];
  assign t[112] = t[133] ^ x[8];
  assign t[113] = t[134] ^ x[36];
  assign t[114] = t[135] ^ x[6];
  assign t[115] = t[136] ^ x[14];
  assign t[116] = t[137] ^ x[16];
  assign t[117] = t[138] ^ x[15];
  assign t[118] = t[139] ^ x[17];
  assign t[119] = t[140] ^ x[18];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[19];
  assign t[121] = t[142] ^ x[13];
  assign t[122] = t[143] ^ x[25];
  assign t[123] = t[144] ^ x[27];
  assign t[124] = t[145] ^ x[26];
  assign t[125] = t[146] ^ x[28];
  assign t[126] = t[147] ^ x[29];
  assign t[127] = t[148] ^ x[30];
  assign t[128] = t[149] ^ x[24];
  assign t[129] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[131] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[132] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[133] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[134] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[135] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[136] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[137] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[138] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[139] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[141] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[142] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[143] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[144] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[145] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[146] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[147] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[148] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[149] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[63]);
  assign t[15] = ~(t[62] ^ t[14]);
  assign t[16] = t[64] ^ t[63];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[62] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[62] ^ t[27];
  assign t[23] = t[65] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[63] ^ t[66];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[67]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[65] ^ t[29]);
  assign t[31] = t[68] ^ t[67];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[65] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[65] ^ t[36];
  assign t[36] = t[67] ^ t[69];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[70]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[62] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[61]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[65] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[71]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[62] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[63] = (t[74] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[74] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[64] = (t[74] & ~t[78]) | (~t[74] & t[78]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[74] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[74] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[67] = (t[80] & ~t[83] & ~t[85]) | (~t[82] & t[83] & ~t[84]) | (~t[80] & ~t[83] & t[85]) | (t[82] & t[83] & t[84]);
  assign t[68] = (t[80] & ~t[84]) | (~t[80] & t[84]);
  assign t[69] = (t[80] & ~t[83] & ~t[84]) | (~t[82] & t[83] & ~t[85]) | (~t[80] & ~t[83] & t[84]) | (t[82] & t[83] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[72] & ~t[86]) | (~t[72] & t[86]);
  assign t[71] = (t[72] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[73]) | (~t[72] & ~t[88] & t[89]) | (t[87] & t[88] & t[73]);
  assign t[72] = t[90] ^ x[7];
  assign t[73] = t[91] ^ x[8];
  assign t[74] = t[92] ^ x[14];
  assign t[75] = t[93] ^ x[15];
  assign t[76] = t[94] ^ x[16];
  assign t[77] = t[95] ^ x[17];
  assign t[78] = t[96] ^ x[18];
  assign t[79] = t[97] ^ x[19];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[25];
  assign t[81] = t[99] ^ x[26];
  assign t[82] = t[100] ^ x[27];
  assign t[83] = t[101] ^ x[28];
  assign t[84] = t[102] ^ x[29];
  assign t[85] = t[103] ^ x[30];
  assign t[86] = t[104] ^ x[32];
  assign t[87] = t[105] ^ x[34];
  assign t[88] = t[106] ^ x[35];
  assign t[89] = t[107] ^ x[36];
  assign t[8] = t[62] & t[13];
  assign t[90] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[91] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[92] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[93] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[94] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[95] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[96] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[97] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[98] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[99] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind71(x, y);
 input [36:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[101] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[102] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[103] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[104] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[105] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[106] = t[127] ^ x[7];
  assign t[107] = t[128] ^ x[34];
  assign t[108] = t[129] ^ x[32];
  assign t[109] = t[130] ^ x[35];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[8];
  assign t[111] = t[132] ^ x[36];
  assign t[112] = t[133] ^ x[6];
  assign t[113] = t[134] ^ x[14];
  assign t[114] = t[135] ^ x[16];
  assign t[115] = t[136] ^ x[15];
  assign t[116] = t[137] ^ x[17];
  assign t[117] = t[138] ^ x[18];
  assign t[118] = t[139] ^ x[19];
  assign t[119] = t[140] ^ x[13];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[25];
  assign t[121] = t[142] ^ x[27];
  assign t[122] = t[143] ^ x[26];
  assign t[123] = t[144] ^ x[28];
  assign t[124] = t[145] ^ x[29];
  assign t[125] = t[146] ^ x[30];
  assign t[126] = t[147] ^ x[24];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[135] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[136] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[137] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[138] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[139] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[141] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[142] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[143] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[144] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[145] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[146] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[147] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[61]);
  assign t[15] = ~(t[60] ^ t[14]);
  assign t[16] = t[62] ^ t[61];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[60] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[60] ^ t[27];
  assign t[23] = t[63] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[61] ^ t[64];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[65]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[63] ^ t[29]);
  assign t[31] = t[66] ^ t[65];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[63] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[63] ^ t[36];
  assign t[36] = t[65] ^ t[67];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[68]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[60] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[59]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[63] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[42]);
  assign t[56] = ~(t[57] ^ t[69]);
  assign t[57] = ~t[58];
  assign t[58] = ~(t[48]);
  assign t[59] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[61] = (t[72] & ~t[75] & ~t[77]) | (~t[74] & t[75] & ~t[76]) | (~t[72] & ~t[75] & t[77]) | (t[74] & t[75] & t[76]);
  assign t[62] = (t[72] & ~t[76]) | (~t[72] & t[76]);
  assign t[63] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[64] = (t[72] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[77]) | (~t[72] & ~t[75] & t[76]) | (t[74] & t[75] & t[77]);
  assign t[65] = (t[78] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[78] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[66] = (t[78] & ~t[82]) | (~t[78] & t[82]);
  assign t[67] = (t[78] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[78] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[68] = (t[70] & ~t[84]) | (~t[70] & t[84]);
  assign t[69] = (t[70] & ~t[86] & ~t[71]) | (~t[85] & t[86] & ~t[87]) | (~t[70] & ~t[86] & t[71]) | (t[85] & t[86] & t[87]);
  assign t[6] = t[10] & t[11];
  assign t[70] = t[88] ^ x[7];
  assign t[71] = t[89] ^ x[8];
  assign t[72] = t[90] ^ x[14];
  assign t[73] = t[91] ^ x[15];
  assign t[74] = t[92] ^ x[16];
  assign t[75] = t[93] ^ x[17];
  assign t[76] = t[94] ^ x[18];
  assign t[77] = t[95] ^ x[19];
  assign t[78] = t[96] ^ x[25];
  assign t[79] = t[97] ^ x[26];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[27];
  assign t[81] = t[99] ^ x[28];
  assign t[82] = t[100] ^ x[29];
  assign t[83] = t[101] ^ x[30];
  assign t[84] = t[102] ^ x[32];
  assign t[85] = t[103] ^ x[34];
  assign t[86] = t[104] ^ x[35];
  assign t[87] = t[105] ^ x[36];
  assign t[88] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[89] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[8] = t[60] & t[13];
  assign t[90] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[93] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[96] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[97] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[98] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[99] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind72(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[19];
  assign t[102] = t[123] ^ x[20];
  assign t[103] = t[124] ^ x[14];
  assign t[104] = t[125] ^ x[26];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[27];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[30];
  assign t[109] = t[130] ^ x[31];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[25];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[119] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[121] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[122] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[123] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[124] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[125] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[126] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[127] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[128] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[129] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[131] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[48]);
  assign t[15] = ~(t[47] ^ t[14]);
  assign t[16] = t[49] ^ t[48];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[47] ^ t[27];
  assign t[23] = t[50] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[48] ^ t[51];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[52]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[50] ^ t[29]);
  assign t[31] = t[53] ^ t[52];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[50] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[50] ^ t[36];
  assign t[36] = t[52] ^ t[54];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[27] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[36] ^ t[24];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[58] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[49] = (t[58] & ~t[62]) | (~t[58] & t[62]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[58] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[52] = (t[64] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[64] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[64] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[57]) | (~t[56] & ~t[71] & t[72]) | (t[70] & t[71] & t[57]);
  assign t[56] = t[73] ^ x[8];
  assign t[57] = t[74] ^ x[9];
  assign t[58] = t[75] ^ x[15];
  assign t[59] = t[76] ^ x[16];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[17];
  assign t[61] = t[78] ^ x[18];
  assign t[62] = t[79] ^ x[19];
  assign t[63] = t[80] ^ x[20];
  assign t[64] = t[81] ^ x[26];
  assign t[65] = t[82] ^ x[27];
  assign t[66] = t[83] ^ x[28];
  assign t[67] = t[84] ^ x[29];
  assign t[68] = t[85] ^ x[30];
  assign t[69] = t[86] ^ x[31];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[33];
  assign t[71] = t[88] ^ x[34];
  assign t[72] = t[89] ^ x[35];
  assign t[73] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[86] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[87] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[88] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[47] & t[13];
  assign t[90] = t[111] ^ x[8];
  assign t[91] = t[112] ^ x[33];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[9];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[15];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[16];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind73(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[20];
  assign t[105] = t[126] ^ x[14];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[31];
  assign t[112] = t[133] ^ x[25];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[121] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[122] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[123] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[126] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[127] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[128] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[129] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[132] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[133] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[50]);
  assign t[15] = ~(t[49] ^ t[14]);
  assign t[16] = t[51] ^ t[50];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[49] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[49] ^ t[27];
  assign t[23] = t[52] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[50] ^ t[53];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[54]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[52] ^ t[29]);
  assign t[31] = t[55] ^ t[54];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[52] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[52] ^ t[36];
  assign t[36] = t[54] ^ t[56];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[57]);
  assign t[42] = t[44] ^ t[9];
  assign t[43] = ~t[45];
  assign t[44] = t[16] ^ t[21];
  assign t[45] = ~(t[46]);
  assign t[46] = t[47] ^ t[24];
  assign t[47] = t[31] ^ t[34];
  assign t[48] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[49] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[60] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[60] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[51] = (t[60] & ~t[64]) | (~t[60] & t[64]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[60] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[60] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[54] = (t[66] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[66] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[55] = (t[66] & ~t[70]) | (~t[66] & t[70]);
  assign t[56] = (t[66] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[66] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[57] = (t[58] & ~t[73] & ~t[59]) | (~t[72] & t[73] & ~t[74]) | (~t[58] & ~t[73] & t[59]) | (t[72] & t[73] & t[74]);
  assign t[58] = t[75] ^ x[8];
  assign t[59] = t[76] ^ x[9];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[15];
  assign t[61] = t[78] ^ x[16];
  assign t[62] = t[79] ^ x[17];
  assign t[63] = t[80] ^ x[18];
  assign t[64] = t[81] ^ x[19];
  assign t[65] = t[82] ^ x[20];
  assign t[66] = t[83] ^ x[26];
  assign t[67] = t[84] ^ x[27];
  assign t[68] = t[85] ^ x[28];
  assign t[69] = t[86] ^ x[29];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[30];
  assign t[71] = t[88] ^ x[31];
  assign t[72] = t[89] ^ x[33];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[35];
  assign t[75] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[76] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[77] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[8] = t[49] & t[13];
  assign t[90] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[7];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind74(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[15];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[16];
  assign t[104] = t[125] ^ x[19];
  assign t[105] = t[126] ^ x[13];
  assign t[106] = t[127] ^ x[25];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[26];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[27];
  assign t[111] = t[132] ^ x[30];
  assign t[112] = t[133] ^ x[24];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[47] ^ t[15];
  assign t[120] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[121] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[122] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[123] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[124] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[125] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[126] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[127] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[128] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[129] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[131] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[132] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[133] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[48] ^ t[49];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[49]);
  assign t[16] = ~(t[47] ^ t[15]);
  assign t[17] = t[47] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[50] ^ t[30];
  assign t[26] = t[49] ^ t[51];
  assign t[27] = t[47] ^ t[13];
  assign t[28] = t[52] ^ t[53];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[50] ^ t[30]);
  assign t[32] = t[50] & t[34];
  assign t[33] = t[50] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[53] ^ t[54];
  assign t[36] = t[50] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[26] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[35] ^ t[23];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[60]) | (~t[58] & t[60]);
  assign t[49] = (t[58] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[60]) | (~t[58] & ~t[62] & t[63]) | (t[61] & t[62] & t[60]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[62] & ~t[60]) | (~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[62] & t[60]) | (t[61] & t[62] & t[63]);
  assign t[52] = (t[64] & ~t[66]) | (~t[64] & t[66]);
  assign t[53] = (t[64] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[66]) | (~t[64] & ~t[68] & t[69]) | (t[67] & t[68] & t[66]);
  assign t[54] = (t[64] & ~t[68] & ~t[66]) | (~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[68] & t[66]) | (t[67] & t[68] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[56] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = t[74] ^ x[7];
  assign t[57] = t[75] ^ x[8];
  assign t[58] = t[76] ^ x[14];
  assign t[59] = t[77] ^ x[15];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[16];
  assign t[61] = t[79] ^ x[17];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[19];
  assign t[64] = t[82] ^ x[25];
  assign t[65] = t[83] ^ x[26];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[29];
  assign t[69] = t[87] ^ x[30];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[32];
  assign t[71] = t[89] ^ x[33];
  assign t[72] = t[90] ^ x[34];
  assign t[73] = t[91] ^ x[35];
  assign t[74] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[83] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[89] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[7];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[8];
  assign t[95] = t[116] ^ x[33];
  assign t[96] = t[117] ^ x[34];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[6];
  assign t[99] = t[120] ^ x[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind75(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[19];
  assign t[103] = t[124] ^ x[13];
  assign t[104] = t[125] ^ x[25];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[30];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[24];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[119] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[11] = t[45] ^ t[15];
  assign t[120] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[121] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[122] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[123] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[126] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[127] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[128] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[129] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[46] ^ t[47];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[47]);
  assign t[16] = ~(t[45] ^ t[15]);
  assign t[17] = t[45] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[45] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[48] ^ t[30];
  assign t[26] = t[47] ^ t[49];
  assign t[27] = t[45] ^ t[13];
  assign t[28] = t[50] ^ t[51];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[51]);
  assign t[31] = ~(t[48] ^ t[30]);
  assign t[32] = t[48] & t[34];
  assign t[33] = t[48] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[51] ^ t[52];
  assign t[36] = t[48] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[5]);
  assign t[41] = ~(t[42] ^ t[53]);
  assign t[42] = ~t[43];
  assign t[43] = ~(t[18]);
  assign t[44] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[56] & ~t[58]) | (~t[56] & t[58]);
  assign t[47] = (t[56] & ~t[60] & ~t[61]) | (~t[59] & t[60] & ~t[58]) | (~t[56] & ~t[60] & t[61]) | (t[59] & t[60] & t[58]);
  assign t[48] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[49] = (t[56] & ~t[60] & ~t[58]) | (~t[59] & t[60] & ~t[61]) | (~t[56] & ~t[60] & t[58]) | (t[59] & t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[44]);
  assign t[50] = (t[62] & ~t[64]) | (~t[62] & t[64]);
  assign t[51] = (t[62] & ~t[66] & ~t[67]) | (~t[65] & t[66] & ~t[64]) | (~t[62] & ~t[66] & t[67]) | (t[65] & t[66] & t[64]);
  assign t[52] = (t[62] & ~t[66] & ~t[64]) | (~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[66] & t[64]) | (t[65] & t[66] & t[67]);
  assign t[53] = (t[54] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[54] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[54] = t[72] ^ x[7];
  assign t[55] = t[73] ^ x[8];
  assign t[56] = t[74] ^ x[14];
  assign t[57] = t[75] ^ x[15];
  assign t[58] = t[76] ^ x[16];
  assign t[59] = t[77] ^ x[17];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[25];
  assign t[63] = t[81] ^ x[26];
  assign t[64] = t[82] ^ x[27];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[29];
  assign t[67] = t[85] ^ x[30];
  assign t[68] = t[86] ^ x[32];
  assign t[69] = t[87] ^ x[33];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[34];
  assign t[71] = t[89] ^ x[35];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[81] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[86] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[87] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[88] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[111] ^ x[7];
  assign t[91] = t[112] ^ x[32];
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[6];
  assign t[97] = t[118] ^ x[14];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind76(x, y);
 input [35:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[101] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[102] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[103] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[104] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[105] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[35]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[114] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[115] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[116] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[118] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[119] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[11] = ~(t[37] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[38] ^ t[39];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = x[0] ? x[35] : t[18];
  assign t[18] = ~(t[19] ^ t[20]);
  assign t[19] = ~t[21];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[23] ^ t[41]);
  assign t[22] = t[24] ^ t[8];
  assign t[23] = ~t[25];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = ~(t[28]);
  assign t[26] = t[42] ^ t[35];
  assign t[27] = t[10] & t[29];
  assign t[28] = t[30] ^ t[14];
  assign t[29] = t[37] ^ t[7];
  assign t[2] = ~t[4];
  assign t[30] = t[31] ^ t[32];
  assign t[31] = t[43] ^ t[38];
  assign t[32] = t[15] & t[33];
  assign t[33] = t[40] ^ t[13];
  assign t[34] = (t[44] & ~t[46] & ~t[48]) | (~t[45] & t[46] & ~t[47]) | (~t[44] & ~t[46] & t[48]) | (t[45] & t[46] & t[47]);
  assign t[35] = (t[49] & ~t[51] & ~t[53]) | (~t[50] & t[51] & ~t[52]) | (~t[49] & ~t[51] & t[53]) | (t[50] & t[51] & t[52]);
  assign t[36] = (t[49] & ~t[51] & ~t[52]) | (~t[50] & t[51] & ~t[53]) | (~t[49] & ~t[51] & t[52]) | (t[50] & t[51] & t[53]);
  assign t[37] = (t[49] & ~t[54]) | (~t[49] & t[54]);
  assign t[38] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[39] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[60]) | (~t[55] & t[60]);
  assign t[41] = (t[44] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[44] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[42] = (t[49] & ~t[52]) | (~t[49] & t[52]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = t[61] ^ x[8];
  assign t[45] = t[62] ^ x[9];
  assign t[46] = t[63] ^ x[10];
  assign t[47] = t[64] ^ x[11];
  assign t[48] = t[65] ^ x[12];
  assign t[49] = t[66] ^ x[18];
  assign t[4] = ~(t[6] ^ t[34]);
  assign t[50] = t[67] ^ x[19];
  assign t[51] = t[68] ^ x[20];
  assign t[52] = t[69] ^ x[21];
  assign t[53] = t[70] ^ x[22];
  assign t[54] = t[71] ^ x[23];
  assign t[55] = t[72] ^ x[29];
  assign t[56] = t[73] ^ x[30];
  assign t[57] = t[74] ^ x[31];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[34];
  assign t[61] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[62] = (t[79] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (~t[78] & t[79] & ~t[81] & ~t[82] & ~t[84]) | (~t[78] & t[79] & ~t[80] & ~t[83] & ~t[84]) | (t[78] & ~t[79] & t[80] & t[81] & ~t[84]) | (t[78] & ~t[79] & t[82] & t[83] & ~t[84]) | (t[79] & ~t[81] & ~t[83] & t[84]) | (~t[79] & t[81] & t[83] & t[84]);
  assign t[63] = (t[78] & t[79] & t[80] & ~t[81] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & ~t[81] & ~t[82] & t[83] & t[84]) | (~t[79] & ~t[80] & t[81] & ~t[82] & ~t[83]) | (~t[78] & ~t[80] & t[81] & ~t[83] & ~t[84]) | (~t[78] & ~t[79] & t[81] & ~t[82] & ~t[84]) | (~t[79] & t[80] & t[81] & t[82] & ~t[83]) | (~t[80] & t[81] & t[82] & ~t[84]);
  assign t[64] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[65] = (t[78] & t[79] & ~t[81] & t[82] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & ~t[81] & ~t[82] & t[83]) | (~t[78] & ~t[81] & ~t[82] & t[83] & ~t[84]) | (~t[78] & ~t[79] & ~t[80] & t[83] & ~t[84]) | (~t[79] & t[80] & ~t[81] & t[82] & t[83]) | (t[80] & ~t[82] & t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = ~t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[72] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[73] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[74] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[8];
  assign t[79] = t[100] ^ x[9];
  assign t[7] = t[35] ^ t[36];
  assign t[80] = t[101] ^ x[6];
  assign t[81] = t[102] ^ x[10];
  assign t[82] = t[103] ^ x[11];
  assign t[83] = t[104] ^ x[12];
  assign t[84] = t[105] ^ x[7];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[23];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[29];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[32];
  assign t[97] = t[118] ^ x[33];
  assign t[98] = t[119] ^ x[28];
  assign t[99] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~t[17]) | (~t[0] & t[17]);
endmodule

module R2ind77(x, y);
 input [60:0] x;
 output y;

 wire [212:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[50];
  assign t[101] = t[125] ^ x[51];
  assign t[102] = t[126] ^ x[52];
  assign t[103] = t[127] ^ x[59];
  assign t[104] = t[128] ^ x[60];
  assign t[105] = (t[129] & ~t[131] & ~t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[132] & ~t[133] & ~t[135]) | (t[129] & ~t[130] & ~t[131] & ~t[134] & ~t[135]) | (~t[129] & t[130] & t[131] & t[132] & ~t[135]) | (~t[129] & t[130] & t[133] & t[134] & ~t[135]) | (t[129] & ~t[131] & ~t[133] & t[135]) | (~t[129] & t[131] & t[133] & t[135]);
  assign t[106] = (t[129] & t[130] & ~t[131] & ~t[133] & t[134] & ~t[135]) | (t[129] & t[131] & ~t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[131] & t[133] & ~t[134] & ~t[135]) | (~t[129] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[129] & ~t[130] & ~t[132] & t[133] & ~t[135]) | (~t[129] & ~t[131] & t[132] & t[133] & t[134]) | (t[132] & t[133] & ~t[134] & ~t[135]);
  assign t[107] = (t[136] & ~t[138] & ~t[139] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & ~t[139] & ~t[140] & ~t[142]) | (t[136] & ~t[137] & ~t[138] & ~t[141] & ~t[142]) | (~t[136] & t[137] & t[138] & t[139] & ~t[142]) | (~t[136] & t[137] & t[140] & t[141] & ~t[142]) | (t[136] & ~t[138] & ~t[140] & t[142]) | (~t[136] & t[138] & t[140] & t[142]);
  assign t[108] = (t[136] & t[137] & ~t[138] & t[139] & ~t[140] & ~t[142]) | (t[136] & ~t[138] & ~t[139] & t[140] & ~t[141] & t[142]) | (~t[137] & t[138] & ~t[139] & ~t[140] & ~t[142]) | (~t[136] & t[138] & ~t[139] & ~t[140] & ~t[141]) | (~t[136] & ~t[137] & t[138] & ~t[141] & ~t[142]) | (~t[136] & t[138] & t[139] & ~t[140] & t[141]) | (t[138] & ~t[139] & t[141] & ~t[142]);
  assign t[109] = (t[143] & ~t[145] & ~t[146] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & ~t[146] & ~t[147] & ~t[149]) | (t[143] & ~t[144] & ~t[145] & ~t[148] & ~t[149]) | (~t[143] & t[144] & t[145] & t[146] & ~t[149]) | (~t[143] & t[144] & t[147] & t[148] & ~t[149]) | (t[143] & ~t[145] & ~t[147] & t[149]) | (~t[143] & t[145] & t[147] & t[149]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (t[143] & t[144] & ~t[145] & ~t[147] & t[148] & ~t[149]) | (t[143] & t[145] & ~t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[145] & t[147] & ~t[148] & ~t[149]) | (~t[143] & ~t[145] & ~t[146] & t[147] & ~t[148]) | (~t[143] & ~t[144] & ~t[146] & t[147] & ~t[149]) | (~t[143] & ~t[145] & t[146] & t[147] & t[148]) | (t[146] & t[147] & ~t[148] & ~t[149]);
  assign t[111] = (t[137] & ~t[138] & ~t[139] & ~t[140] & ~t[141]) | (~t[136] & t[137] & ~t[139] & ~t[140] & ~t[142]) | (~t[136] & t[137] & ~t[138] & ~t[141] & ~t[142]) | (t[136] & ~t[137] & t[138] & t[139] & ~t[142]) | (t[136] & ~t[137] & t[140] & t[141] & ~t[142]) | (t[137] & ~t[139] & ~t[141] & t[142]) | (~t[137] & t[139] & t[141] & t[142]);
  assign t[112] = (t[136] & t[137] & t[138] & ~t[139] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & ~t[139] & ~t[140] & t[141] & t[142]) | (~t[137] & ~t[138] & t[139] & ~t[140] & ~t[141]) | (~t[136] & ~t[138] & t[139] & ~t[141] & ~t[142]) | (~t[136] & ~t[137] & t[139] & ~t[140] & ~t[142]) | (~t[137] & t[138] & t[139] & t[140] & ~t[141]) | (~t[138] & t[139] & t[140] & ~t[142]);
  assign t[113] = (t[136] & t[137] & ~t[138] & ~t[140] & t[141] & ~t[142]) | (t[136] & t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[142]) | (~t[136] & ~t[138] & ~t[139] & t[140] & ~t[141]) | (~t[136] & ~t[137] & ~t[139] & t[140] & ~t[142]) | (~t[136] & ~t[138] & t[139] & t[140] & t[141]) | (t[139] & t[140] & ~t[141] & ~t[142]);
  assign t[114] = (t[136] & t[137] & ~t[139] & t[140] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[138] & ~t[139] & ~t[140] & t[141]) | (~t[136] & ~t[139] & ~t[140] & t[141] & ~t[142]) | (~t[136] & ~t[137] & ~t[138] & t[141] & ~t[142]) | (~t[137] & t[138] & ~t[139] & t[140] & t[141]) | (t[138] & ~t[140] & t[141] & ~t[142]);
  assign t[115] = (t[150] & ~t[152] & ~t[153] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & ~t[153] & ~t[154] & ~t[156]) | (t[150] & ~t[151] & ~t[152] & ~t[155] & ~t[156]) | (~t[150] & t[151] & t[152] & t[153] & ~t[156]) | (~t[150] & t[151] & t[154] & t[155] & ~t[156]) | (t[150] & ~t[152] & ~t[154] & t[156]) | (~t[150] & t[152] & t[154] & t[156]);
  assign t[116] = (t[150] & t[151] & ~t[152] & t[153] & ~t[154] & ~t[156]) | (t[150] & ~t[152] & ~t[153] & t[154] & ~t[155] & t[156]) | (~t[151] & t[152] & ~t[153] & ~t[154] & ~t[156]) | (~t[150] & t[152] & ~t[153] & ~t[154] & ~t[155]) | (~t[150] & ~t[151] & t[152] & ~t[155] & ~t[156]) | (~t[150] & t[152] & t[153] & ~t[154] & t[155]) | (t[152] & ~t[153] & t[155] & ~t[156]);
  assign t[117] = (t[151] & ~t[152] & ~t[153] & ~t[154] & ~t[155]) | (~t[150] & t[151] & ~t[153] & ~t[154] & ~t[156]) | (~t[150] & t[151] & ~t[152] & ~t[155] & ~t[156]) | (t[150] & ~t[151] & t[152] & t[153] & ~t[156]) | (t[150] & ~t[151] & t[154] & t[155] & ~t[156]) | (t[151] & ~t[153] & ~t[155] & t[156]) | (~t[151] & t[153] & t[155] & t[156]);
  assign t[118] = (t[150] & t[151] & t[152] & ~t[153] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & ~t[153] & ~t[154] & t[155] & t[156]) | (~t[151] & ~t[152] & t[153] & ~t[154] & ~t[155]) | (~t[150] & ~t[152] & t[153] & ~t[155] & ~t[156]) | (~t[150] & ~t[151] & t[153] & ~t[154] & ~t[156]) | (~t[151] & t[152] & t[153] & t[154] & ~t[155]) | (~t[152] & t[153] & t[154] & ~t[156]);
  assign t[119] = (t[150] & t[151] & ~t[152] & ~t[154] & t[155] & ~t[156]) | (t[150] & t[152] & ~t[153] & ~t[154] & ~t[155] & t[156]) | (~t[151] & ~t[152] & t[154] & ~t[155] & ~t[156]) | (~t[150] & ~t[152] & ~t[153] & t[154] & ~t[155]) | (~t[150] & ~t[151] & ~t[153] & t[154] & ~t[156]) | (~t[150] & ~t[152] & t[153] & t[154] & t[155]) | (t[153] & t[154] & ~t[155] & ~t[156]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (t[150] & t[151] & ~t[153] & t[154] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & t[153] & ~t[154] & ~t[155] & t[156]) | (~t[151] & ~t[152] & ~t[153] & ~t[154] & t[155]) | (~t[150] & ~t[153] & ~t[154] & t[155] & ~t[156]) | (~t[150] & ~t[151] & ~t[152] & t[155] & ~t[156]) | (~t[151] & t[152] & ~t[153] & t[154] & t[155]) | (t[152] & ~t[154] & t[155] & ~t[156]);
  assign t[121] = (t[129] & t[130] & ~t[131] & t[132] & ~t[133] & ~t[135]) | (t[129] & ~t[131] & ~t[132] & t[133] & ~t[134] & t[135]) | (~t[130] & t[131] & ~t[132] & ~t[133] & ~t[135]) | (~t[129] & t[131] & ~t[132] & ~t[133] & ~t[134]) | (~t[129] & ~t[130] & t[131] & ~t[134] & ~t[135]) | (~t[129] & t[131] & t[132] & ~t[133] & t[134]) | (t[131] & ~t[132] & t[134] & ~t[135]);
  assign t[122] = (t[157] & ~t[159] & ~t[160] & ~t[161] & ~t[162]) | (t[157] & ~t[158] & ~t[160] & ~t[161] & ~t[163]) | (t[157] & ~t[158] & ~t[159] & ~t[162] & ~t[163]) | (~t[157] & t[158] & t[159] & t[160] & ~t[163]) | (~t[157] & t[158] & t[161] & t[162] & ~t[163]) | (t[157] & ~t[159] & ~t[161] & t[163]) | (~t[157] & t[159] & t[161] & t[163]);
  assign t[123] = (t[157] & t[158] & ~t[159] & ~t[161] & t[162] & ~t[163]) | (t[157] & t[159] & ~t[160] & ~t[161] & ~t[162] & t[163]) | (~t[158] & ~t[159] & t[161] & ~t[162] & ~t[163]) | (~t[157] & ~t[159] & ~t[160] & t[161] & ~t[162]) | (~t[157] & ~t[158] & ~t[160] & t[161] & ~t[163]) | (~t[157] & ~t[159] & t[160] & t[161] & t[162]) | (t[160] & t[161] & ~t[162] & ~t[163]);
  assign t[124] = (t[130] & ~t[131] & ~t[132] & ~t[133] & ~t[134]) | (~t[129] & t[130] & ~t[132] & ~t[133] & ~t[135]) | (~t[129] & t[130] & ~t[131] & ~t[134] & ~t[135]) | (t[129] & ~t[130] & t[131] & t[132] & ~t[135]) | (t[129] & ~t[130] & t[133] & t[134] & ~t[135]) | (t[130] & ~t[132] & ~t[134] & t[135]) | (~t[130] & t[132] & t[134] & t[135]);
  assign t[125] = (t[129] & t[130] & t[131] & ~t[132] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[132] & ~t[133] & t[134] & t[135]) | (~t[130] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (~t[129] & ~t[131] & t[132] & ~t[134] & ~t[135]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[135]) | (~t[130] & t[131] & t[132] & t[133] & ~t[134]) | (~t[131] & t[132] & t[133] & ~t[135]);
  assign t[126] = (t[129] & t[130] & ~t[132] & t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[129] & ~t[130] & ~t[131] & t[134] & ~t[135]) | (~t[130] & t[131] & ~t[132] & t[133] & t[134]) | (t[131] & ~t[133] & t[134] & ~t[135]);
  assign t[127] = (t[164] & ~t[166] & ~t[167] & ~t[168] & ~t[169]) | (t[164] & ~t[165] & ~t[167] & ~t[168] & ~t[170]) | (t[164] & ~t[165] & ~t[166] & ~t[169] & ~t[170]) | (~t[164] & t[165] & t[166] & t[167] & ~t[170]) | (~t[164] & t[165] & t[168] & t[169] & ~t[170]) | (t[164] & ~t[166] & ~t[168] & t[170]) | (~t[164] & t[166] & t[168] & t[170]);
  assign t[128] = (t[164] & t[165] & ~t[166] & ~t[168] & t[169] & ~t[170]) | (t[164] & t[166] & ~t[167] & ~t[168] & ~t[169] & t[170]) | (~t[165] & ~t[166] & t[168] & ~t[169] & ~t[170]) | (~t[164] & ~t[166] & ~t[167] & t[168] & ~t[169]) | (~t[164] & ~t[165] & ~t[167] & t[168] & ~t[170]) | (~t[164] & ~t[166] & t[167] & t[168] & t[169]) | (t[167] & t[168] & ~t[169] & ~t[170]);
  assign t[129] = t[171] ^ x[7];
  assign t[12] = ~(t[18] ^ t[69]);
  assign t[130] = t[172] ^ x[50];
  assign t[131] = t[173] ^ x[40];
  assign t[132] = t[174] ^ x[51];
  assign t[133] = t[175] ^ x[8];
  assign t[134] = t[176] ^ x[52];
  assign t[135] = t[177] ^ x[6];
  assign t[136] = t[178] ^ x[14];
  assign t[137] = t[179] ^ x[24];
  assign t[138] = t[180] ^ x[15];
  assign t[139] = t[181] ^ x[25];
  assign t[13] = t[19] ^ t[20];
  assign t[140] = t[182] ^ x[26];
  assign t[141] = t[183] ^ x[27];
  assign t[142] = t[184] ^ x[13];
  assign t[143] = t[185] ^ x[22];
  assign t[144] = t[186] ^ x[17];
  assign t[145] = t[187] ^ x[18];
  assign t[146] = t[188] ^ x[19];
  assign t[147] = t[189] ^ x[23];
  assign t[148] = t[190] ^ x[20];
  assign t[149] = t[191] ^ x[21];
  assign t[14] = ~(t[70]);
  assign t[150] = t[192] ^ x[33];
  assign t[151] = t[193] ^ x[35];
  assign t[152] = t[194] ^ x[34];
  assign t[153] = t[195] ^ x[36];
  assign t[154] = t[196] ^ x[37];
  assign t[155] = t[197] ^ x[38];
  assign t[156] = t[198] ^ x[32];
  assign t[157] = t[199] ^ x[47];
  assign t[158] = t[200] ^ x[42];
  assign t[159] = t[201] ^ x[43];
  assign t[15] = ~(t[68] ^ t[14]);
  assign t[160] = t[202] ^ x[44];
  assign t[161] = t[203] ^ x[48];
  assign t[162] = t[204] ^ x[45];
  assign t[163] = t[205] ^ x[46];
  assign t[164] = t[206] ^ x[59];
  assign t[165] = t[207] ^ x[54];
  assign t[166] = t[208] ^ x[55];
  assign t[167] = t[209] ^ x[56];
  assign t[168] = t[210] ^ x[60];
  assign t[169] = t[211] ^ x[57];
  assign t[16] = t[71] ^ t[70];
  assign t[170] = t[212] ^ x[58];
  assign t[171] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[172] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[173] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[174] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[175] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[176] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[177] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[178] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[179] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[180] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[181] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[182] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[183] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[184] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[185] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[186] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[187] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[188] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[189] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = ~t[22];
  assign t[190] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[192] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[193] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[194] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[195] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[196] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[197] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[198] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[199] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[19] = t[68] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[201] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[202] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[203] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[204] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[205] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[206] = (x[53] & ~1'b0 & ~1'b0) | (~x[53] & 1'b0 & ~1'b0) | (~x[53] & ~1'b0 & 1'b0) | (x[53] & 1'b0 & 1'b0);
  assign t[207] = (x[53] & ~1'b0 & ~1'b0) | (~x[53] & 1'b0 & ~1'b0) | (~x[53] & ~1'b0 & 1'b0) | (x[53] & 1'b0 & 1'b0);
  assign t[208] = (x[53] & ~1'b0) | (~x[53] & 1'b0);
  assign t[209] = (x[53] & ~1'b0) | (~x[53] & 1'b0);
  assign t[20] = t[14] & t[21];
  assign t[210] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[211] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[212] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[21] = t[68] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[70] ^ t[72];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[73] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[74]);
  assign t[32] = ~(t[73] ^ t[31]);
  assign t[33] = t[75] ^ t[74];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[73] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[73] ^ t[38];
  assign t[38] = t[74] ^ t[76];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~(t[46] ^ t[77]);
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~t[49];
  assign t[47] = t[16] ^ t[20];
  assign t[48] = t[68] ^ t[14];
  assign t[49] = ~(t[50] ^ t[78]);
  assign t[4] = ~(t[7] ^ t[67]);
  assign t[50] = ~t[51];
  assign t[51] = ~(t[52] ^ t[53]);
  assign t[52] = t[54] ^ t[27];
  assign t[53] = t[24] ^ t[55];
  assign t[54] = t[33] ^ t[36];
  assign t[55] = t[73] ^ t[31];
  assign t[56] = x[0] ? x[49] : t[57];
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = ~(t[61]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[62] ^ t[79]);
  assign t[61] = t[23] ^ t[9];
  assign t[62] = ~t[63];
  assign t[63] = ~(t[64] ^ t[80]);
  assign t[64] = ~t[65];
  assign t[65] = ~(t[66]);
  assign t[66] = t[38] ^ t[27];
  assign t[67] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[68] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[69] = (t[85] & ~t[86]) | (~t[85] & t[86]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[83] & ~t[88] & ~t[90]) | (~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[88] & t[90]) | (t[87] & t[88] & t[89]);
  assign t[71] = (t[83] & ~t[89]) | (~t[83] & t[89]);
  assign t[72] = (t[83] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[90]) | (~t[83] & ~t[88] & t[89]) | (t[87] & t[88] & t[90]);
  assign t[73] = (t[91] & ~t[92]) | (~t[91] & t[92]);
  assign t[74] = (t[91] & ~t[94] & ~t[96]) | (~t[93] & t[94] & ~t[95]) | (~t[91] & ~t[94] & t[96]) | (t[93] & t[94] & t[95]);
  assign t[75] = (t[91] & ~t[95]) | (~t[91] & t[95]);
  assign t[76] = (t[91] & ~t[94] & ~t[95]) | (~t[93] & t[94] & ~t[96]) | (~t[91] & ~t[94] & t[95]) | (t[93] & t[94] & t[96]);
  assign t[77] = (t[81] & ~t[97]) | (~t[81] & t[97]);
  assign t[78] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[79] = (t[81] & ~t[101] & ~t[102]) | (~t[100] & t[101] & ~t[82]) | (~t[81] & ~t[101] & t[102]) | (t[100] & t[101] & t[82]);
  assign t[7] = ~t[12];
  assign t[80] = (t[103] & ~t[104]) | (~t[103] & t[104]);
  assign t[81] = t[105] ^ x[7];
  assign t[82] = t[106] ^ x[8];
  assign t[83] = t[107] ^ x[14];
  assign t[84] = t[108] ^ x[15];
  assign t[85] = t[109] ^ x[22];
  assign t[86] = t[110] ^ x[23];
  assign t[87] = t[111] ^ x[24];
  assign t[88] = t[112] ^ x[25];
  assign t[89] = t[113] ^ x[26];
  assign t[8] = t[68] & t[13];
  assign t[90] = t[114] ^ x[27];
  assign t[91] = t[115] ^ x[33];
  assign t[92] = t[116] ^ x[34];
  assign t[93] = t[117] ^ x[35];
  assign t[94] = t[118] ^ x[36];
  assign t[95] = t[119] ^ x[37];
  assign t[96] = t[120] ^ x[38];
  assign t[97] = t[121] ^ x[40];
  assign t[98] = t[122] ^ x[47];
  assign t[99] = t[123] ^ x[48];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39] & ~t[56]) | (~t[0] & t[39] & ~t[56]) | (~t[0] & ~t[39] & t[56]) | (t[0] & t[39] & t[56]);
endmodule

module R2ind78(x, y);
 input [60:0] x;
 output y;

 wire [210:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[52];
  assign t[101] = t[125] ^ x[59];
  assign t[102] = t[126] ^ x[60];
  assign t[103] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[104] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[105] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[106] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[107] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[108] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[109] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[111] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[112] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[113] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[114] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[115] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[116] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[117] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[118] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[119] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[121] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[122] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[123] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[124] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[125] = (t[162] & ~t[164] & ~t[165] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & ~t[165] & ~t[166] & ~t[168]) | (t[162] & ~t[163] & ~t[164] & ~t[167] & ~t[168]) | (~t[162] & t[163] & t[164] & t[165] & ~t[168]) | (~t[162] & t[163] & t[166] & t[167] & ~t[168]) | (t[162] & ~t[164] & ~t[166] & t[168]) | (~t[162] & t[164] & t[166] & t[168]);
  assign t[126] = (t[162] & t[163] & ~t[164] & ~t[166] & t[167] & ~t[168]) | (t[162] & t[164] & ~t[165] & ~t[166] & ~t[167] & t[168]) | (~t[163] & ~t[164] & t[166] & ~t[167] & ~t[168]) | (~t[162] & ~t[164] & ~t[165] & t[166] & ~t[167]) | (~t[162] & ~t[163] & ~t[165] & t[166] & ~t[168]) | (~t[162] & ~t[164] & t[165] & t[166] & t[167]) | (t[165] & t[166] & ~t[167] & ~t[168]);
  assign t[127] = t[169] ^ x[7];
  assign t[128] = t[170] ^ x[50];
  assign t[129] = t[171] ^ x[40];
  assign t[12] = ~(t[18] ^ t[67]);
  assign t[130] = t[172] ^ x[51];
  assign t[131] = t[173] ^ x[8];
  assign t[132] = t[174] ^ x[52];
  assign t[133] = t[175] ^ x[6];
  assign t[134] = t[176] ^ x[14];
  assign t[135] = t[177] ^ x[24];
  assign t[136] = t[178] ^ x[15];
  assign t[137] = t[179] ^ x[25];
  assign t[138] = t[180] ^ x[26];
  assign t[139] = t[181] ^ x[27];
  assign t[13] = t[19] ^ t[20];
  assign t[140] = t[182] ^ x[13];
  assign t[141] = t[183] ^ x[22];
  assign t[142] = t[184] ^ x[17];
  assign t[143] = t[185] ^ x[18];
  assign t[144] = t[186] ^ x[19];
  assign t[145] = t[187] ^ x[23];
  assign t[146] = t[188] ^ x[20];
  assign t[147] = t[189] ^ x[21];
  assign t[148] = t[190] ^ x[33];
  assign t[149] = t[191] ^ x[35];
  assign t[14] = ~(t[68]);
  assign t[150] = t[192] ^ x[34];
  assign t[151] = t[193] ^ x[36];
  assign t[152] = t[194] ^ x[37];
  assign t[153] = t[195] ^ x[38];
  assign t[154] = t[196] ^ x[32];
  assign t[155] = t[197] ^ x[47];
  assign t[156] = t[198] ^ x[42];
  assign t[157] = t[199] ^ x[43];
  assign t[158] = t[200] ^ x[44];
  assign t[159] = t[201] ^ x[48];
  assign t[15] = ~(t[66] ^ t[14]);
  assign t[160] = t[202] ^ x[45];
  assign t[161] = t[203] ^ x[46];
  assign t[162] = t[204] ^ x[59];
  assign t[163] = t[205] ^ x[54];
  assign t[164] = t[206] ^ x[55];
  assign t[165] = t[207] ^ x[56];
  assign t[166] = t[208] ^ x[60];
  assign t[167] = t[209] ^ x[57];
  assign t[168] = t[210] ^ x[58];
  assign t[169] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[16] = t[69] ^ t[68];
  assign t[170] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[171] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[172] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[173] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[174] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[175] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[176] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[177] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[178] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[179] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[180] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[181] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[182] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[183] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[184] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[185] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[186] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[187] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[188] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[189] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = ~t[22];
  assign t[190] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[191] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[192] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[193] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[194] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[195] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[196] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[197] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[198] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[199] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[19] = t[66] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[201] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[202] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[203] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[204] = (x[53] & ~1'b0 & ~1'b0) | (~x[53] & 1'b0 & ~1'b0) | (~x[53] & ~1'b0 & 1'b0) | (x[53] & 1'b0 & 1'b0);
  assign t[205] = (x[53] & ~1'b0 & ~1'b0) | (~x[53] & 1'b0 & ~1'b0) | (~x[53] & ~1'b0 & 1'b0) | (x[53] & 1'b0 & 1'b0);
  assign t[206] = (x[53] & ~1'b0) | (~x[53] & 1'b0);
  assign t[207] = (x[53] & ~1'b0) | (~x[53] & 1'b0);
  assign t[208] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[209] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[20] = t[14] & t[21];
  assign t[210] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[21] = t[66] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[68] ^ t[70];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[71] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[72]);
  assign t[32] = ~(t[71] ^ t[31]);
  assign t[33] = t[73] ^ t[72];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[71] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[71] ^ t[38];
  assign t[38] = t[72] ^ t[74];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~(t[46] ^ t[75]);
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~t[49];
  assign t[47] = t[16] ^ t[20];
  assign t[48] = t[66] ^ t[14];
  assign t[49] = ~(t[50] ^ t[76]);
  assign t[4] = ~(t[7] ^ t[65]);
  assign t[50] = ~t[51];
  assign t[51] = ~(t[52] ^ t[53]);
  assign t[52] = t[54] ^ t[27];
  assign t[53] = t[24] ^ t[55];
  assign t[54] = t[33] ^ t[36];
  assign t[55] = t[71] ^ t[31];
  assign t[56] = x[0] ? x[49] : t[57];
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = ~(t[44]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[61] ^ t[77]);
  assign t[61] = ~t[62];
  assign t[62] = ~(t[63] ^ t[78]);
  assign t[63] = ~t[64];
  assign t[64] = ~(t[52]);
  assign t[65] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[66] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[67] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[68] = (t[81] & ~t[86] & ~t[88]) | (~t[85] & t[86] & ~t[87]) | (~t[81] & ~t[86] & t[88]) | (t[85] & t[86] & t[87]);
  assign t[69] = (t[81] & ~t[87]) | (~t[81] & t[87]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[81] & ~t[86] & ~t[87]) | (~t[85] & t[86] & ~t[88]) | (~t[81] & ~t[86] & t[87]) | (t[85] & t[86] & t[88]);
  assign t[71] = (t[89] & ~t[90]) | (~t[89] & t[90]);
  assign t[72] = (t[89] & ~t[92] & ~t[94]) | (~t[91] & t[92] & ~t[93]) | (~t[89] & ~t[92] & t[94]) | (t[91] & t[92] & t[93]);
  assign t[73] = (t[89] & ~t[93]) | (~t[89] & t[93]);
  assign t[74] = (t[89] & ~t[92] & ~t[93]) | (~t[91] & t[92] & ~t[94]) | (~t[89] & ~t[92] & t[93]) | (t[91] & t[92] & t[94]);
  assign t[75] = (t[79] & ~t[95]) | (~t[79] & t[95]);
  assign t[76] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[77] = (t[79] & ~t[99] & ~t[80]) | (~t[98] & t[99] & ~t[100]) | (~t[79] & ~t[99] & t[80]) | (t[98] & t[99] & t[100]);
  assign t[78] = (t[101] & ~t[102]) | (~t[101] & t[102]);
  assign t[79] = t[103] ^ x[7];
  assign t[7] = ~t[12];
  assign t[80] = t[104] ^ x[8];
  assign t[81] = t[105] ^ x[14];
  assign t[82] = t[106] ^ x[15];
  assign t[83] = t[107] ^ x[22];
  assign t[84] = t[108] ^ x[23];
  assign t[85] = t[109] ^ x[24];
  assign t[86] = t[110] ^ x[25];
  assign t[87] = t[111] ^ x[26];
  assign t[88] = t[112] ^ x[27];
  assign t[89] = t[113] ^ x[33];
  assign t[8] = t[66] & t[13];
  assign t[90] = t[114] ^ x[34];
  assign t[91] = t[115] ^ x[35];
  assign t[92] = t[116] ^ x[36];
  assign t[93] = t[117] ^ x[37];
  assign t[94] = t[118] ^ x[38];
  assign t[95] = t[119] ^ x[40];
  assign t[96] = t[120] ^ x[47];
  assign t[97] = t[121] ^ x[48];
  assign t[98] = t[122] ^ x[50];
  assign t[99] = t[123] ^ x[51];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39] & ~t[56]) | (~t[0] & t[39] & ~t[56]) | (~t[0] & ~t[39] & t[56]) | (t[0] & t[39] & t[56]);
endmodule

module R2ind79(x, y);
 input [51:0] x;
 output y;

 wire [173:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[101] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[102] = (t[132] & ~t[134] & ~t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[135] & ~t[136] & ~t[138]) | (t[132] & ~t[133] & ~t[134] & ~t[137] & ~t[138]) | (~t[132] & t[133] & t[134] & t[135] & ~t[138]) | (~t[132] & t[133] & t[136] & t[137] & ~t[138]) | (t[132] & ~t[134] & ~t[136] & t[138]) | (~t[132] & t[134] & t[136] & t[138]);
  assign t[103] = (t[132] & t[133] & ~t[134] & ~t[136] & t[137] & ~t[138]) | (t[132] & t[134] & ~t[135] & ~t[136] & ~t[137] & t[138]) | (~t[133] & ~t[134] & t[136] & ~t[137] & ~t[138]) | (~t[132] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[132] & ~t[133] & ~t[135] & t[136] & ~t[138]) | (~t[132] & ~t[134] & t[135] & t[136] & t[137]) | (t[135] & t[136] & ~t[137] & ~t[138]);
  assign t[104] = t[139] ^ x[8];
  assign t[105] = t[140] ^ x[41];
  assign t[106] = t[141] ^ x[6];
  assign t[107] = t[142] ^ x[42];
  assign t[108] = t[143] ^ x[9];
  assign t[109] = t[144] ^ x[43];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[145] ^ x[7];
  assign t[111] = t[146] ^ x[15];
  assign t[112] = t[147] ^ x[25];
  assign t[113] = t[148] ^ x[16];
  assign t[114] = t[149] ^ x[26];
  assign t[115] = t[150] ^ x[27];
  assign t[116] = t[151] ^ x[28];
  assign t[117] = t[152] ^ x[14];
  assign t[118] = t[153] ^ x[23];
  assign t[119] = t[154] ^ x[18];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[155] ^ x[19];
  assign t[121] = t[156] ^ x[20];
  assign t[122] = t[157] ^ x[24];
  assign t[123] = t[158] ^ x[21];
  assign t[124] = t[159] ^ x[22];
  assign t[125] = t[160] ^ x[34];
  assign t[126] = t[161] ^ x[36];
  assign t[127] = t[162] ^ x[35];
  assign t[128] = t[163] ^ x[37];
  assign t[129] = t[164] ^ x[38];
  assign t[12] = ~(t[18] ^ t[52]);
  assign t[130] = t[165] ^ x[39];
  assign t[131] = t[166] ^ x[33];
  assign t[132] = t[167] ^ x[50];
  assign t[133] = t[168] ^ x[45];
  assign t[134] = t[169] ^ x[46];
  assign t[135] = t[170] ^ x[47];
  assign t[136] = t[171] ^ x[51];
  assign t[137] = t[172] ^ x[48];
  assign t[138] = t[173] ^ x[49];
  assign t[139] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[141] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[142] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[143] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[144] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[145] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[146] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[147] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[148] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[149] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[14] = ~(t[53]);
  assign t[150] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[151] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[152] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[153] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[154] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[155] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[156] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[157] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[158] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~(t[51] ^ t[14]);
  assign t[160] = (x[29] & ~x[30] & ~x[31]) | (~x[29] & x[30] & ~x[31]) | (~x[29] & ~x[30] & x[31]) | (x[29] & x[30] & x[31]);
  assign t[161] = (x[29] & ~x[30] & ~x[32]) | (~x[29] & x[30] & ~x[32]) | (~x[29] & ~x[30] & x[32]) | (x[29] & x[30] & x[32]);
  assign t[162] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[163] = (x[29] & ~x[32]) | (~x[29] & x[32]);
  assign t[164] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[165] = (x[30] & ~x[32]) | (~x[30] & x[32]);
  assign t[166] = (x[31] & ~x[32]) | (~x[31] & x[32]);
  assign t[167] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[168] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[169] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[16] = t[54] ^ t[53];
  assign t[170] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[171] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[172] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[51] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[51] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[53] ^ t[55];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[56] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[57]);
  assign t[32] = ~(t[56] ^ t[31]);
  assign t[33] = t[58] ^ t[57];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[56] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[56] ^ t[38];
  assign t[38] = t[57] ^ t[59];
  assign t[39] = x[0] ? x[40] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44]);
  assign t[43] = ~(t[45] ^ t[60]);
  assign t[44] = t[23] ^ t[9];
  assign t[45] = ~t[46];
  assign t[46] = ~(t[47] ^ t[61]);
  assign t[47] = ~t[48];
  assign t[48] = ~(t[49]);
  assign t[49] = t[38] ^ t[27];
  assign t[4] = ~(t[7] ^ t[50]);
  assign t[50] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[51] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[64] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[64] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[54] = (t[64] & ~t[70]) | (~t[64] & t[70]);
  assign t[55] = (t[64] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[64] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[56] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[57] = (t[72] & ~t[75] & ~t[77]) | (~t[74] & t[75] & ~t[76]) | (~t[72] & ~t[75] & t[77]) | (t[74] & t[75] & t[76]);
  assign t[58] = (t[72] & ~t[76]) | (~t[72] & t[76]);
  assign t[59] = (t[72] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[77]) | (~t[72] & ~t[75] & t[76]) | (t[74] & t[75] & t[77]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[62] & ~t[79] & ~t[80]) | (~t[78] & t[79] & ~t[63]) | (~t[62] & ~t[79] & t[80]) | (t[78] & t[79] & t[63]);
  assign t[61] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[62] = t[83] ^ x[8];
  assign t[63] = t[84] ^ x[9];
  assign t[64] = t[85] ^ x[15];
  assign t[65] = t[86] ^ x[16];
  assign t[66] = t[87] ^ x[23];
  assign t[67] = t[88] ^ x[24];
  assign t[68] = t[89] ^ x[25];
  assign t[69] = t[90] ^ x[26];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[91] ^ x[27];
  assign t[71] = t[92] ^ x[28];
  assign t[72] = t[93] ^ x[34];
  assign t[73] = t[94] ^ x[35];
  assign t[74] = t[95] ^ x[36];
  assign t[75] = t[96] ^ x[37];
  assign t[76] = t[97] ^ x[38];
  assign t[77] = t[98] ^ x[39];
  assign t[78] = t[99] ^ x[41];
  assign t[79] = t[100] ^ x[42];
  assign t[7] = ~t[12];
  assign t[80] = t[101] ^ x[43];
  assign t[81] = t[102] ^ x[50];
  assign t[82] = t[103] ^ x[51];
  assign t[83] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[84] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (t[111] & ~t[112] & ~t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[112] & ~t[113] & ~t[116] & ~t[117]) | (~t[111] & t[112] & t[113] & t[114] & ~t[117]) | (~t[111] & t[112] & t[115] & t[116] & ~t[117]) | (t[111] & ~t[113] & ~t[115] & t[117]) | (~t[111] & t[113] & t[115] & t[117]);
  assign t[86] = (t[111] & t[112] & ~t[113] & t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[113] & ~t[114] & t[115] & ~t[116] & t[117]) | (~t[112] & t[113] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[112] & t[113] & ~t[116] & ~t[117]) | (~t[111] & t[113] & t[114] & ~t[115] & t[116]) | (t[113] & ~t[114] & t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[120] & ~t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[121] & ~t[122] & ~t[124]) | (t[118] & ~t[119] & ~t[120] & ~t[123] & ~t[124]) | (~t[118] & t[119] & t[120] & t[121] & ~t[124]) | (~t[118] & t[119] & t[122] & t[123] & ~t[124]) | (t[118] & ~t[120] & ~t[122] & t[124]) | (~t[118] & t[120] & t[122] & t[124]);
  assign t[88] = (t[118] & t[119] & ~t[120] & ~t[122] & t[123] & ~t[124]) | (t[118] & t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[124]) | (~t[118] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[118] & ~t[119] & ~t[121] & t[122] & ~t[124]) | (~t[118] & ~t[120] & t[121] & t[122] & t[123]) | (t[121] & t[122] & ~t[123] & ~t[124]);
  assign t[89] = (t[112] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & t[112] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[112] & ~t[113] & ~t[116] & ~t[117]) | (t[111] & ~t[112] & t[113] & t[114] & ~t[117]) | (t[111] & ~t[112] & t[115] & t[116] & ~t[117]) | (t[112] & ~t[114] & ~t[116] & t[117]) | (~t[112] & t[114] & t[116] & t[117]);
  assign t[8] = t[51] & t[13];
  assign t[90] = (t[111] & t[112] & t[113] & ~t[114] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[114] & ~t[115] & t[116] & t[117]) | (~t[112] & ~t[113] & t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[113] & t[114] & ~t[116] & ~t[117]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[117]) | (~t[112] & t[113] & t[114] & t[115] & ~t[116]) | (~t[113] & t[114] & t[115] & ~t[117]);
  assign t[91] = (t[111] & t[112] & ~t[113] & ~t[115] & t[116] & ~t[117]) | (t[111] & t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[117]) | (~t[111] & ~t[113] & ~t[114] & t[115] & ~t[116]) | (~t[111] & ~t[112] & ~t[114] & t[115] & ~t[117]) | (~t[111] & ~t[113] & t[114] & t[115] & t[116]) | (t[114] & t[115] & ~t[116] & ~t[117]);
  assign t[92] = (t[111] & t[112] & ~t[114] & t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[111] & ~t[112] & ~t[113] & t[116] & ~t[117]) | (~t[112] & t[113] & ~t[114] & t[115] & t[116]) | (t[113] & ~t[115] & t[116] & ~t[117]);
  assign t[93] = (t[125] & ~t[127] & ~t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[128] & ~t[129] & ~t[131]) | (t[125] & ~t[126] & ~t[127] & ~t[130] & ~t[131]) | (~t[125] & t[126] & t[127] & t[128] & ~t[131]) | (~t[125] & t[126] & t[129] & t[130] & ~t[131]) | (t[125] & ~t[127] & ~t[129] & t[131]) | (~t[125] & t[127] & t[129] & t[131]);
  assign t[94] = (t[125] & t[126] & ~t[127] & t[128] & ~t[129] & ~t[131]) | (t[125] & ~t[127] & ~t[128] & t[129] & ~t[130] & t[131]) | (~t[126] & t[127] & ~t[128] & ~t[129] & ~t[131]) | (~t[125] & t[127] & ~t[128] & ~t[129] & ~t[130]) | (~t[125] & ~t[126] & t[127] & ~t[130] & ~t[131]) | (~t[125] & t[127] & t[128] & ~t[129] & t[130]) | (t[127] & ~t[128] & t[130] & ~t[131]);
  assign t[95] = (t[126] & ~t[127] & ~t[128] & ~t[129] & ~t[130]) | (~t[125] & t[126] & ~t[128] & ~t[129] & ~t[131]) | (~t[125] & t[126] & ~t[127] & ~t[130] & ~t[131]) | (t[125] & ~t[126] & t[127] & t[128] & ~t[131]) | (t[125] & ~t[126] & t[129] & t[130] & ~t[131]) | (t[126] & ~t[128] & ~t[130] & t[131]) | (~t[126] & t[128] & t[130] & t[131]);
  assign t[96] = (t[125] & t[126] & t[127] & ~t[128] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & ~t[128] & ~t[129] & t[130] & t[131]) | (~t[126] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (~t[125] & ~t[127] & t[128] & ~t[130] & ~t[131]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[131]) | (~t[126] & t[127] & t[128] & t[129] & ~t[130]) | (~t[127] & t[128] & t[129] & ~t[131]);
  assign t[97] = (t[125] & t[126] & ~t[127] & ~t[129] & t[130] & ~t[131]) | (t[125] & t[127] & ~t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[127] & t[129] & ~t[130] & ~t[131]) | (~t[125] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[125] & ~t[126] & ~t[128] & t[129] & ~t[131]) | (~t[125] & ~t[127] & t[128] & t[129] & t[130]) | (t[128] & t[129] & ~t[130] & ~t[131]);
  assign t[98] = (t[125] & t[126] & ~t[128] & t[129] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[128] & ~t[129] & t[130] & ~t[131]) | (~t[125] & ~t[126] & ~t[127] & t[130] & ~t[131]) | (~t[126] & t[127] & ~t[128] & t[129] & t[130]) | (t[127] & ~t[129] & t[130] & ~t[131]);
  assign t[99] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind80(x, y);
 input [51:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[101] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[102] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[103] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[104] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[105] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[106] = t[141] ^ x[8];
  assign t[107] = t[142] ^ x[41];
  assign t[108] = t[143] ^ x[6];
  assign t[109] = t[144] ^ x[42];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[145] ^ x[9];
  assign t[111] = t[146] ^ x[43];
  assign t[112] = t[147] ^ x[7];
  assign t[113] = t[148] ^ x[15];
  assign t[114] = t[149] ^ x[25];
  assign t[115] = t[150] ^ x[16];
  assign t[116] = t[151] ^ x[26];
  assign t[117] = t[152] ^ x[27];
  assign t[118] = t[153] ^ x[28];
  assign t[119] = t[154] ^ x[14];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[155] ^ x[23];
  assign t[121] = t[156] ^ x[18];
  assign t[122] = t[157] ^ x[19];
  assign t[123] = t[158] ^ x[20];
  assign t[124] = t[159] ^ x[24];
  assign t[125] = t[160] ^ x[21];
  assign t[126] = t[161] ^ x[22];
  assign t[127] = t[162] ^ x[34];
  assign t[128] = t[163] ^ x[36];
  assign t[129] = t[164] ^ x[35];
  assign t[12] = ~(t[18] ^ t[54]);
  assign t[130] = t[165] ^ x[37];
  assign t[131] = t[166] ^ x[38];
  assign t[132] = t[167] ^ x[39];
  assign t[133] = t[168] ^ x[33];
  assign t[134] = t[169] ^ x[50];
  assign t[135] = t[170] ^ x[45];
  assign t[136] = t[171] ^ x[46];
  assign t[137] = t[172] ^ x[47];
  assign t[138] = t[173] ^ x[51];
  assign t[139] = t[174] ^ x[48];
  assign t[13] = t[19] ^ t[20];
  assign t[140] = t[175] ^ x[49];
  assign t[141] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[142] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[143] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[144] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[145] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[146] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[147] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[148] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[149] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[14] = ~(t[55]);
  assign t[150] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[151] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[152] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[153] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[154] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[155] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[156] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[157] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[158] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~(t[53] ^ t[14]);
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (x[29] & ~x[30] & ~x[31]) | (~x[29] & x[30] & ~x[31]) | (~x[29] & ~x[30] & x[31]) | (x[29] & x[30] & x[31]);
  assign t[163] = (x[29] & ~x[30] & ~x[32]) | (~x[29] & x[30] & ~x[32]) | (~x[29] & ~x[30] & x[32]) | (x[29] & x[30] & x[32]);
  assign t[164] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[165] = (x[29] & ~x[32]) | (~x[29] & x[32]);
  assign t[166] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[167] = (x[30] & ~x[32]) | (~x[30] & x[32]);
  assign t[168] = (x[31] & ~x[32]) | (~x[31] & x[32]);
  assign t[169] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[16] = t[56] ^ t[55];
  assign t[170] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[171] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[172] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[174] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[175] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[53] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[53] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[55] ^ t[57];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[58] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[59]);
  assign t[32] = ~(t[58] ^ t[31]);
  assign t[33] = t[60] ^ t[59];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[58] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[58] ^ t[38];
  assign t[38] = t[59] ^ t[61];
  assign t[39] = x[0] ? x[40] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44]);
  assign t[43] = ~(t[45] ^ t[62]);
  assign t[44] = t[46] ^ t[9];
  assign t[45] = ~t[47];
  assign t[46] = t[16] ^ t[20];
  assign t[47] = ~(t[48] ^ t[63]);
  assign t[48] = ~t[49];
  assign t[49] = ~(t[50]);
  assign t[4] = ~(t[7] ^ t[52]);
  assign t[50] = t[51] ^ t[27];
  assign t[51] = t[33] ^ t[36];
  assign t[52] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[53] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[54] = (t[68] & ~t[69]) | (~t[68] & t[69]);
  assign t[55] = (t[66] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[66] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = (t[66] & ~t[72]) | (~t[66] & t[72]);
  assign t[57] = (t[66] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[73]) | (~t[66] & ~t[71] & t[72]) | (t[70] & t[71] & t[73]);
  assign t[58] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[59] = (t[74] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[74] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[74] & ~t[78]) | (~t[74] & t[78]);
  assign t[61] = (t[74] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[74] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[62] = (t[64] & ~t[81] & ~t[65]) | (~t[80] & t[81] & ~t[82]) | (~t[64] & ~t[81] & t[65]) | (t[80] & t[81] & t[82]);
  assign t[63] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[64] = t[85] ^ x[8];
  assign t[65] = t[86] ^ x[9];
  assign t[66] = t[87] ^ x[15];
  assign t[67] = t[88] ^ x[16];
  assign t[68] = t[89] ^ x[23];
  assign t[69] = t[90] ^ x[24];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[91] ^ x[25];
  assign t[71] = t[92] ^ x[26];
  assign t[72] = t[93] ^ x[27];
  assign t[73] = t[94] ^ x[28];
  assign t[74] = t[95] ^ x[34];
  assign t[75] = t[96] ^ x[35];
  assign t[76] = t[97] ^ x[36];
  assign t[77] = t[98] ^ x[37];
  assign t[78] = t[99] ^ x[38];
  assign t[79] = t[100] ^ x[39];
  assign t[7] = ~t[12];
  assign t[80] = t[101] ^ x[41];
  assign t[81] = t[102] ^ x[42];
  assign t[82] = t[103] ^ x[43];
  assign t[83] = t[104] ^ x[50];
  assign t[84] = t[105] ^ x[51];
  assign t[85] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[86] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[87] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[88] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[8] = t[53] & t[13];
  assign t[90] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[91] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[92] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[93] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[94] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[95] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[96] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[97] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[98] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[99] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind81(x, y);
 input [51:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[101] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[102] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[103] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[104] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[105] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[106] = t[141] ^ x[7];
  assign t[107] = t[142] ^ x[40];
  assign t[108] = t[143] ^ x[8];
  assign t[109] = t[144] ^ x[41];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[145] ^ x[42];
  assign t[111] = t[146] ^ x[43];
  assign t[112] = t[147] ^ x[6];
  assign t[113] = t[148] ^ x[14];
  assign t[114] = t[149] ^ x[25];
  assign t[115] = t[150] ^ x[15];
  assign t[116] = t[151] ^ x[26];
  assign t[117] = t[152] ^ x[24];
  assign t[118] = t[153] ^ x[27];
  assign t[119] = t[154] ^ x[13];
  assign t[11] = t[51] ^ t[15];
  assign t[120] = t[155] ^ x[22];
  assign t[121] = t[156] ^ x[17];
  assign t[122] = t[157] ^ x[18];
  assign t[123] = t[158] ^ x[19];
  assign t[124] = t[159] ^ x[23];
  assign t[125] = t[160] ^ x[20];
  assign t[126] = t[161] ^ x[21];
  assign t[127] = t[162] ^ x[33];
  assign t[128] = t[163] ^ x[36];
  assign t[129] = t[164] ^ x[34];
  assign t[12] = ~(t[18] ^ t[52]);
  assign t[130] = t[165] ^ x[37];
  assign t[131] = t[166] ^ x[35];
  assign t[132] = t[167] ^ x[38];
  assign t[133] = t[168] ^ x[32];
  assign t[134] = t[169] ^ x[50];
  assign t[135] = t[170] ^ x[45];
  assign t[136] = t[171] ^ x[46];
  assign t[137] = t[172] ^ x[47];
  assign t[138] = t[173] ^ x[51];
  assign t[139] = t[174] ^ x[48];
  assign t[13] = t[53] ^ t[54];
  assign t[140] = t[175] ^ x[49];
  assign t[141] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[142] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[143] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[144] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[145] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[146] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[147] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[148] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[149] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[14] = t[15] & t[19];
  assign t[150] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[151] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[152] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[153] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[154] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[155] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[156] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[157] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[158] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~(t[54]);
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[162] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[163] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[164] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[165] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[166] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[167] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[168] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[169] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[16] = ~(t[51] ^ t[15]);
  assign t[170] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[171] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[172] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[174] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[175] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[17] = t[51] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[51] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[54] ^ t[55];
  assign t[23] = t[51] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[56] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[57] ^ t[58];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[58]);
  assign t[33] = ~(t[56] ^ t[32]);
  assign t[34] = t[56] & t[36];
  assign t[35] = t[56] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[56] ^ t[30];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44]);
  assign t[43] = ~(t[45] ^ t[60]);
  assign t[44] = t[22] ^ t[9];
  assign t[45] = ~t[46];
  assign t[46] = ~(t[47] ^ t[61]);
  assign t[47] = ~t[48];
  assign t[48] = ~(t[49]);
  assign t[49] = t[37] ^ t[27];
  assign t[4] = ~(t[7] ^ t[50]);
  assign t[50] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[51] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[70] & ~t[71]) | (~t[69] & t[70] & ~t[68]) | (~t[64] & ~t[70] & t[71]) | (t[69] & t[70] & t[68]);
  assign t[55] = (t[64] & ~t[70] & ~t[68]) | (~t[69] & t[70] & ~t[71]) | (~t[64] & ~t[70] & t[68]) | (t[69] & t[70] & t[71]);
  assign t[56] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[57] = (t[72] & ~t[74]) | (~t[72] & t[74]);
  assign t[58] = (t[72] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[74]) | (~t[72] & ~t[76] & t[77]) | (t[75] & t[76] & t[74]);
  assign t[59] = (t[72] & ~t[76] & ~t[74]) | (~t[75] & t[76] & ~t[77]) | (~t[72] & ~t[76] & t[74]) | (t[75] & t[76] & t[77]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[62] & ~t[79] & ~t[81]) | (~t[78] & t[79] & ~t[80]) | (~t[62] & ~t[79] & t[81]) | (t[78] & t[79] & t[80]);
  assign t[61] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[62] = t[84] ^ x[7];
  assign t[63] = t[85] ^ x[8];
  assign t[64] = t[86] ^ x[14];
  assign t[65] = t[87] ^ x[15];
  assign t[66] = t[88] ^ x[22];
  assign t[67] = t[89] ^ x[23];
  assign t[68] = t[90] ^ x[24];
  assign t[69] = t[91] ^ x[25];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[92] ^ x[26];
  assign t[71] = t[93] ^ x[27];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[34];
  assign t[74] = t[96] ^ x[35];
  assign t[75] = t[97] ^ x[36];
  assign t[76] = t[98] ^ x[37];
  assign t[77] = t[99] ^ x[38];
  assign t[78] = t[100] ^ x[40];
  assign t[79] = t[101] ^ x[41];
  assign t[7] = ~t[12];
  assign t[80] = t[102] ^ x[42];
  assign t[81] = t[103] ^ x[43];
  assign t[82] = t[104] ^ x[50];
  assign t[83] = t[105] ^ x[51];
  assign t[84] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[85] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[87] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[89] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[91] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[92] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[93] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[94] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[95] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[96] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[97] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[98] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[99] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind82(x, y);
 input [51:0] x;
 output y;

 wire [173:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[101] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[102] = (t[132] & ~t[134] & ~t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[135] & ~t[136] & ~t[138]) | (t[132] & ~t[133] & ~t[134] & ~t[137] & ~t[138]) | (~t[132] & t[133] & t[134] & t[135] & ~t[138]) | (~t[132] & t[133] & t[136] & t[137] & ~t[138]) | (t[132] & ~t[134] & ~t[136] & t[138]) | (~t[132] & t[134] & t[136] & t[138]);
  assign t[103] = (t[132] & t[133] & ~t[134] & ~t[136] & t[137] & ~t[138]) | (t[132] & t[134] & ~t[135] & ~t[136] & ~t[137] & t[138]) | (~t[133] & ~t[134] & t[136] & ~t[137] & ~t[138]) | (~t[132] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[132] & ~t[133] & ~t[135] & t[136] & ~t[138]) | (~t[132] & ~t[134] & t[135] & t[136] & t[137]) | (t[135] & t[136] & ~t[137] & ~t[138]);
  assign t[104] = t[139] ^ x[7];
  assign t[105] = t[140] ^ x[40];
  assign t[106] = t[141] ^ x[8];
  assign t[107] = t[142] ^ x[41];
  assign t[108] = t[143] ^ x[42];
  assign t[109] = t[144] ^ x[43];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[145] ^ x[6];
  assign t[111] = t[146] ^ x[14];
  assign t[112] = t[147] ^ x[25];
  assign t[113] = t[148] ^ x[15];
  assign t[114] = t[149] ^ x[26];
  assign t[115] = t[150] ^ x[24];
  assign t[116] = t[151] ^ x[27];
  assign t[117] = t[152] ^ x[13];
  assign t[118] = t[153] ^ x[22];
  assign t[119] = t[154] ^ x[17];
  assign t[11] = t[49] ^ t[15];
  assign t[120] = t[155] ^ x[18];
  assign t[121] = t[156] ^ x[19];
  assign t[122] = t[157] ^ x[23];
  assign t[123] = t[158] ^ x[20];
  assign t[124] = t[159] ^ x[21];
  assign t[125] = t[160] ^ x[33];
  assign t[126] = t[161] ^ x[36];
  assign t[127] = t[162] ^ x[34];
  assign t[128] = t[163] ^ x[37];
  assign t[129] = t[164] ^ x[35];
  assign t[12] = ~(t[18] ^ t[50]);
  assign t[130] = t[165] ^ x[38];
  assign t[131] = t[166] ^ x[32];
  assign t[132] = t[167] ^ x[50];
  assign t[133] = t[168] ^ x[45];
  assign t[134] = t[169] ^ x[46];
  assign t[135] = t[170] ^ x[47];
  assign t[136] = t[171] ^ x[51];
  assign t[137] = t[172] ^ x[48];
  assign t[138] = t[173] ^ x[49];
  assign t[139] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[13] = t[51] ^ t[52];
  assign t[140] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[141] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[142] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[143] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[144] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[145] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[146] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[147] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[148] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[149] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[14] = t[15] & t[19];
  assign t[150] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[151] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[152] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[153] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[154] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[155] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[156] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[157] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[158] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = ~(t[52]);
  assign t[160] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[161] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[162] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[163] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[164] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[165] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[166] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[167] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[168] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[169] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[16] = ~(t[49] ^ t[15]);
  assign t[170] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[171] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[172] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[17] = t[49] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[49] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[52] ^ t[53];
  assign t[23] = t[49] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[54] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[55] ^ t[56];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[56]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[36];
  assign t[35] = t[54] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[56] ^ t[57];
  assign t[38] = t[54] ^ t[30];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[5]);
  assign t[43] = ~(t[44] ^ t[58]);
  assign t[44] = ~t[45];
  assign t[45] = ~(t[46] ^ t[59]);
  assign t[46] = ~t[47];
  assign t[47] = ~(t[24]);
  assign t[48] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[49] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[62] & ~t[66]) | (~t[62] & t[66]);
  assign t[52] = (t[62] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[66]) | (~t[62] & ~t[68] & t[69]) | (t[67] & t[68] & t[66]);
  assign t[53] = (t[62] & ~t[68] & ~t[66]) | (~t[67] & t[68] & ~t[69]) | (~t[62] & ~t[68] & t[66]) | (t[67] & t[68] & t[69]);
  assign t[54] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[55] = (t[70] & ~t[72]) | (~t[70] & t[72]);
  assign t[56] = (t[70] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[72]) | (~t[70] & ~t[74] & t[75]) | (t[73] & t[74] & t[72]);
  assign t[57] = (t[70] & ~t[74] & ~t[72]) | (~t[73] & t[74] & ~t[75]) | (~t[70] & ~t[74] & t[72]) | (t[73] & t[74] & t[75]);
  assign t[58] = (t[60] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[60] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[59] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[82] ^ x[7];
  assign t[61] = t[83] ^ x[8];
  assign t[62] = t[84] ^ x[14];
  assign t[63] = t[85] ^ x[15];
  assign t[64] = t[86] ^ x[22];
  assign t[65] = t[87] ^ x[23];
  assign t[66] = t[88] ^ x[24];
  assign t[67] = t[89] ^ x[25];
  assign t[68] = t[90] ^ x[26];
  assign t[69] = t[91] ^ x[27];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[34];
  assign t[72] = t[94] ^ x[35];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[37];
  assign t[75] = t[97] ^ x[38];
  assign t[76] = t[98] ^ x[40];
  assign t[77] = t[99] ^ x[41];
  assign t[78] = t[100] ^ x[42];
  assign t[79] = t[101] ^ x[43];
  assign t[7] = ~t[12];
  assign t[80] = t[102] ^ x[50];
  assign t[81] = t[103] ^ x[51];
  assign t[82] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[83] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[84] = (t[111] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (t[111] & ~t[112] & ~t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[112] & ~t[113] & ~t[116] & ~t[117]) | (~t[111] & t[112] & t[113] & t[114] & ~t[117]) | (~t[111] & t[112] & t[115] & t[116] & ~t[117]) | (t[111] & ~t[113] & ~t[115] & t[117]) | (~t[111] & t[113] & t[115] & t[117]);
  assign t[85] = (t[111] & t[112] & ~t[113] & t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[113] & ~t[114] & t[115] & ~t[116] & t[117]) | (~t[112] & t[113] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[112] & t[113] & ~t[116] & ~t[117]) | (~t[111] & t[113] & t[114] & ~t[115] & t[116]) | (t[113] & ~t[114] & t[116] & ~t[117]);
  assign t[86] = (t[118] & ~t[120] & ~t[121] & ~t[122] & ~t[123]) | (t[118] & ~t[119] & ~t[121] & ~t[122] & ~t[124]) | (t[118] & ~t[119] & ~t[120] & ~t[123] & ~t[124]) | (~t[118] & t[119] & t[120] & t[121] & ~t[124]) | (~t[118] & t[119] & t[122] & t[123] & ~t[124]) | (t[118] & ~t[120] & ~t[122] & t[124]) | (~t[118] & t[120] & t[122] & t[124]);
  assign t[87] = (t[118] & t[119] & ~t[120] & ~t[122] & t[123] & ~t[124]) | (t[118] & t[120] & ~t[121] & ~t[122] & ~t[123] & t[124]) | (~t[119] & ~t[120] & t[122] & ~t[123] & ~t[124]) | (~t[118] & ~t[120] & ~t[121] & t[122] & ~t[123]) | (~t[118] & ~t[119] & ~t[121] & t[122] & ~t[124]) | (~t[118] & ~t[120] & t[121] & t[122] & t[123]) | (t[121] & t[122] & ~t[123] & ~t[124]);
  assign t[88] = (t[111] & t[112] & ~t[113] & ~t[115] & t[116] & ~t[117]) | (t[111] & t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[117]) | (~t[111] & ~t[113] & ~t[114] & t[115] & ~t[116]) | (~t[111] & ~t[112] & ~t[114] & t[115] & ~t[117]) | (~t[111] & ~t[113] & t[114] & t[115] & t[116]) | (t[114] & t[115] & ~t[116] & ~t[117]);
  assign t[89] = (t[112] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (~t[111] & t[112] & ~t[114] & ~t[115] & ~t[117]) | (~t[111] & t[112] & ~t[113] & ~t[116] & ~t[117]) | (t[111] & ~t[112] & t[113] & t[114] & ~t[117]) | (t[111] & ~t[112] & t[115] & t[116] & ~t[117]) | (t[112] & ~t[114] & ~t[116] & t[117]) | (~t[112] & t[114] & t[116] & t[117]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[111] & t[112] & t[113] & ~t[114] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[114] & ~t[115] & t[116] & t[117]) | (~t[112] & ~t[113] & t[114] & ~t[115] & ~t[116]) | (~t[111] & ~t[113] & t[114] & ~t[116] & ~t[117]) | (~t[111] & ~t[112] & t[114] & ~t[115] & ~t[117]) | (~t[112] & t[113] & t[114] & t[115] & ~t[116]) | (~t[113] & t[114] & t[115] & ~t[117]);
  assign t[91] = (t[111] & t[112] & ~t[114] & t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & ~t[114] & ~t[115] & t[116]) | (~t[111] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[111] & ~t[112] & ~t[113] & t[116] & ~t[117]) | (~t[112] & t[113] & ~t[114] & t[115] & t[116]) | (t[113] & ~t[115] & t[116] & ~t[117]);
  assign t[92] = (t[125] & ~t[127] & ~t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[128] & ~t[129] & ~t[131]) | (t[125] & ~t[126] & ~t[127] & ~t[130] & ~t[131]) | (~t[125] & t[126] & t[127] & t[128] & ~t[131]) | (~t[125] & t[126] & t[129] & t[130] & ~t[131]) | (t[125] & ~t[127] & ~t[129] & t[131]) | (~t[125] & t[127] & t[129] & t[131]);
  assign t[93] = (t[125] & t[126] & ~t[127] & t[128] & ~t[129] & ~t[131]) | (t[125] & ~t[127] & ~t[128] & t[129] & ~t[130] & t[131]) | (~t[126] & t[127] & ~t[128] & ~t[129] & ~t[131]) | (~t[125] & t[127] & ~t[128] & ~t[129] & ~t[130]) | (~t[125] & ~t[126] & t[127] & ~t[130] & ~t[131]) | (~t[125] & t[127] & t[128] & ~t[129] & t[130]) | (t[127] & ~t[128] & t[130] & ~t[131]);
  assign t[94] = (t[125] & t[126] & ~t[127] & ~t[129] & t[130] & ~t[131]) | (t[125] & t[127] & ~t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[127] & t[129] & ~t[130] & ~t[131]) | (~t[125] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[125] & ~t[126] & ~t[128] & t[129] & ~t[131]) | (~t[125] & ~t[127] & t[128] & t[129] & t[130]) | (t[128] & t[129] & ~t[130] & ~t[131]);
  assign t[95] = (t[126] & ~t[127] & ~t[128] & ~t[129] & ~t[130]) | (~t[125] & t[126] & ~t[128] & ~t[129] & ~t[131]) | (~t[125] & t[126] & ~t[127] & ~t[130] & ~t[131]) | (t[125] & ~t[126] & t[127] & t[128] & ~t[131]) | (t[125] & ~t[126] & t[129] & t[130] & ~t[131]) | (t[126] & ~t[128] & ~t[130] & t[131]) | (~t[126] & t[128] & t[130] & t[131]);
  assign t[96] = (t[125] & t[126] & t[127] & ~t[128] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & ~t[128] & ~t[129] & t[130] & t[131]) | (~t[126] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (~t[125] & ~t[127] & t[128] & ~t[130] & ~t[131]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[131]) | (~t[126] & t[127] & t[128] & t[129] & ~t[130]) | (~t[127] & t[128] & t[129] & ~t[131]);
  assign t[97] = (t[125] & t[126] & ~t[128] & t[129] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[128] & ~t[129] & t[130] & ~t[131]) | (~t[125] & ~t[126] & ~t[127] & t[130] & ~t[131]) | (~t[126] & t[127] & ~t[128] & t[129] & t[130]) | (t[127] & ~t[129] & t[130] & ~t[131]);
  assign t[98] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[99] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind83(x, y);
 input [51:0] x;
 output y;

 wire [161:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[135] ^ x[19];
  assign t[101] = t[136] ^ x[31];
  assign t[102] = t[137] ^ x[20];
  assign t[103] = t[138] ^ x[21];
  assign t[104] = t[139] ^ x[22];
  assign t[105] = t[140] ^ x[17];
  assign t[106] = t[141] ^ x[29];
  assign t[107] = t[142] ^ x[24];
  assign t[108] = t[143] ^ x[25];
  assign t[109] = t[144] ^ x[26];
  assign t[10] = ~(t[39]);
  assign t[110] = t[145] ^ x[30];
  assign t[111] = t[146] ^ x[27];
  assign t[112] = t[147] ^ x[28];
  assign t[113] = t[148] ^ x[37];
  assign t[114] = t[149] ^ x[38];
  assign t[115] = t[150] ^ x[42];
  assign t[116] = t[151] ^ x[39];
  assign t[117] = t[152] ^ x[40];
  assign t[118] = t[153] ^ x[41];
  assign t[119] = t[154] ^ x[36];
  assign t[11] = ~(t[42] ^ t[10]);
  assign t[120] = t[155] ^ x[50];
  assign t[121] = t[156] ^ x[45];
  assign t[122] = t[157] ^ x[46];
  assign t[123] = t[158] ^ x[47];
  assign t[124] = t[159] ^ x[51];
  assign t[125] = t[160] ^ x[48];
  assign t[126] = t[161] ^ x[49];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = ~t[13];
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[135] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[136] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[137] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[138] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[139] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[13] = ~(t[14]);
  assign t[140] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[141] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[142] = (x[23] & ~1'b0 & ~1'b0) | (~x[23] & 1'b0 & ~1'b0) | (~x[23] & ~1'b0 & 1'b0) | (x[23] & 1'b0 & 1'b0);
  assign t[143] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[144] = (x[23] & ~1'b0) | (~x[23] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[32] & ~x[33] & ~x[34]) | (~x[32] & x[33] & ~x[34]) | (~x[32] & ~x[33] & x[34]) | (x[32] & x[33] & x[34]);
  assign t[149] = (x[32] & ~x[33] & ~x[35]) | (~x[32] & x[33] & ~x[35]) | (~x[32] & ~x[33] & x[35]) | (x[32] & x[33] & x[35]);
  assign t[14] = t[15] ^ t[16];
  assign t[150] = (x[32] & ~x[34]) | (~x[32] & x[34]);
  assign t[151] = (x[32] & ~x[35]) | (~x[32] & x[35]);
  assign t[152] = (x[33] & ~x[34]) | (~x[33] & x[34]);
  assign t[153] = (x[33] & ~x[35]) | (~x[33] & x[35]);
  assign t[154] = (x[34] & ~x[35]) | (~x[34] & x[35]);
  assign t[155] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[156] = (x[44] & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0);
  assign t[157] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[158] = (x[44] & ~1'b0) | (~x[44] & 1'b0);
  assign t[159] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = t[43] ^ t[44];
  assign t[160] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[161] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[43]);
  assign t[18] = ~(t[45] ^ t[17]);
  assign t[19] = x[0] ? x[43] : t[20];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = ~t[23];
  assign t[22] = ~(t[24]);
  assign t[23] = ~(t[25] ^ t[46]);
  assign t[24] = t[26] ^ t[8];
  assign t[25] = ~t[27];
  assign t[26] = t[28] ^ t[29];
  assign t[27] = ~(t[30] ^ t[47]);
  assign t[28] = t[48] ^ t[39];
  assign t[29] = t[10] & t[31];
  assign t[2] = ~t[4];
  assign t[30] = ~t[32];
  assign t[31] = t[42] ^ t[7];
  assign t[32] = ~(t[33]);
  assign t[33] = t[34] ^ t[16];
  assign t[34] = t[35] ^ t[36];
  assign t[35] = t[49] ^ t[43];
  assign t[36] = t[17] & t[37];
  assign t[37] = t[45] ^ t[15];
  assign t[38] = (t[50] & ~t[52] & ~t[54]) | (~t[51] & t[52] & ~t[53]) | (~t[50] & ~t[52] & t[54]) | (t[51] & t[52] & t[53]);
  assign t[39] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[41] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[42] = (t[55] & ~t[62]) | (~t[55] & t[62]);
  assign t[43] = (t[63] & ~t[65] & ~t[67]) | (~t[64] & t[65] & ~t[66]) | (~t[63] & ~t[65] & t[67]) | (t[64] & t[65] & t[66]);
  assign t[44] = (t[63] & ~t[65] & ~t[66]) | (~t[64] & t[65] & ~t[67]) | (~t[63] & ~t[65] & t[66]) | (t[64] & t[65] & t[67]);
  assign t[45] = (t[63] & ~t[68]) | (~t[63] & t[68]);
  assign t[46] = (t[50] & ~t[52] & ~t[53]) | (~t[51] & t[52] & ~t[54]) | (~t[50] & ~t[52] & t[53]) | (t[51] & t[52] & t[54]);
  assign t[47] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[48] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[49] = (t[63] & ~t[66]) | (~t[63] & t[66]);
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[71] ^ x[8];
  assign t[51] = t[72] ^ x[9];
  assign t[52] = t[73] ^ x[10];
  assign t[53] = t[74] ^ x[11];
  assign t[54] = t[75] ^ x[12];
  assign t[55] = t[76] ^ x[18];
  assign t[56] = t[77] ^ x[19];
  assign t[57] = t[78] ^ x[20];
  assign t[58] = t[79] ^ x[21];
  assign t[59] = t[80] ^ x[22];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[81] ^ x[29];
  assign t[61] = t[82] ^ x[30];
  assign t[62] = t[83] ^ x[31];
  assign t[63] = t[84] ^ x[37];
  assign t[64] = t[85] ^ x[38];
  assign t[65] = t[86] ^ x[39];
  assign t[66] = t[87] ^ x[40];
  assign t[67] = t[88] ^ x[41];
  assign t[68] = t[89] ^ x[42];
  assign t[69] = t[90] ^ x[50];
  assign t[6] = ~t[9];
  assign t[70] = t[91] ^ x[51];
  assign t[71] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[72] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[73] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[74] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[78] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[79] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[7] = t[39] ^ t[40];
  assign t[80] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[82] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[83] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[84] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[85] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[86] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[87] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[88] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[89] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[8] = t[10] & t[11];
  assign t[90] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[91] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[92] = t[127] ^ x[8];
  assign t[93] = t[128] ^ x[9];
  assign t[94] = t[129] ^ x[6];
  assign t[95] = t[130] ^ x[10];
  assign t[96] = t[131] ^ x[11];
  assign t[97] = t[132] ^ x[12];
  assign t[98] = t[133] ^ x[7];
  assign t[99] = t[134] ^ x[18];
  assign t[9] = ~(t[12] ^ t[41]);
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind84(x, y);
 input [36:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[101] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[102] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[103] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[104] = (t[108] & t[109] & ~t[110] & t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[110] & ~t[111] & t[112] & ~t[113] & t[114]) | (~t[109] & t[110] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[109] & t[110] & ~t[113] & ~t[114]) | (~t[108] & t[110] & t[111] & ~t[112] & t[113]) | (t[110] & ~t[111] & t[113] & ~t[114]);
  assign t[105] = (t[109] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & t[109] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[109] & ~t[110] & ~t[113] & ~t[114]) | (t[108] & ~t[109] & t[110] & t[111] & ~t[114]) | (t[108] & ~t[109] & t[112] & t[113] & ~t[114]) | (t[109] & ~t[111] & ~t[113] & t[114]) | (~t[109] & t[111] & t[113] & t[114]);
  assign t[106] = (t[108] & t[109] & t[110] & ~t[111] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[111] & ~t[112] & t[113] & t[114]) | (~t[109] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[110] & t[111] & ~t[113] & ~t[114]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[114]) | (~t[109] & t[110] & t[111] & t[112] & ~t[113]) | (~t[110] & t[111] & t[112] & ~t[114]);
  assign t[107] = (t[108] & t[109] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[108] & ~t[109] & ~t[110] & t[113] & ~t[114]) | (~t[109] & t[110] & ~t[111] & t[112] & t[113]) | (t[110] & ~t[112] & t[113] & ~t[114]);
  assign t[108] = t[129] ^ x[7];
  assign t[109] = t[130] ^ x[34];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[32];
  assign t[111] = t[132] ^ x[35];
  assign t[112] = t[133] ^ x[8];
  assign t[113] = t[134] ^ x[36];
  assign t[114] = t[135] ^ x[6];
  assign t[115] = t[136] ^ x[14];
  assign t[116] = t[137] ^ x[16];
  assign t[117] = t[138] ^ x[15];
  assign t[118] = t[139] ^ x[17];
  assign t[119] = t[140] ^ x[18];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[19];
  assign t[121] = t[142] ^ x[13];
  assign t[122] = t[143] ^ x[25];
  assign t[123] = t[144] ^ x[27];
  assign t[124] = t[145] ^ x[26];
  assign t[125] = t[146] ^ x[28];
  assign t[126] = t[147] ^ x[29];
  assign t[127] = t[148] ^ x[30];
  assign t[128] = t[149] ^ x[24];
  assign t[129] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[131] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[132] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[133] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[134] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[135] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[136] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[137] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[138] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[139] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[141] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[142] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[143] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[144] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[145] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[146] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[147] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[148] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[149] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[63]);
  assign t[15] = ~(t[62] ^ t[14]);
  assign t[16] = t[64] ^ t[63];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[62] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[62] ^ t[27];
  assign t[23] = t[65] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[63] ^ t[66];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[67]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[65] ^ t[29]);
  assign t[31] = t[68] ^ t[67];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[65] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[65] ^ t[36];
  assign t[36] = t[67] ^ t[69];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[70]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[62] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[61]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[65] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[71]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[62] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[63] = (t[74] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[74] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[64] = (t[74] & ~t[78]) | (~t[74] & t[78]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[74] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[74] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[67] = (t[80] & ~t[83] & ~t[85]) | (~t[82] & t[83] & ~t[84]) | (~t[80] & ~t[83] & t[85]) | (t[82] & t[83] & t[84]);
  assign t[68] = (t[80] & ~t[84]) | (~t[80] & t[84]);
  assign t[69] = (t[80] & ~t[83] & ~t[84]) | (~t[82] & t[83] & ~t[85]) | (~t[80] & ~t[83] & t[84]) | (t[82] & t[83] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[72] & ~t[86]) | (~t[72] & t[86]);
  assign t[71] = (t[72] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[73]) | (~t[72] & ~t[88] & t[89]) | (t[87] & t[88] & t[73]);
  assign t[72] = t[90] ^ x[7];
  assign t[73] = t[91] ^ x[8];
  assign t[74] = t[92] ^ x[14];
  assign t[75] = t[93] ^ x[15];
  assign t[76] = t[94] ^ x[16];
  assign t[77] = t[95] ^ x[17];
  assign t[78] = t[96] ^ x[18];
  assign t[79] = t[97] ^ x[19];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[25];
  assign t[81] = t[99] ^ x[26];
  assign t[82] = t[100] ^ x[27];
  assign t[83] = t[101] ^ x[28];
  assign t[84] = t[102] ^ x[29];
  assign t[85] = t[103] ^ x[30];
  assign t[86] = t[104] ^ x[32];
  assign t[87] = t[105] ^ x[34];
  assign t[88] = t[106] ^ x[35];
  assign t[89] = t[107] ^ x[36];
  assign t[8] = t[62] & t[13];
  assign t[90] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[91] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[92] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[93] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[94] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[95] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[96] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[97] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[98] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[99] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind85(x, y);
 input [36:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[101] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[102] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[103] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[104] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[105] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[106] = t[127] ^ x[7];
  assign t[107] = t[128] ^ x[34];
  assign t[108] = t[129] ^ x[32];
  assign t[109] = t[130] ^ x[35];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[8];
  assign t[111] = t[132] ^ x[36];
  assign t[112] = t[133] ^ x[6];
  assign t[113] = t[134] ^ x[14];
  assign t[114] = t[135] ^ x[16];
  assign t[115] = t[136] ^ x[15];
  assign t[116] = t[137] ^ x[17];
  assign t[117] = t[138] ^ x[18];
  assign t[118] = t[139] ^ x[19];
  assign t[119] = t[140] ^ x[13];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[25];
  assign t[121] = t[142] ^ x[27];
  assign t[122] = t[143] ^ x[26];
  assign t[123] = t[144] ^ x[28];
  assign t[124] = t[145] ^ x[29];
  assign t[125] = t[146] ^ x[30];
  assign t[126] = t[147] ^ x[24];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[135] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[136] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[137] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[138] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[139] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[141] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[142] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[143] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[144] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[145] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[146] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[147] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[61]);
  assign t[15] = ~(t[60] ^ t[14]);
  assign t[16] = t[62] ^ t[61];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[60] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[60] ^ t[27];
  assign t[23] = t[63] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[61] ^ t[64];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[65]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[63] ^ t[29]);
  assign t[31] = t[66] ^ t[65];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[63] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[63] ^ t[36];
  assign t[36] = t[65] ^ t[67];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[68]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[60] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[59]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[63] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[42]);
  assign t[56] = ~(t[57] ^ t[69]);
  assign t[57] = ~t[58];
  assign t[58] = ~(t[48]);
  assign t[59] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[61] = (t[72] & ~t[75] & ~t[77]) | (~t[74] & t[75] & ~t[76]) | (~t[72] & ~t[75] & t[77]) | (t[74] & t[75] & t[76]);
  assign t[62] = (t[72] & ~t[76]) | (~t[72] & t[76]);
  assign t[63] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[64] = (t[72] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[77]) | (~t[72] & ~t[75] & t[76]) | (t[74] & t[75] & t[77]);
  assign t[65] = (t[78] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[78] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[66] = (t[78] & ~t[82]) | (~t[78] & t[82]);
  assign t[67] = (t[78] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[78] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[68] = (t[70] & ~t[84]) | (~t[70] & t[84]);
  assign t[69] = (t[70] & ~t[86] & ~t[71]) | (~t[85] & t[86] & ~t[87]) | (~t[70] & ~t[86] & t[71]) | (t[85] & t[86] & t[87]);
  assign t[6] = t[10] & t[11];
  assign t[70] = t[88] ^ x[7];
  assign t[71] = t[89] ^ x[8];
  assign t[72] = t[90] ^ x[14];
  assign t[73] = t[91] ^ x[15];
  assign t[74] = t[92] ^ x[16];
  assign t[75] = t[93] ^ x[17];
  assign t[76] = t[94] ^ x[18];
  assign t[77] = t[95] ^ x[19];
  assign t[78] = t[96] ^ x[25];
  assign t[79] = t[97] ^ x[26];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[27];
  assign t[81] = t[99] ^ x[28];
  assign t[82] = t[100] ^ x[29];
  assign t[83] = t[101] ^ x[30];
  assign t[84] = t[102] ^ x[32];
  assign t[85] = t[103] ^ x[34];
  assign t[86] = t[104] ^ x[35];
  assign t[87] = t[105] ^ x[36];
  assign t[88] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[89] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[8] = t[60] & t[13];
  assign t[90] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[93] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[96] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[97] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[98] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[99] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind86(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[19];
  assign t[102] = t[123] ^ x[20];
  assign t[103] = t[124] ^ x[14];
  assign t[104] = t[125] ^ x[26];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[27];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[30];
  assign t[109] = t[130] ^ x[31];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[25];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[119] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[121] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[122] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[123] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[124] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[125] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[126] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[127] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[128] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[129] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[131] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[48]);
  assign t[15] = ~(t[47] ^ t[14]);
  assign t[16] = t[49] ^ t[48];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[47] ^ t[27];
  assign t[23] = t[50] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[48] ^ t[51];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[52]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[50] ^ t[29]);
  assign t[31] = t[53] ^ t[52];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[50] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[50] ^ t[36];
  assign t[36] = t[52] ^ t[54];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[27] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[36] ^ t[24];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[58] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[49] = (t[58] & ~t[62]) | (~t[58] & t[62]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[58] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[52] = (t[64] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[64] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[64] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[57]) | (~t[56] & ~t[71] & t[72]) | (t[70] & t[71] & t[57]);
  assign t[56] = t[73] ^ x[8];
  assign t[57] = t[74] ^ x[9];
  assign t[58] = t[75] ^ x[15];
  assign t[59] = t[76] ^ x[16];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[17];
  assign t[61] = t[78] ^ x[18];
  assign t[62] = t[79] ^ x[19];
  assign t[63] = t[80] ^ x[20];
  assign t[64] = t[81] ^ x[26];
  assign t[65] = t[82] ^ x[27];
  assign t[66] = t[83] ^ x[28];
  assign t[67] = t[84] ^ x[29];
  assign t[68] = t[85] ^ x[30];
  assign t[69] = t[86] ^ x[31];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[33];
  assign t[71] = t[88] ^ x[34];
  assign t[72] = t[89] ^ x[35];
  assign t[73] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[86] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[87] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[88] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[47] & t[13];
  assign t[90] = t[111] ^ x[8];
  assign t[91] = t[112] ^ x[33];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[9];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[15];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[16];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind87(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[20];
  assign t[105] = t[126] ^ x[14];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[31];
  assign t[112] = t[133] ^ x[25];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[121] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[122] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[123] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[126] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[127] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[128] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[129] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[132] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[133] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[50]);
  assign t[15] = ~(t[49] ^ t[14]);
  assign t[16] = t[51] ^ t[50];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[49] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[49] ^ t[27];
  assign t[23] = t[52] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[50] ^ t[53];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[54]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[52] ^ t[29]);
  assign t[31] = t[55] ^ t[54];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[52] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[52] ^ t[36];
  assign t[36] = t[54] ^ t[56];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[57]);
  assign t[42] = t[44] ^ t[9];
  assign t[43] = ~t[45];
  assign t[44] = t[16] ^ t[21];
  assign t[45] = ~(t[46]);
  assign t[46] = t[47] ^ t[24];
  assign t[47] = t[31] ^ t[34];
  assign t[48] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[49] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[60] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[60] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[51] = (t[60] & ~t[64]) | (~t[60] & t[64]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[60] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[60] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[54] = (t[66] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[66] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[55] = (t[66] & ~t[70]) | (~t[66] & t[70]);
  assign t[56] = (t[66] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[66] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[57] = (t[58] & ~t[73] & ~t[59]) | (~t[72] & t[73] & ~t[74]) | (~t[58] & ~t[73] & t[59]) | (t[72] & t[73] & t[74]);
  assign t[58] = t[75] ^ x[8];
  assign t[59] = t[76] ^ x[9];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[15];
  assign t[61] = t[78] ^ x[16];
  assign t[62] = t[79] ^ x[17];
  assign t[63] = t[80] ^ x[18];
  assign t[64] = t[81] ^ x[19];
  assign t[65] = t[82] ^ x[20];
  assign t[66] = t[83] ^ x[26];
  assign t[67] = t[84] ^ x[27];
  assign t[68] = t[85] ^ x[28];
  assign t[69] = t[86] ^ x[29];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[30];
  assign t[71] = t[88] ^ x[31];
  assign t[72] = t[89] ^ x[33];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[35];
  assign t[75] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[76] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[77] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[8] = t[49] & t[13];
  assign t[90] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[7];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind88(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[15];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[16];
  assign t[104] = t[125] ^ x[19];
  assign t[105] = t[126] ^ x[13];
  assign t[106] = t[127] ^ x[25];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[26];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[27];
  assign t[111] = t[132] ^ x[30];
  assign t[112] = t[133] ^ x[24];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[47] ^ t[15];
  assign t[120] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[121] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[122] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[123] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[124] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[125] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[126] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[127] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[128] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[129] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[131] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[132] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[133] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[48] ^ t[49];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[49]);
  assign t[16] = ~(t[47] ^ t[15]);
  assign t[17] = t[47] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[50] ^ t[30];
  assign t[26] = t[49] ^ t[51];
  assign t[27] = t[47] ^ t[13];
  assign t[28] = t[52] ^ t[53];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[50] ^ t[30]);
  assign t[32] = t[50] & t[34];
  assign t[33] = t[50] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[53] ^ t[54];
  assign t[36] = t[50] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[26] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[35] ^ t[23];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[60]) | (~t[58] & t[60]);
  assign t[49] = (t[58] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[60]) | (~t[58] & ~t[62] & t[63]) | (t[61] & t[62] & t[60]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[62] & ~t[60]) | (~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[62] & t[60]) | (t[61] & t[62] & t[63]);
  assign t[52] = (t[64] & ~t[66]) | (~t[64] & t[66]);
  assign t[53] = (t[64] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[66]) | (~t[64] & ~t[68] & t[69]) | (t[67] & t[68] & t[66]);
  assign t[54] = (t[64] & ~t[68] & ~t[66]) | (~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[68] & t[66]) | (t[67] & t[68] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[56] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = t[74] ^ x[7];
  assign t[57] = t[75] ^ x[8];
  assign t[58] = t[76] ^ x[14];
  assign t[59] = t[77] ^ x[15];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[16];
  assign t[61] = t[79] ^ x[17];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[19];
  assign t[64] = t[82] ^ x[25];
  assign t[65] = t[83] ^ x[26];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[29];
  assign t[69] = t[87] ^ x[30];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[32];
  assign t[71] = t[89] ^ x[33];
  assign t[72] = t[90] ^ x[34];
  assign t[73] = t[91] ^ x[35];
  assign t[74] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[83] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[89] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[7];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[8];
  assign t[95] = t[116] ^ x[33];
  assign t[96] = t[117] ^ x[34];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[6];
  assign t[99] = t[120] ^ x[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind89(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[19];
  assign t[103] = t[124] ^ x[13];
  assign t[104] = t[125] ^ x[25];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[30];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[24];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[119] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[11] = t[45] ^ t[15];
  assign t[120] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[121] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[122] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[123] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[126] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[127] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[128] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[129] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[46] ^ t[47];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[47]);
  assign t[16] = ~(t[45] ^ t[15]);
  assign t[17] = t[45] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[45] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[48] ^ t[30];
  assign t[26] = t[47] ^ t[49];
  assign t[27] = t[45] ^ t[13];
  assign t[28] = t[50] ^ t[51];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[51]);
  assign t[31] = ~(t[48] ^ t[30]);
  assign t[32] = t[48] & t[34];
  assign t[33] = t[48] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[51] ^ t[52];
  assign t[36] = t[48] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[5]);
  assign t[41] = ~(t[42] ^ t[53]);
  assign t[42] = ~t[43];
  assign t[43] = ~(t[18]);
  assign t[44] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[56] & ~t[58]) | (~t[56] & t[58]);
  assign t[47] = (t[56] & ~t[60] & ~t[61]) | (~t[59] & t[60] & ~t[58]) | (~t[56] & ~t[60] & t[61]) | (t[59] & t[60] & t[58]);
  assign t[48] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[49] = (t[56] & ~t[60] & ~t[58]) | (~t[59] & t[60] & ~t[61]) | (~t[56] & ~t[60] & t[58]) | (t[59] & t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[44]);
  assign t[50] = (t[62] & ~t[64]) | (~t[62] & t[64]);
  assign t[51] = (t[62] & ~t[66] & ~t[67]) | (~t[65] & t[66] & ~t[64]) | (~t[62] & ~t[66] & t[67]) | (t[65] & t[66] & t[64]);
  assign t[52] = (t[62] & ~t[66] & ~t[64]) | (~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[66] & t[64]) | (t[65] & t[66] & t[67]);
  assign t[53] = (t[54] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[54] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[54] = t[72] ^ x[7];
  assign t[55] = t[73] ^ x[8];
  assign t[56] = t[74] ^ x[14];
  assign t[57] = t[75] ^ x[15];
  assign t[58] = t[76] ^ x[16];
  assign t[59] = t[77] ^ x[17];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[25];
  assign t[63] = t[81] ^ x[26];
  assign t[64] = t[82] ^ x[27];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[29];
  assign t[67] = t[85] ^ x[30];
  assign t[68] = t[86] ^ x[32];
  assign t[69] = t[87] ^ x[33];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[34];
  assign t[71] = t[89] ^ x[35];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[81] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[86] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[87] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[88] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[111] ^ x[7];
  assign t[91] = t[112] ^ x[32];
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[6];
  assign t[97] = t[118] ^ x[14];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind90(x, y);
 input [35:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[101] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[102] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[103] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[104] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[105] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[35]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[114] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[115] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[116] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[118] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[119] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[11] = ~(t[37] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[38] ^ t[39];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = x[0] ? x[35] : t[18];
  assign t[18] = ~(t[19] ^ t[20]);
  assign t[19] = ~t[21];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[23] ^ t[41]);
  assign t[22] = t[24] ^ t[8];
  assign t[23] = ~t[25];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = ~(t[28]);
  assign t[26] = t[42] ^ t[35];
  assign t[27] = t[10] & t[29];
  assign t[28] = t[30] ^ t[14];
  assign t[29] = t[37] ^ t[7];
  assign t[2] = ~t[4];
  assign t[30] = t[31] ^ t[32];
  assign t[31] = t[43] ^ t[38];
  assign t[32] = t[15] & t[33];
  assign t[33] = t[40] ^ t[13];
  assign t[34] = (t[44] & ~t[46] & ~t[48]) | (~t[45] & t[46] & ~t[47]) | (~t[44] & ~t[46] & t[48]) | (t[45] & t[46] & t[47]);
  assign t[35] = (t[49] & ~t[51] & ~t[53]) | (~t[50] & t[51] & ~t[52]) | (~t[49] & ~t[51] & t[53]) | (t[50] & t[51] & t[52]);
  assign t[36] = (t[49] & ~t[51] & ~t[52]) | (~t[50] & t[51] & ~t[53]) | (~t[49] & ~t[51] & t[52]) | (t[50] & t[51] & t[53]);
  assign t[37] = (t[49] & ~t[54]) | (~t[49] & t[54]);
  assign t[38] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[39] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[60]) | (~t[55] & t[60]);
  assign t[41] = (t[44] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[44] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[42] = (t[49] & ~t[52]) | (~t[49] & t[52]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = t[61] ^ x[8];
  assign t[45] = t[62] ^ x[9];
  assign t[46] = t[63] ^ x[10];
  assign t[47] = t[64] ^ x[11];
  assign t[48] = t[65] ^ x[12];
  assign t[49] = t[66] ^ x[18];
  assign t[4] = ~(t[6] ^ t[34]);
  assign t[50] = t[67] ^ x[19];
  assign t[51] = t[68] ^ x[20];
  assign t[52] = t[69] ^ x[21];
  assign t[53] = t[70] ^ x[22];
  assign t[54] = t[71] ^ x[23];
  assign t[55] = t[72] ^ x[29];
  assign t[56] = t[73] ^ x[30];
  assign t[57] = t[74] ^ x[31];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[34];
  assign t[61] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[62] = (t[79] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (~t[78] & t[79] & ~t[81] & ~t[82] & ~t[84]) | (~t[78] & t[79] & ~t[80] & ~t[83] & ~t[84]) | (t[78] & ~t[79] & t[80] & t[81] & ~t[84]) | (t[78] & ~t[79] & t[82] & t[83] & ~t[84]) | (t[79] & ~t[81] & ~t[83] & t[84]) | (~t[79] & t[81] & t[83] & t[84]);
  assign t[63] = (t[78] & t[79] & t[80] & ~t[81] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & ~t[81] & ~t[82] & t[83] & t[84]) | (~t[79] & ~t[80] & t[81] & ~t[82] & ~t[83]) | (~t[78] & ~t[80] & t[81] & ~t[83] & ~t[84]) | (~t[78] & ~t[79] & t[81] & ~t[82] & ~t[84]) | (~t[79] & t[80] & t[81] & t[82] & ~t[83]) | (~t[80] & t[81] & t[82] & ~t[84]);
  assign t[64] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[65] = (t[78] & t[79] & ~t[81] & t[82] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & ~t[81] & ~t[82] & t[83]) | (~t[78] & ~t[81] & ~t[82] & t[83] & ~t[84]) | (~t[78] & ~t[79] & ~t[80] & t[83] & ~t[84]) | (~t[79] & t[80] & ~t[81] & t[82] & t[83]) | (t[80] & ~t[82] & t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = ~t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[72] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[73] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[74] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[8];
  assign t[79] = t[100] ^ x[9];
  assign t[7] = t[35] ^ t[36];
  assign t[80] = t[101] ^ x[6];
  assign t[81] = t[102] ^ x[10];
  assign t[82] = t[103] ^ x[11];
  assign t[83] = t[104] ^ x[12];
  assign t[84] = t[105] ^ x[7];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[23];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[29];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[32];
  assign t[97] = t[118] ^ x[33];
  assign t[98] = t[119] ^ x[28];
  assign t[99] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~t[17]) | (~t[0] & t[17]);
endmodule

module R2ind91(x, y);
 input [36:0] x;
 output y;

 wire [150:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & t[124] & ~t[125] & t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[125] & ~t[126] & t[127] & ~t[128] & t[129]) | (~t[124] & t[125] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[124] & t[125] & ~t[128] & ~t[129]) | (~t[123] & t[125] & t[126] & ~t[127] & t[128]) | (t[125] & ~t[126] & t[128] & ~t[129]);
  assign t[101] = (t[124] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & t[124] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[124] & ~t[125] & ~t[128] & ~t[129]) | (t[123] & ~t[124] & t[125] & t[126] & ~t[129]) | (t[123] & ~t[124] & t[127] & t[128] & ~t[129]) | (t[124] & ~t[126] & ~t[128] & t[129]) | (~t[124] & t[126] & t[128] & t[129]);
  assign t[102] = (t[123] & t[124] & t[125] & ~t[126] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[126] & ~t[127] & t[128] & t[129]) | (~t[124] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[125] & t[126] & ~t[128] & ~t[129]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[129]) | (~t[124] & t[125] & t[126] & t[127] & ~t[128]) | (~t[125] & t[126] & t[127] & ~t[129]);
  assign t[103] = (t[123] & t[124] & ~t[125] & ~t[127] & t[128] & ~t[129]) | (t[123] & t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[129]) | (~t[123] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[123] & ~t[124] & ~t[126] & t[127] & ~t[129]) | (~t[123] & ~t[125] & t[126] & t[127] & t[128]) | (t[126] & t[127] & ~t[128] & ~t[129]);
  assign t[104] = (t[123] & t[124] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[123] & ~t[124] & ~t[125] & t[128] & ~t[129]) | (~t[124] & t[125] & ~t[126] & t[127] & t[128]) | (t[125] & ~t[127] & t[128] & ~t[129]);
  assign t[105] = (t[109] & t[110] & ~t[111] & t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[111] & ~t[112] & t[113] & ~t[114] & t[115]) | (~t[110] & t[111] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[110] & t[111] & ~t[114] & ~t[115]) | (~t[109] & t[111] & t[112] & ~t[113] & t[114]) | (t[111] & ~t[112] & t[114] & ~t[115]);
  assign t[106] = (t[110] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (~t[109] & t[110] & ~t[112] & ~t[113] & ~t[115]) | (~t[109] & t[110] & ~t[111] & ~t[114] & ~t[115]) | (t[109] & ~t[110] & t[111] & t[112] & ~t[115]) | (t[109] & ~t[110] & t[113] & t[114] & ~t[115]) | (t[110] & ~t[112] & ~t[114] & t[115]) | (~t[110] & t[112] & t[114] & t[115]);
  assign t[107] = (t[109] & t[110] & t[111] & ~t[112] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & ~t[112] & ~t[113] & t[114] & t[115]) | (~t[110] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (~t[109] & ~t[111] & t[112] & ~t[114] & ~t[115]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[115]) | (~t[110] & t[111] & t[112] & t[113] & ~t[114]) | (~t[111] & t[112] & t[113] & ~t[115]);
  assign t[108] = (t[109] & t[110] & ~t[112] & t[113] & ~t[114] & ~t[115]) | (t[110] & ~t[111] & t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[112] & ~t[113] & t[114] & ~t[115]) | (~t[109] & ~t[110] & ~t[111] & t[114] & ~t[115]) | (~t[110] & t[111] & ~t[112] & t[113] & t[114]) | (t[111] & ~t[113] & t[114] & ~t[115]);
  assign t[109] = t[130] ^ x[7];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[34];
  assign t[111] = t[132] ^ x[32];
  assign t[112] = t[133] ^ x[35];
  assign t[113] = t[134] ^ x[8];
  assign t[114] = t[135] ^ x[36];
  assign t[115] = t[136] ^ x[6];
  assign t[116] = t[137] ^ x[14];
  assign t[117] = t[138] ^ x[16];
  assign t[118] = t[139] ^ x[15];
  assign t[119] = t[140] ^ x[17];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[18];
  assign t[121] = t[142] ^ x[19];
  assign t[122] = t[143] ^ x[13];
  assign t[123] = t[144] ^ x[25];
  assign t[124] = t[145] ^ x[27];
  assign t[125] = t[146] ^ x[26];
  assign t[126] = t[147] ^ x[28];
  assign t[127] = t[148] ^ x[29];
  assign t[128] = t[149] ^ x[30];
  assign t[129] = t[150] ^ x[24];
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[131] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[132] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[133] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[134] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[135] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[136] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[137] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[138] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[139] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[141] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[142] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[143] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[144] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[145] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[146] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[147] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[148] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[149] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[14] = ~(t[64]);
  assign t[150] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[15] = ~(t[63] ^ t[14]);
  assign t[16] = t[65] ^ t[64];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[63] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[63] ^ t[27];
  assign t[23] = t[66] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[64] ^ t[67];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[68]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[66] ^ t[29]);
  assign t[31] = t[69] ^ t[68];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[66] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[66] ^ t[36];
  assign t[36] = t[68] ^ t[70];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[71]);
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~t[46];
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~(t[49] ^ t[50]);
  assign t[47] = t[16] ^ t[21];
  assign t[48] = t[63] ^ t[14];
  assign t[49] = t[51] ^ t[24];
  assign t[4] = ~(t[7] ^ t[62]);
  assign t[50] = t[18] ^ t[52];
  assign t[51] = t[31] ^ t[34];
  assign t[52] = t[66] ^ t[29];
  assign t[53] = x[0] ? x[33] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~t[57];
  assign t[56] = ~(t[58]);
  assign t[57] = ~(t[59] ^ t[72]);
  assign t[58] = t[27] ^ t[9];
  assign t[59] = ~t[60];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[61]);
  assign t[61] = t[36] ^ t[24];
  assign t[62] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[63] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[64] = (t[75] & ~t[78] & ~t[80]) | (~t[77] & t[78] & ~t[79]) | (~t[75] & ~t[78] & t[80]) | (t[77] & t[78] & t[79]);
  assign t[65] = (t[75] & ~t[79]) | (~t[75] & t[79]);
  assign t[66] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[67] = (t[75] & ~t[78] & ~t[79]) | (~t[77] & t[78] & ~t[80]) | (~t[75] & ~t[78] & t[79]) | (t[77] & t[78] & t[80]);
  assign t[68] = (t[81] & ~t[84] & ~t[86]) | (~t[83] & t[84] & ~t[85]) | (~t[81] & ~t[84] & t[86]) | (t[83] & t[84] & t[85]);
  assign t[69] = (t[81] & ~t[85]) | (~t[81] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[81] & ~t[84] & ~t[85]) | (~t[83] & t[84] & ~t[86]) | (~t[81] & ~t[84] & t[85]) | (t[83] & t[84] & t[86]);
  assign t[71] = (t[73] & ~t[87]) | (~t[73] & t[87]);
  assign t[72] = (t[73] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[74]) | (~t[73] & ~t[89] & t[90]) | (t[88] & t[89] & t[74]);
  assign t[73] = t[91] ^ x[7];
  assign t[74] = t[92] ^ x[8];
  assign t[75] = t[93] ^ x[14];
  assign t[76] = t[94] ^ x[15];
  assign t[77] = t[95] ^ x[16];
  assign t[78] = t[96] ^ x[17];
  assign t[79] = t[97] ^ x[18];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[19];
  assign t[81] = t[99] ^ x[25];
  assign t[82] = t[100] ^ x[26];
  assign t[83] = t[101] ^ x[27];
  assign t[84] = t[102] ^ x[28];
  assign t[85] = t[103] ^ x[29];
  assign t[86] = t[104] ^ x[30];
  assign t[87] = t[105] ^ x[32];
  assign t[88] = t[106] ^ x[34];
  assign t[89] = t[107] ^ x[35];
  assign t[8] = t[63] & t[13];
  assign t[90] = t[108] ^ x[36];
  assign t[91] = (t[109] & ~t[111] & ~t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[112] & ~t[113] & ~t[115]) | (t[109] & ~t[110] & ~t[111] & ~t[114] & ~t[115]) | (~t[109] & t[110] & t[111] & t[112] & ~t[115]) | (~t[109] & t[110] & t[113] & t[114] & ~t[115]) | (t[109] & ~t[111] & ~t[113] & t[115]) | (~t[109] & t[111] & t[113] & t[115]);
  assign t[92] = (t[109] & t[110] & ~t[111] & ~t[113] & t[114] & ~t[115]) | (t[109] & t[111] & ~t[112] & ~t[113] & ~t[114] & t[115]) | (~t[110] & ~t[111] & t[113] & ~t[114] & ~t[115]) | (~t[109] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[109] & ~t[110] & ~t[112] & t[113] & ~t[115]) | (~t[109] & ~t[111] & t[112] & t[113] & t[114]) | (t[112] & t[113] & ~t[114] & ~t[115]);
  assign t[93] = (t[116] & ~t[118] & ~t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[119] & ~t[120] & ~t[122]) | (t[116] & ~t[117] & ~t[118] & ~t[121] & ~t[122]) | (~t[116] & t[117] & t[118] & t[119] & ~t[122]) | (~t[116] & t[117] & t[120] & t[121] & ~t[122]) | (t[116] & ~t[118] & ~t[120] & t[122]) | (~t[116] & t[118] & t[120] & t[122]);
  assign t[94] = (t[116] & t[117] & ~t[118] & t[119] & ~t[120] & ~t[122]) | (t[116] & ~t[118] & ~t[119] & t[120] & ~t[121] & t[122]) | (~t[117] & t[118] & ~t[119] & ~t[120] & ~t[122]) | (~t[116] & t[118] & ~t[119] & ~t[120] & ~t[121]) | (~t[116] & ~t[117] & t[118] & ~t[121] & ~t[122]) | (~t[116] & t[118] & t[119] & ~t[120] & t[121]) | (t[118] & ~t[119] & t[121] & ~t[122]);
  assign t[95] = (t[117] & ~t[118] & ~t[119] & ~t[120] & ~t[121]) | (~t[116] & t[117] & ~t[119] & ~t[120] & ~t[122]) | (~t[116] & t[117] & ~t[118] & ~t[121] & ~t[122]) | (t[116] & ~t[117] & t[118] & t[119] & ~t[122]) | (t[116] & ~t[117] & t[120] & t[121] & ~t[122]) | (t[117] & ~t[119] & ~t[121] & t[122]) | (~t[117] & t[119] & t[121] & t[122]);
  assign t[96] = (t[116] & t[117] & t[118] & ~t[119] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & ~t[119] & ~t[120] & t[121] & t[122]) | (~t[117] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (~t[116] & ~t[118] & t[119] & ~t[121] & ~t[122]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[122]) | (~t[117] & t[118] & t[119] & t[120] & ~t[121]) | (~t[118] & t[119] & t[120] & ~t[122]);
  assign t[97] = (t[116] & t[117] & ~t[118] & ~t[120] & t[121] & ~t[122]) | (t[116] & t[118] & ~t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[118] & t[120] & ~t[121] & ~t[122]) | (~t[116] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[116] & ~t[117] & ~t[119] & t[120] & ~t[122]) | (~t[116] & ~t[118] & t[119] & t[120] & t[121]) | (t[119] & t[120] & ~t[121] & ~t[122]);
  assign t[98] = (t[116] & t[117] & ~t[119] & t[120] & ~t[121] & ~t[122]) | (t[117] & ~t[118] & t[119] & ~t[120] & ~t[121] & t[122]) | (~t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[119] & ~t[120] & t[121] & ~t[122]) | (~t[116] & ~t[117] & ~t[118] & t[121] & ~t[122]) | (~t[117] & t[118] & ~t[119] & t[120] & t[121]) | (t[118] & ~t[120] & t[121] & ~t[122]);
  assign t[99] = (t[123] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[124] & ~t[125] & ~t[128] & ~t[129]) | (~t[123] & t[124] & t[125] & t[126] & ~t[129]) | (~t[123] & t[124] & t[127] & t[128] & ~t[129]) | (t[123] & ~t[125] & ~t[127] & t[129]) | (~t[123] & t[125] & t[127] & t[129]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[53]) | (~t[0] & t[37] & ~t[53]) | (~t[0] & ~t[37] & t[53]) | (t[0] & t[37] & t[53]);
endmodule

module R2ind92(x, y);
 input [36:0] x;
 output y;

 wire [148:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[121] & t[122] & t[123] & ~t[124] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[124] & ~t[125] & t[126] & t[127]) | (~t[122] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[123] & t[124] & ~t[126] & ~t[127]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[127]) | (~t[122] & t[123] & t[124] & t[125] & ~t[126]) | (~t[123] & t[124] & t[125] & ~t[127]);
  assign t[101] = (t[121] & t[122] & ~t[123] & ~t[125] & t[126] & ~t[127]) | (t[121] & t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[127]) | (~t[121] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[121] & ~t[122] & ~t[124] & t[125] & ~t[127]) | (~t[121] & ~t[123] & t[124] & t[125] & t[126]) | (t[124] & t[125] & ~t[126] & ~t[127]);
  assign t[102] = (t[121] & t[122] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[121] & ~t[122] & ~t[123] & t[126] & ~t[127]) | (~t[122] & t[123] & ~t[124] & t[125] & t[126]) | (t[123] & ~t[125] & t[126] & ~t[127]);
  assign t[103] = (t[107] & t[108] & ~t[109] & t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[109] & ~t[110] & t[111] & ~t[112] & t[113]) | (~t[108] & t[109] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[108] & t[109] & ~t[112] & ~t[113]) | (~t[107] & t[109] & t[110] & ~t[111] & t[112]) | (t[109] & ~t[110] & t[112] & ~t[113]);
  assign t[104] = (t[108] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & t[108] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[108] & ~t[109] & ~t[112] & ~t[113]) | (t[107] & ~t[108] & t[109] & t[110] & ~t[113]) | (t[107] & ~t[108] & t[111] & t[112] & ~t[113]) | (t[108] & ~t[110] & ~t[112] & t[113]) | (~t[108] & t[110] & t[112] & t[113]);
  assign t[105] = (t[107] & t[108] & t[109] & ~t[110] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[110] & ~t[111] & t[112] & t[113]) | (~t[108] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[109] & t[110] & ~t[112] & ~t[113]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[113]) | (~t[108] & t[109] & t[110] & t[111] & ~t[112]) | (~t[109] & t[110] & t[111] & ~t[113]);
  assign t[106] = (t[107] & t[108] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[107] & ~t[108] & ~t[109] & t[112] & ~t[113]) | (~t[108] & t[109] & ~t[110] & t[111] & t[112]) | (t[109] & ~t[111] & t[112] & ~t[113]);
  assign t[107] = t[128] ^ x[7];
  assign t[108] = t[129] ^ x[34];
  assign t[109] = t[130] ^ x[32];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[35];
  assign t[111] = t[132] ^ x[8];
  assign t[112] = t[133] ^ x[36];
  assign t[113] = t[134] ^ x[6];
  assign t[114] = t[135] ^ x[14];
  assign t[115] = t[136] ^ x[16];
  assign t[116] = t[137] ^ x[15];
  assign t[117] = t[138] ^ x[17];
  assign t[118] = t[139] ^ x[18];
  assign t[119] = t[140] ^ x[19];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[13];
  assign t[121] = t[142] ^ x[25];
  assign t[122] = t[143] ^ x[27];
  assign t[123] = t[144] ^ x[26];
  assign t[124] = t[145] ^ x[28];
  assign t[125] = t[146] ^ x[29];
  assign t[126] = t[147] ^ x[30];
  assign t[127] = t[148] ^ x[24];
  assign t[128] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[129] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[131] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[132] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[133] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[134] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[135] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[136] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[137] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[138] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[139] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[141] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[142] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[143] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[144] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[145] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[146] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[147] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[148] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[62]);
  assign t[15] = ~(t[61] ^ t[14]);
  assign t[16] = t[63] ^ t[62];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[61] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[61] ^ t[27];
  assign t[23] = t[64] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[62] ^ t[65];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[66]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[64] ^ t[29]);
  assign t[31] = t[67] ^ t[66];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[64] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[64] ^ t[36];
  assign t[36] = t[66] ^ t[68];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[69]);
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~t[46];
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~(t[49] ^ t[50]);
  assign t[47] = t[16] ^ t[21];
  assign t[48] = t[61] ^ t[14];
  assign t[49] = t[51] ^ t[24];
  assign t[4] = ~(t[7] ^ t[60]);
  assign t[50] = t[18] ^ t[52];
  assign t[51] = t[31] ^ t[34];
  assign t[52] = t[64] ^ t[29];
  assign t[53] = x[0] ? x[33] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~t[57];
  assign t[56] = ~(t[44]);
  assign t[57] = ~(t[58] ^ t[70]);
  assign t[58] = ~t[59];
  assign t[59] = ~(t[49]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[61] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[62] = (t[73] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[73] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[63] = (t[73] & ~t[77]) | (~t[73] & t[77]);
  assign t[64] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[65] = (t[73] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[73] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[66] = (t[79] & ~t[82] & ~t[84]) | (~t[81] & t[82] & ~t[83]) | (~t[79] & ~t[82] & t[84]) | (t[81] & t[82] & t[83]);
  assign t[67] = (t[79] & ~t[83]) | (~t[79] & t[83]);
  assign t[68] = (t[79] & ~t[82] & ~t[83]) | (~t[81] & t[82] & ~t[84]) | (~t[79] & ~t[82] & t[83]) | (t[81] & t[82] & t[84]);
  assign t[69] = (t[71] & ~t[85]) | (~t[71] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[71] & ~t[87] & ~t[72]) | (~t[86] & t[87] & ~t[88]) | (~t[71] & ~t[87] & t[72]) | (t[86] & t[87] & t[88]);
  assign t[71] = t[89] ^ x[7];
  assign t[72] = t[90] ^ x[8];
  assign t[73] = t[91] ^ x[14];
  assign t[74] = t[92] ^ x[15];
  assign t[75] = t[93] ^ x[16];
  assign t[76] = t[94] ^ x[17];
  assign t[77] = t[95] ^ x[18];
  assign t[78] = t[96] ^ x[19];
  assign t[79] = t[97] ^ x[25];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[26];
  assign t[81] = t[99] ^ x[27];
  assign t[82] = t[100] ^ x[28];
  assign t[83] = t[101] ^ x[29];
  assign t[84] = t[102] ^ x[30];
  assign t[85] = t[103] ^ x[32];
  assign t[86] = t[104] ^ x[34];
  assign t[87] = t[105] ^ x[35];
  assign t[88] = t[106] ^ x[36];
  assign t[89] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[8] = t[61] & t[13];
  assign t[90] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[91] = (t[114] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[115] & ~t[116] & ~t[119] & ~t[120]) | (~t[114] & t[115] & t[116] & t[117] & ~t[120]) | (~t[114] & t[115] & t[118] & t[119] & ~t[120]) | (t[114] & ~t[116] & ~t[118] & t[120]) | (~t[114] & t[116] & t[118] & t[120]);
  assign t[92] = (t[114] & t[115] & ~t[116] & t[117] & ~t[118] & ~t[120]) | (t[114] & ~t[116] & ~t[117] & t[118] & ~t[119] & t[120]) | (~t[115] & t[116] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[115] & t[116] & ~t[119] & ~t[120]) | (~t[114] & t[116] & t[117] & ~t[118] & t[119]) | (t[116] & ~t[117] & t[119] & ~t[120]);
  assign t[93] = (t[115] & ~t[116] & ~t[117] & ~t[118] & ~t[119]) | (~t[114] & t[115] & ~t[117] & ~t[118] & ~t[120]) | (~t[114] & t[115] & ~t[116] & ~t[119] & ~t[120]) | (t[114] & ~t[115] & t[116] & t[117] & ~t[120]) | (t[114] & ~t[115] & t[118] & t[119] & ~t[120]) | (t[115] & ~t[117] & ~t[119] & t[120]) | (~t[115] & t[117] & t[119] & t[120]);
  assign t[94] = (t[114] & t[115] & t[116] & ~t[117] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[117] & ~t[118] & t[119] & t[120]) | (~t[115] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (~t[114] & ~t[116] & t[117] & ~t[119] & ~t[120]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[120]) | (~t[115] & t[116] & t[117] & t[118] & ~t[119]) | (~t[116] & t[117] & t[118] & ~t[120]);
  assign t[95] = (t[114] & t[115] & ~t[116] & ~t[118] & t[119] & ~t[120]) | (t[114] & t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[120]) | (~t[114] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[114] & ~t[115] & ~t[117] & t[118] & ~t[120]) | (~t[114] & ~t[116] & t[117] & t[118] & t[119]) | (t[117] & t[118] & ~t[119] & ~t[120]);
  assign t[96] = (t[114] & t[115] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[114] & ~t[115] & ~t[116] & t[119] & ~t[120]) | (~t[115] & t[116] & ~t[117] & t[118] & t[119]) | (t[116] & ~t[118] & t[119] & ~t[120]);
  assign t[97] = (t[121] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[122] & ~t[123] & ~t[126] & ~t[127]) | (~t[121] & t[122] & t[123] & t[124] & ~t[127]) | (~t[121] & t[122] & t[125] & t[126] & ~t[127]) | (t[121] & ~t[123] & ~t[125] & t[127]) | (~t[121] & t[123] & t[125] & t[127]);
  assign t[98] = (t[121] & t[122] & ~t[123] & t[124] & ~t[125] & ~t[127]) | (t[121] & ~t[123] & ~t[124] & t[125] & ~t[126] & t[127]) | (~t[122] & t[123] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & ~t[122] & t[123] & ~t[126] & ~t[127]) | (~t[121] & t[123] & t[124] & ~t[125] & t[126]) | (t[123] & ~t[124] & t[126] & ~t[127]);
  assign t[99] = (t[122] & ~t[123] & ~t[124] & ~t[125] & ~t[126]) | (~t[121] & t[122] & ~t[124] & ~t[125] & ~t[127]) | (~t[121] & t[122] & ~t[123] & ~t[126] & ~t[127]) | (t[121] & ~t[122] & t[123] & t[124] & ~t[127]) | (t[121] & ~t[122] & t[125] & t[126] & ~t[127]) | (t[122] & ~t[124] & ~t[126] & t[127]) | (~t[122] & t[124] & t[126] & t[127]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[53]) | (~t[0] & t[37] & ~t[53]) | (~t[0] & ~t[37] & t[53]) | (t[0] & t[37] & t[53]);
endmodule

module R2ind93(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[19];
  assign t[102] = t[123] ^ x[20];
  assign t[103] = t[124] ^ x[14];
  assign t[104] = t[125] ^ x[26];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[27];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[30];
  assign t[109] = t[130] ^ x[31];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[25];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[119] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[121] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[122] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[123] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[124] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[125] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[126] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[127] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[128] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[129] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[131] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[48]);
  assign t[15] = ~(t[47] ^ t[14]);
  assign t[16] = t[49] ^ t[48];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[47] ^ t[27];
  assign t[23] = t[50] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[48] ^ t[51];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[52]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[50] ^ t[29]);
  assign t[31] = t[53] ^ t[52];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[50] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[50] ^ t[36];
  assign t[36] = t[52] ^ t[54];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[27] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[36] ^ t[24];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[58] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[49] = (t[58] & ~t[62]) | (~t[58] & t[62]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[58] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[52] = (t[64] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[64] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[64] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[57]) | (~t[56] & ~t[71] & t[72]) | (t[70] & t[71] & t[57]);
  assign t[56] = t[73] ^ x[8];
  assign t[57] = t[74] ^ x[9];
  assign t[58] = t[75] ^ x[15];
  assign t[59] = t[76] ^ x[16];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[17];
  assign t[61] = t[78] ^ x[18];
  assign t[62] = t[79] ^ x[19];
  assign t[63] = t[80] ^ x[20];
  assign t[64] = t[81] ^ x[26];
  assign t[65] = t[82] ^ x[27];
  assign t[66] = t[83] ^ x[28];
  assign t[67] = t[84] ^ x[29];
  assign t[68] = t[85] ^ x[30];
  assign t[69] = t[86] ^ x[31];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[33];
  assign t[71] = t[88] ^ x[34];
  assign t[72] = t[89] ^ x[35];
  assign t[73] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[86] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[87] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[88] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[47] & t[13];
  assign t[90] = t[111] ^ x[8];
  assign t[91] = t[112] ^ x[33];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[9];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[15];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[16];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind94(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[20];
  assign t[105] = t[126] ^ x[14];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[31];
  assign t[112] = t[133] ^ x[25];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[121] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[122] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[123] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[126] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[127] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[128] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[129] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[132] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[133] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[50]);
  assign t[15] = ~(t[49] ^ t[14]);
  assign t[16] = t[51] ^ t[50];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[49] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[49] ^ t[27];
  assign t[23] = t[52] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[50] ^ t[53];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[54]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[52] ^ t[29]);
  assign t[31] = t[55] ^ t[54];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[52] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[52] ^ t[36];
  assign t[36] = t[54] ^ t[56];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[57]);
  assign t[42] = t[44] ^ t[9];
  assign t[43] = ~t[45];
  assign t[44] = t[16] ^ t[21];
  assign t[45] = ~(t[46]);
  assign t[46] = t[47] ^ t[24];
  assign t[47] = t[31] ^ t[34];
  assign t[48] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[49] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[60] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[60] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[51] = (t[60] & ~t[64]) | (~t[60] & t[64]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[60] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[60] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[54] = (t[66] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[66] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[55] = (t[66] & ~t[70]) | (~t[66] & t[70]);
  assign t[56] = (t[66] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[66] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[57] = (t[58] & ~t[73] & ~t[59]) | (~t[72] & t[73] & ~t[74]) | (~t[58] & ~t[73] & t[59]) | (t[72] & t[73] & t[74]);
  assign t[58] = t[75] ^ x[8];
  assign t[59] = t[76] ^ x[9];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[15];
  assign t[61] = t[78] ^ x[16];
  assign t[62] = t[79] ^ x[17];
  assign t[63] = t[80] ^ x[18];
  assign t[64] = t[81] ^ x[19];
  assign t[65] = t[82] ^ x[20];
  assign t[66] = t[83] ^ x[26];
  assign t[67] = t[84] ^ x[27];
  assign t[68] = t[85] ^ x[28];
  assign t[69] = t[86] ^ x[29];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[30];
  assign t[71] = t[88] ^ x[31];
  assign t[72] = t[89] ^ x[33];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[35];
  assign t[75] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[76] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[77] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[8] = t[49] & t[13];
  assign t[90] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[7];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind95(x, y);
 input [35:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[14];
  assign t[101] = t[122] ^ x[17];
  assign t[102] = t[123] ^ x[15];
  assign t[103] = t[124] ^ x[18];
  assign t[104] = t[125] ^ x[16];
  assign t[105] = t[126] ^ x[19];
  assign t[106] = t[127] ^ x[13];
  assign t[107] = t[128] ^ x[25];
  assign t[108] = t[129] ^ x[28];
  assign t[109] = t[130] ^ x[26];
  assign t[10] = t[16] ^ t[17];
  assign t[110] = t[131] ^ x[29];
  assign t[111] = t[132] ^ x[27];
  assign t[112] = t[133] ^ x[30];
  assign t[113] = t[134] ^ x[24];
  assign t[114] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[115] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[116] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[117] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[118] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[119] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[121] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[122] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[123] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[124] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[125] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[126] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[127] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[128] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[129] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[131] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[132] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[133] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[134] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[48] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[49] ^ t[50];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[50]);
  assign t[19] = ~(t[48] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[48] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[51] ^ t[29];
  assign t[25] = t[48] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[52] ^ t[53];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[53]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[51] ^ t[29]);
  assign t[31] = t[51] & t[35];
  assign t[32] = t[50] ^ t[54];
  assign t[33] = t[48] ^ t[16];
  assign t[34] = t[51] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[53] ^ t[55];
  assign t[37] = t[51] ^ t[27];
  assign t[38] = x[0] ? x[31] : t[39];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5]);
  assign t[40] = ~t[42];
  assign t[41] = ~(t[43]);
  assign t[42] = ~(t[44] ^ t[56]);
  assign t[43] = t[32] ^ t[11];
  assign t[44] = ~t[45];
  assign t[45] = ~(t[46]);
  assign t[46] = t[36] ^ t[22];
  assign t[47] = (t[57] & ~t[58]) | (~t[57] & t[58]);
  assign t[48] = (t[59] & ~t[60]) | (~t[59] & t[60]);
  assign t[49] = (t[59] & ~t[61]) | (~t[59] & t[61]);
  assign t[4] = ~(t[6] ^ t[47]);
  assign t[50] = (t[59] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[61]) | (~t[59] & ~t[63] & t[64]) | (t[62] & t[63] & t[61]);
  assign t[51] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[52] = (t[65] & ~t[67]) | (~t[65] & t[67]);
  assign t[53] = (t[65] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[67]) | (~t[65] & ~t[69] & t[70]) | (t[68] & t[69] & t[67]);
  assign t[54] = (t[59] & ~t[63] & ~t[61]) | (~t[62] & t[63] & ~t[64]) | (~t[59] & ~t[63] & t[61]) | (t[62] & t[63] & t[64]);
  assign t[55] = (t[65] & ~t[69] & ~t[67]) | (~t[68] & t[69] & ~t[70]) | (~t[65] & ~t[69] & t[67]) | (t[68] & t[69] & t[70]);
  assign t[56] = (t[57] & ~t[72] & ~t[74]) | (~t[71] & t[72] & ~t[73]) | (~t[57] & ~t[72] & t[74]) | (t[71] & t[72] & t[73]);
  assign t[57] = t[75] ^ x[7];
  assign t[58] = t[76] ^ x[8];
  assign t[59] = t[77] ^ x[14];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = t[78] ^ x[15];
  assign t[61] = t[79] ^ x[16];
  assign t[62] = t[80] ^ x[17];
  assign t[63] = t[81] ^ x[18];
  assign t[64] = t[82] ^ x[19];
  assign t[65] = t[83] ^ x[25];
  assign t[66] = t[84] ^ x[26];
  assign t[67] = t[85] ^ x[27];
  assign t[68] = t[86] ^ x[28];
  assign t[69] = t[87] ^ x[29];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[30];
  assign t[71] = t[89] ^ x[32];
  assign t[72] = t[90] ^ x[33];
  assign t[73] = t[91] ^ x[34];
  assign t[74] = t[92] ^ x[35];
  assign t[75] = (t[93] & ~t[95] & ~t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[96] & ~t[97] & ~t[99]) | (t[93] & ~t[94] & ~t[95] & ~t[98] & ~t[99]) | (~t[93] & t[94] & t[95] & t[96] & ~t[99]) | (~t[93] & t[94] & t[97] & t[98] & ~t[99]) | (t[93] & ~t[95] & ~t[97] & t[99]) | (~t[93] & t[95] & t[97] & t[99]);
  assign t[76] = (t[93] & t[94] & ~t[95] & t[96] & ~t[97] & ~t[99]) | (t[93] & ~t[95] & ~t[96] & t[97] & ~t[98] & t[99]) | (~t[94] & t[95] & ~t[96] & ~t[97] & ~t[99]) | (~t[93] & t[95] & ~t[96] & ~t[97] & ~t[98]) | (~t[93] & ~t[94] & t[95] & ~t[98] & ~t[99]) | (~t[93] & t[95] & t[96] & ~t[97] & t[98]) | (t[95] & ~t[96] & t[98] & ~t[99]);
  assign t[77] = (t[100] & ~t[102] & ~t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[103] & ~t[104] & ~t[106]) | (t[100] & ~t[101] & ~t[102] & ~t[105] & ~t[106]) | (~t[100] & t[101] & t[102] & t[103] & ~t[106]) | (~t[100] & t[101] & t[104] & t[105] & ~t[106]) | (t[100] & ~t[102] & ~t[104] & t[106]) | (~t[100] & t[102] & t[104] & t[106]);
  assign t[78] = (t[100] & t[101] & ~t[102] & t[103] & ~t[104] & ~t[106]) | (t[100] & ~t[102] & ~t[103] & t[104] & ~t[105] & t[106]) | (~t[101] & t[102] & ~t[103] & ~t[104] & ~t[106]) | (~t[100] & t[102] & ~t[103] & ~t[104] & ~t[105]) | (~t[100] & ~t[101] & t[102] & ~t[105] & ~t[106]) | (~t[100] & t[102] & t[103] & ~t[104] & t[105]) | (t[102] & ~t[103] & t[105] & ~t[106]);
  assign t[79] = (t[100] & t[101] & ~t[102] & ~t[104] & t[105] & ~t[106]) | (t[100] & t[102] & ~t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[102] & t[104] & ~t[105] & ~t[106]) | (~t[100] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[100] & ~t[101] & ~t[103] & t[104] & ~t[106]) | (~t[100] & ~t[102] & t[103] & t[104] & t[105]) | (t[103] & t[104] & ~t[105] & ~t[106]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (t[101] & ~t[102] & ~t[103] & ~t[104] & ~t[105]) | (~t[100] & t[101] & ~t[103] & ~t[104] & ~t[106]) | (~t[100] & t[101] & ~t[102] & ~t[105] & ~t[106]) | (t[100] & ~t[101] & t[102] & t[103] & ~t[106]) | (t[100] & ~t[101] & t[104] & t[105] & ~t[106]) | (t[101] & ~t[103] & ~t[105] & t[106]) | (~t[101] & t[103] & t[105] & t[106]);
  assign t[81] = (t[100] & t[101] & t[102] & ~t[103] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & ~t[103] & ~t[104] & t[105] & t[106]) | (~t[101] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (~t[100] & ~t[102] & t[103] & ~t[105] & ~t[106]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[106]) | (~t[101] & t[102] & t[103] & t[104] & ~t[105]) | (~t[102] & t[103] & t[104] & ~t[106]);
  assign t[82] = (t[100] & t[101] & ~t[103] & t[104] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[103] & ~t[104] & t[105] & ~t[106]) | (~t[100] & ~t[101] & ~t[102] & t[105] & ~t[106]) | (~t[101] & t[102] & ~t[103] & t[104] & t[105]) | (t[102] & ~t[104] & t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[108] & ~t[109] & ~t[112] & ~t[113]) | (~t[107] & t[108] & t[109] & t[110] & ~t[113]) | (~t[107] & t[108] & t[111] & t[112] & ~t[113]) | (t[107] & ~t[109] & ~t[111] & t[113]) | (~t[107] & t[109] & t[111] & t[113]);
  assign t[84] = (t[107] & t[108] & ~t[109] & t[110] & ~t[111] & ~t[113]) | (t[107] & ~t[109] & ~t[110] & t[111] & ~t[112] & t[113]) | (~t[108] & t[109] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[108] & t[109] & ~t[112] & ~t[113]) | (~t[107] & t[109] & t[110] & ~t[111] & t[112]) | (t[109] & ~t[110] & t[112] & ~t[113]);
  assign t[85] = (t[107] & t[108] & ~t[109] & ~t[111] & t[112] & ~t[113]) | (t[107] & t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[113]) | (~t[107] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[107] & ~t[108] & ~t[110] & t[111] & ~t[113]) | (~t[107] & ~t[109] & t[110] & t[111] & t[112]) | (t[110] & t[111] & ~t[112] & ~t[113]);
  assign t[86] = (t[108] & ~t[109] & ~t[110] & ~t[111] & ~t[112]) | (~t[107] & t[108] & ~t[110] & ~t[111] & ~t[113]) | (~t[107] & t[108] & ~t[109] & ~t[112] & ~t[113]) | (t[107] & ~t[108] & t[109] & t[110] & ~t[113]) | (t[107] & ~t[108] & t[111] & t[112] & ~t[113]) | (t[108] & ~t[110] & ~t[112] & t[113]) | (~t[108] & t[110] & t[112] & t[113]);
  assign t[87] = (t[107] & t[108] & t[109] & ~t[110] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[110] & ~t[111] & t[112] & t[113]) | (~t[108] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (~t[107] & ~t[109] & t[110] & ~t[112] & ~t[113]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[113]) | (~t[108] & t[109] & t[110] & t[111] & ~t[112]) | (~t[109] & t[110] & t[111] & ~t[113]);
  assign t[88] = (t[107] & t[108] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[107] & ~t[108] & ~t[109] & t[112] & ~t[113]) | (~t[108] & t[109] & ~t[110] & t[111] & t[112]) | (t[109] & ~t[111] & t[112] & ~t[113]);
  assign t[89] = (t[94] & ~t[95] & ~t[96] & ~t[97] & ~t[98]) | (~t[93] & t[94] & ~t[96] & ~t[97] & ~t[99]) | (~t[93] & t[94] & ~t[95] & ~t[98] & ~t[99]) | (t[93] & ~t[94] & t[95] & t[96] & ~t[99]) | (t[93] & ~t[94] & t[97] & t[98] & ~t[99]) | (t[94] & ~t[96] & ~t[98] & t[99]) | (~t[94] & t[96] & t[98] & t[99]);
  assign t[8] = t[12] ^ t[13];
  assign t[90] = (t[93] & t[94] & t[95] & ~t[96] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & ~t[96] & ~t[97] & t[98] & t[99]) | (~t[94] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (~t[93] & ~t[95] & t[96] & ~t[98] & ~t[99]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[99]) | (~t[94] & t[95] & t[96] & t[97] & ~t[98]) | (~t[95] & t[96] & t[97] & ~t[99]);
  assign t[91] = (t[93] & t[94] & ~t[95] & ~t[97] & t[98] & ~t[99]) | (t[93] & t[95] & ~t[96] & ~t[97] & ~t[98] & t[99]) | (~t[94] & ~t[95] & t[97] & ~t[98] & ~t[99]) | (~t[93] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[93] & ~t[94] & ~t[96] & t[97] & ~t[99]) | (~t[93] & ~t[95] & t[96] & t[97] & t[98]) | (t[96] & t[97] & ~t[98] & ~t[99]);
  assign t[92] = (t[93] & t[94] & ~t[96] & t[97] & ~t[98] & ~t[99]) | (t[94] & ~t[95] & t[96] & ~t[97] & ~t[98] & t[99]) | (~t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[96] & ~t[97] & t[98] & ~t[99]) | (~t[93] & ~t[94] & ~t[95] & t[98] & ~t[99]) | (~t[94] & t[95] & ~t[96] & t[97] & t[98]) | (t[95] & ~t[97] & t[98] & ~t[99]);
  assign t[93] = t[114] ^ x[7];
  assign t[94] = t[115] ^ x[32];
  assign t[95] = t[116] ^ x[8];
  assign t[96] = t[117] ^ x[33];
  assign t[97] = t[118] ^ x[34];
  assign t[98] = t[119] ^ x[35];
  assign t[99] = t[120] ^ x[6];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0] & ~t[38]) | (~t[0] & t[38]);
endmodule

module R2ind96(x, y);
 input [35:0] x;
 output y;

 wire [132:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[15];
  assign t[101] = t[122] ^ x[18];
  assign t[102] = t[123] ^ x[16];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[13];
  assign t[105] = t[126] ^ x[25];
  assign t[106] = t[127] ^ x[28];
  assign t[107] = t[128] ^ x[26];
  assign t[108] = t[129] ^ x[29];
  assign t[109] = t[130] ^ x[27];
  assign t[10] = t[16] ^ t[17];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[24];
  assign t[112] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[113] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[114] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[115] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[116] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[117] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[118] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[119] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[11] = t[18] & t[19];
  assign t[120] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[121] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[122] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[123] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[124] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[125] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[126] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[127] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[128] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[129] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[12] = t[20] ^ t[11];
  assign t[130] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[131] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[132] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[46] ^ t[18];
  assign t[14] = t[21] ^ t[22];
  assign t[15] = t[23] ^ t[24];
  assign t[16] = t[47] ^ t[48];
  assign t[17] = t[18] & t[25];
  assign t[18] = ~(t[48]);
  assign t[19] = ~(t[46] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[46] & t[26];
  assign t[21] = t[27] ^ t[28];
  assign t[22] = t[29] & t[30];
  assign t[23] = t[31] ^ t[22];
  assign t[24] = t[49] ^ t[29];
  assign t[25] = t[46] ^ t[32];
  assign t[26] = t[33] ^ t[17];
  assign t[27] = t[50] ^ t[51];
  assign t[28] = t[29] & t[34];
  assign t[29] = ~(t[51]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[49] ^ t[29]);
  assign t[31] = t[49] & t[35];
  assign t[32] = t[48] ^ t[52];
  assign t[33] = t[46] ^ t[16];
  assign t[34] = t[49] ^ t[36];
  assign t[35] = t[37] ^ t[28];
  assign t[36] = t[51] ^ t[53];
  assign t[37] = t[49] ^ t[27];
  assign t[38] = x[0] ? x[31] : t[39];
  assign t[39] = ~(t[40] ^ t[41]);
  assign t[3] = ~(t[5]);
  assign t[40] = ~t[42];
  assign t[41] = ~(t[7]);
  assign t[42] = ~(t[43] ^ t[54]);
  assign t[43] = ~t[44];
  assign t[44] = ~(t[14]);
  assign t[45] = (t[55] & ~t[56]) | (~t[55] & t[56]);
  assign t[46] = (t[57] & ~t[58]) | (~t[57] & t[58]);
  assign t[47] = (t[57] & ~t[59]) | (~t[57] & t[59]);
  assign t[48] = (t[57] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[59]) | (~t[57] & ~t[61] & t[62]) | (t[60] & t[61] & t[59]);
  assign t[49] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[4] = ~(t[6] ^ t[45]);
  assign t[50] = (t[63] & ~t[65]) | (~t[63] & t[65]);
  assign t[51] = (t[63] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[65]) | (~t[63] & ~t[67] & t[68]) | (t[66] & t[67] & t[65]);
  assign t[52] = (t[57] & ~t[61] & ~t[59]) | (~t[60] & t[61] & ~t[62]) | (~t[57] & ~t[61] & t[59]) | (t[60] & t[61] & t[62]);
  assign t[53] = (t[63] & ~t[67] & ~t[65]) | (~t[66] & t[67] & ~t[68]) | (~t[63] & ~t[67] & t[65]) | (t[66] & t[67] & t[68]);
  assign t[54] = (t[55] & ~t[70] & ~t[71]) | (~t[69] & t[70] & ~t[72]) | (~t[55] & ~t[70] & t[71]) | (t[69] & t[70] & t[72]);
  assign t[55] = t[73] ^ x[7];
  assign t[56] = t[74] ^ x[8];
  assign t[57] = t[75] ^ x[14];
  assign t[58] = t[76] ^ x[15];
  assign t[59] = t[77] ^ x[16];
  assign t[5] = ~(t[7] ^ t[8]);
  assign t[60] = t[78] ^ x[17];
  assign t[61] = t[79] ^ x[18];
  assign t[62] = t[80] ^ x[19];
  assign t[63] = t[81] ^ x[25];
  assign t[64] = t[82] ^ x[26];
  assign t[65] = t[83] ^ x[27];
  assign t[66] = t[84] ^ x[28];
  assign t[67] = t[85] ^ x[29];
  assign t[68] = t[86] ^ x[30];
  assign t[69] = t[87] ^ x[32];
  assign t[6] = ~t[9];
  assign t[70] = t[88] ^ x[33];
  assign t[71] = t[89] ^ x[34];
  assign t[72] = t[90] ^ x[35];
  assign t[73] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[74] = (t[91] & t[92] & ~t[93] & t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[93] & ~t[94] & t[95] & ~t[96] & t[97]) | (~t[92] & t[93] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[92] & t[93] & ~t[96] & ~t[97]) | (~t[91] & t[93] & t[94] & ~t[95] & t[96]) | (t[93] & ~t[94] & t[96] & ~t[97]);
  assign t[75] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[76] = (t[98] & t[99] & ~t[100] & t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[100] & ~t[101] & t[102] & ~t[103] & t[104]) | (~t[99] & t[100] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[99] & t[100] & ~t[103] & ~t[104]) | (~t[98] & t[100] & t[101] & ~t[102] & t[103]) | (t[100] & ~t[101] & t[103] & ~t[104]);
  assign t[77] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[78] = (t[99] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & t[99] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[99] & ~t[100] & ~t[103] & ~t[104]) | (t[98] & ~t[99] & t[100] & t[101] & ~t[104]) | (t[98] & ~t[99] & t[102] & t[103] & ~t[104]) | (t[99] & ~t[101] & ~t[103] & t[104]) | (~t[99] & t[101] & t[103] & t[104]);
  assign t[79] = (t[98] & t[99] & t[100] & ~t[101] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[101] & ~t[102] & t[103] & t[104]) | (~t[99] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[100] & t[101] & ~t[103] & ~t[104]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[104]) | (~t[99] & t[100] & t[101] & t[102] & ~t[103]) | (~t[100] & t[101] & t[102] & ~t[104]);
  assign t[7] = t[10] ^ t[11];
  assign t[80] = (t[98] & t[99] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[98] & ~t[99] & ~t[100] & t[103] & ~t[104]) | (~t[99] & t[100] & ~t[101] & t[102] & t[103]) | (t[100] & ~t[102] & t[103] & ~t[104]);
  assign t[81] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[82] = (t[105] & t[106] & ~t[107] & t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[107] & ~t[108] & t[109] & ~t[110] & t[111]) | (~t[106] & t[107] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[106] & t[107] & ~t[110] & ~t[111]) | (~t[105] & t[107] & t[108] & ~t[109] & t[110]) | (t[107] & ~t[108] & t[110] & ~t[111]);
  assign t[83] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[84] = (t[106] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (~t[105] & t[106] & ~t[108] & ~t[109] & ~t[111]) | (~t[105] & t[106] & ~t[107] & ~t[110] & ~t[111]) | (t[105] & ~t[106] & t[107] & t[108] & ~t[111]) | (t[105] & ~t[106] & t[109] & t[110] & ~t[111]) | (t[106] & ~t[108] & ~t[110] & t[111]) | (~t[106] & t[108] & t[110] & t[111]);
  assign t[85] = (t[105] & t[106] & t[107] & ~t[108] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[108] & ~t[109] & t[110] & t[111]) | (~t[106] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (~t[105] & ~t[107] & t[108] & ~t[110] & ~t[111]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[111]) | (~t[106] & t[107] & t[108] & t[109] & ~t[110]) | (~t[107] & t[108] & t[109] & ~t[111]);
  assign t[86] = (t[105] & t[106] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[105] & ~t[106] & ~t[107] & t[110] & ~t[111]) | (~t[106] & t[107] & ~t[108] & t[109] & t[110]) | (t[107] & ~t[109] & t[110] & ~t[111]);
  assign t[87] = (t[92] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (~t[91] & t[92] & ~t[94] & ~t[95] & ~t[97]) | (~t[91] & t[92] & ~t[93] & ~t[96] & ~t[97]) | (t[91] & ~t[92] & t[93] & t[94] & ~t[97]) | (t[91] & ~t[92] & t[95] & t[96] & ~t[97]) | (t[92] & ~t[94] & ~t[96] & t[97]) | (~t[92] & t[94] & t[96] & t[97]);
  assign t[88] = (t[91] & t[92] & t[93] & ~t[94] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[94] & ~t[95] & t[96] & t[97]) | (~t[92] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (~t[91] & ~t[93] & t[94] & ~t[96] & ~t[97]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[97]) | (~t[92] & t[93] & t[94] & t[95] & ~t[96]) | (~t[93] & t[94] & t[95] & ~t[97]);
  assign t[89] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[8] = t[12] ^ t[13];
  assign t[90] = (t[91] & t[92] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[91] & ~t[92] & ~t[93] & t[96] & ~t[97]) | (~t[92] & t[93] & ~t[94] & t[95] & t[96]) | (t[93] & ~t[95] & t[96] & ~t[97]);
  assign t[91] = t[112] ^ x[7];
  assign t[92] = t[113] ^ x[32];
  assign t[93] = t[114] ^ x[8];
  assign t[94] = t[115] ^ x[33];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[35];
  assign t[97] = t[118] ^ x[6];
  assign t[98] = t[119] ^ x[14];
  assign t[99] = t[120] ^ x[17];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = (t[0] & ~t[38]) | (~t[0] & t[38]);
endmodule

module R2ind97(x, y);
 input [35:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[101] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[102] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[103] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[104] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[105] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[35]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[114] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[115] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[116] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[118] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[119] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[11] = ~(t[37] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[38] ^ t[39];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = x[0] ? x[35] : t[18];
  assign t[18] = ~(t[19] ^ t[20]);
  assign t[19] = ~t[21];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[23] ^ t[41]);
  assign t[22] = t[24] ^ t[8];
  assign t[23] = ~t[25];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = ~(t[28]);
  assign t[26] = t[42] ^ t[35];
  assign t[27] = t[10] & t[29];
  assign t[28] = t[30] ^ t[14];
  assign t[29] = t[37] ^ t[7];
  assign t[2] = ~t[4];
  assign t[30] = t[31] ^ t[32];
  assign t[31] = t[43] ^ t[38];
  assign t[32] = t[15] & t[33];
  assign t[33] = t[40] ^ t[13];
  assign t[34] = (t[44] & ~t[46] & ~t[48]) | (~t[45] & t[46] & ~t[47]) | (~t[44] & ~t[46] & t[48]) | (t[45] & t[46] & t[47]);
  assign t[35] = (t[49] & ~t[51] & ~t[53]) | (~t[50] & t[51] & ~t[52]) | (~t[49] & ~t[51] & t[53]) | (t[50] & t[51] & t[52]);
  assign t[36] = (t[49] & ~t[51] & ~t[52]) | (~t[50] & t[51] & ~t[53]) | (~t[49] & ~t[51] & t[52]) | (t[50] & t[51] & t[53]);
  assign t[37] = (t[49] & ~t[54]) | (~t[49] & t[54]);
  assign t[38] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[39] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[60]) | (~t[55] & t[60]);
  assign t[41] = (t[44] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[44] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[42] = (t[49] & ~t[52]) | (~t[49] & t[52]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = t[61] ^ x[8];
  assign t[45] = t[62] ^ x[9];
  assign t[46] = t[63] ^ x[10];
  assign t[47] = t[64] ^ x[11];
  assign t[48] = t[65] ^ x[12];
  assign t[49] = t[66] ^ x[18];
  assign t[4] = ~(t[6] ^ t[34]);
  assign t[50] = t[67] ^ x[19];
  assign t[51] = t[68] ^ x[20];
  assign t[52] = t[69] ^ x[21];
  assign t[53] = t[70] ^ x[22];
  assign t[54] = t[71] ^ x[23];
  assign t[55] = t[72] ^ x[29];
  assign t[56] = t[73] ^ x[30];
  assign t[57] = t[74] ^ x[31];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[34];
  assign t[61] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[62] = (t[79] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (~t[78] & t[79] & ~t[81] & ~t[82] & ~t[84]) | (~t[78] & t[79] & ~t[80] & ~t[83] & ~t[84]) | (t[78] & ~t[79] & t[80] & t[81] & ~t[84]) | (t[78] & ~t[79] & t[82] & t[83] & ~t[84]) | (t[79] & ~t[81] & ~t[83] & t[84]) | (~t[79] & t[81] & t[83] & t[84]);
  assign t[63] = (t[78] & t[79] & t[80] & ~t[81] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & ~t[81] & ~t[82] & t[83] & t[84]) | (~t[79] & ~t[80] & t[81] & ~t[82] & ~t[83]) | (~t[78] & ~t[80] & t[81] & ~t[83] & ~t[84]) | (~t[78] & ~t[79] & t[81] & ~t[82] & ~t[84]) | (~t[79] & t[80] & t[81] & t[82] & ~t[83]) | (~t[80] & t[81] & t[82] & ~t[84]);
  assign t[64] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[65] = (t[78] & t[79] & ~t[81] & t[82] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & ~t[81] & ~t[82] & t[83]) | (~t[78] & ~t[81] & ~t[82] & t[83] & ~t[84]) | (~t[78] & ~t[79] & ~t[80] & t[83] & ~t[84]) | (~t[79] & t[80] & ~t[81] & t[82] & t[83]) | (t[80] & ~t[82] & t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = ~t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[72] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[73] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[74] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[8];
  assign t[79] = t[100] ^ x[9];
  assign t[7] = t[35] ^ t[36];
  assign t[80] = t[101] ^ x[6];
  assign t[81] = t[102] ^ x[10];
  assign t[82] = t[103] ^ x[11];
  assign t[83] = t[104] ^ x[12];
  assign t[84] = t[105] ^ x[7];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[23];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[29];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[32];
  assign t[97] = t[118] ^ x[33];
  assign t[98] = t[119] ^ x[28];
  assign t[99] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~t[17]) | (~t[0] & t[17]);
endmodule

module R2ind98(x, y);
 input [52:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[122] ^ x[51];
  assign t[101] = t[123] ^ x[52];
  assign t[102] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[103] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[104] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[105] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[106] = (t[138] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[139] & ~t[140] & ~t[143] & ~t[144]) | (~t[138] & t[139] & t[140] & t[141] & ~t[144]) | (~t[138] & t[139] & t[142] & t[143] & ~t[144]) | (t[138] & ~t[140] & ~t[142] & t[144]) | (~t[138] & t[140] & t[142] & t[144]);
  assign t[107] = (t[138] & t[139] & ~t[140] & ~t[142] & t[143] & ~t[144]) | (t[138] & t[140] & ~t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & t[142] & ~t[143] & ~t[144]) | (~t[138] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[138] & ~t[139] & ~t[141] & t[142] & ~t[144]) | (~t[138] & ~t[140] & t[141] & t[142] & t[143]) | (t[141] & t[142] & ~t[143] & ~t[144]);
  assign t[108] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[109] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[111] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[112] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[113] = (t[145] & t[146] & ~t[147] & t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[147] & ~t[148] & t[149] & ~t[150] & t[151]) | (~t[146] & t[147] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[146] & t[147] & ~t[150] & ~t[151]) | (~t[145] & t[147] & t[148] & ~t[149] & t[150]) | (t[147] & ~t[148] & t[150] & ~t[151]);
  assign t[114] = (t[146] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & t[146] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[146] & ~t[147] & ~t[150] & ~t[151]) | (t[145] & ~t[146] & t[147] & t[148] & ~t[151]) | (t[145] & ~t[146] & t[149] & t[150] & ~t[151]) | (t[146] & ~t[148] & ~t[150] & t[151]) | (~t[146] & t[148] & t[150] & t[151]);
  assign t[115] = (t[145] & t[146] & t[147] & ~t[148] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & ~t[148] & ~t[149] & t[150] & t[151]) | (~t[146] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[147] & t[148] & ~t[150] & ~t[151]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[151]) | (~t[146] & t[147] & t[148] & t[149] & ~t[150]) | (~t[147] & t[148] & t[149] & ~t[151]);
  assign t[116] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[117] = (t[145] & t[146] & ~t[148] & t[149] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[148] & ~t[149] & t[150] & ~t[151]) | (~t[145] & ~t[146] & ~t[147] & t[150] & ~t[151]) | (~t[146] & t[147] & ~t[148] & t[149] & t[150]) | (t[147] & ~t[149] & t[150] & ~t[151]);
  assign t[118] = (t[124] & t[125] & ~t[126] & t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[126] & ~t[127] & t[128] & ~t[129] & t[130]) | (~t[125] & t[126] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[125] & t[126] & ~t[129] & ~t[130]) | (~t[124] & t[126] & t[127] & ~t[128] & t[129]) | (t[126] & ~t[127] & t[129] & ~t[130]);
  assign t[119] = (t[152] & ~t[154] & ~t[155] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & ~t[155] & ~t[156] & ~t[158]) | (t[152] & ~t[153] & ~t[154] & ~t[157] & ~t[158]) | (~t[152] & t[153] & t[154] & t[155] & ~t[158]) | (~t[152] & t[153] & t[156] & t[157] & ~t[158]) | (t[152] & ~t[154] & ~t[156] & t[158]) | (~t[152] & t[154] & t[156] & t[158]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (t[152] & t[153] & ~t[154] & ~t[156] & t[157] & ~t[158]) | (t[152] & t[154] & ~t[155] & ~t[156] & ~t[157] & t[158]) | (~t[153] & ~t[154] & t[156] & ~t[157] & ~t[158]) | (~t[152] & ~t[154] & ~t[155] & t[156] & ~t[157]) | (~t[152] & ~t[153] & ~t[155] & t[156] & ~t[158]) | (~t[152] & ~t[154] & t[155] & t[156] & t[157]) | (t[155] & t[156] & ~t[157] & ~t[158]);
  assign t[121] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[122] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[123] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[124] = t[159] ^ x[7];
  assign t[125] = t[160] ^ x[50];
  assign t[126] = t[161] ^ x[40];
  assign t[127] = t[162] ^ x[51];
  assign t[128] = t[163] ^ x[8];
  assign t[129] = t[164] ^ x[52];
  assign t[12] = ~(t[18] ^ t[69]);
  assign t[130] = t[165] ^ x[6];
  assign t[131] = t[166] ^ x[14];
  assign t[132] = t[167] ^ x[24];
  assign t[133] = t[168] ^ x[15];
  assign t[134] = t[169] ^ x[25];
  assign t[135] = t[170] ^ x[26];
  assign t[136] = t[171] ^ x[27];
  assign t[137] = t[172] ^ x[13];
  assign t[138] = t[173] ^ x[22];
  assign t[139] = t[174] ^ x[17];
  assign t[13] = t[19] ^ t[20];
  assign t[140] = t[175] ^ x[18];
  assign t[141] = t[176] ^ x[19];
  assign t[142] = t[177] ^ x[23];
  assign t[143] = t[178] ^ x[20];
  assign t[144] = t[179] ^ x[21];
  assign t[145] = t[180] ^ x[33];
  assign t[146] = t[181] ^ x[35];
  assign t[147] = t[182] ^ x[34];
  assign t[148] = t[183] ^ x[36];
  assign t[149] = t[184] ^ x[37];
  assign t[14] = ~(t[70]);
  assign t[150] = t[185] ^ x[38];
  assign t[151] = t[186] ^ x[32];
  assign t[152] = t[187] ^ x[47];
  assign t[153] = t[188] ^ x[42];
  assign t[154] = t[189] ^ x[43];
  assign t[155] = t[190] ^ x[44];
  assign t[156] = t[191] ^ x[48];
  assign t[157] = t[192] ^ x[45];
  assign t[158] = t[193] ^ x[46];
  assign t[159] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[15] = ~(t[68] ^ t[14]);
  assign t[160] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[161] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[162] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[163] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[164] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[165] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[166] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[167] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[168] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[169] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[16] = t[71] ^ t[70];
  assign t[170] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[171] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[172] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[173] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[174] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[175] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[176] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[177] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[178] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[179] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[180] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[181] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[182] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[183] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[184] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[185] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[186] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[187] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[188] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[189] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[18] = ~t[22];
  assign t[190] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[192] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[193] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = t[68] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[68] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[70] ^ t[72];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[73] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[74]);
  assign t[32] = ~(t[73] ^ t[31]);
  assign t[33] = t[75] ^ t[74];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[73] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[73] ^ t[38];
  assign t[38] = t[74] ^ t[76];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~(t[46] ^ t[77]);
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~t[49];
  assign t[47] = t[16] ^ t[20];
  assign t[48] = t[68] ^ t[14];
  assign t[49] = ~(t[50] ^ t[78]);
  assign t[4] = ~(t[7] ^ t[67]);
  assign t[50] = ~t[51];
  assign t[51] = ~(t[52] ^ t[53]);
  assign t[52] = t[54] ^ t[27];
  assign t[53] = t[24] ^ t[55];
  assign t[54] = t[33] ^ t[36];
  assign t[55] = t[73] ^ t[31];
  assign t[56] = x[0] ? x[49] : t[57];
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = ~(t[61]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[62] ^ t[79]);
  assign t[61] = t[23] ^ t[9];
  assign t[62] = ~t[63];
  assign t[63] = ~t[64];
  assign t[64] = ~t[65];
  assign t[65] = ~(t[66]);
  assign t[66] = t[38] ^ t[27];
  assign t[67] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[68] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[69] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[82] & ~t[87] & ~t[89]) | (~t[86] & t[87] & ~t[88]) | (~t[82] & ~t[87] & t[89]) | (t[86] & t[87] & t[88]);
  assign t[71] = (t[82] & ~t[88]) | (~t[82] & t[88]);
  assign t[72] = (t[82] & ~t[87] & ~t[88]) | (~t[86] & t[87] & ~t[89]) | (~t[82] & ~t[87] & t[88]) | (t[86] & t[87] & t[89]);
  assign t[73] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[74] = (t[90] & ~t[93] & ~t[95]) | (~t[92] & t[93] & ~t[94]) | (~t[90] & ~t[93] & t[95]) | (t[92] & t[93] & t[94]);
  assign t[75] = (t[90] & ~t[94]) | (~t[90] & t[94]);
  assign t[76] = (t[90] & ~t[93] & ~t[94]) | (~t[92] & t[93] & ~t[95]) | (~t[90] & ~t[93] & t[94]) | (t[92] & t[93] & t[95]);
  assign t[77] = (t[80] & ~t[96]) | (~t[80] & t[96]);
  assign t[78] = (t[97] & ~t[98]) | (~t[97] & t[98]);
  assign t[79] = (t[80] & ~t[100] & ~t[101]) | (~t[99] & t[100] & ~t[81]) | (~t[80] & ~t[100] & t[101]) | (t[99] & t[100] & t[81]);
  assign t[7] = ~t[12];
  assign t[80] = t[102] ^ x[7];
  assign t[81] = t[103] ^ x[8];
  assign t[82] = t[104] ^ x[14];
  assign t[83] = t[105] ^ x[15];
  assign t[84] = t[106] ^ x[22];
  assign t[85] = t[107] ^ x[23];
  assign t[86] = t[108] ^ x[24];
  assign t[87] = t[109] ^ x[25];
  assign t[88] = t[110] ^ x[26];
  assign t[89] = t[111] ^ x[27];
  assign t[8] = t[68] & t[13];
  assign t[90] = t[112] ^ x[33];
  assign t[91] = t[113] ^ x[34];
  assign t[92] = t[114] ^ x[35];
  assign t[93] = t[115] ^ x[36];
  assign t[94] = t[116] ^ x[37];
  assign t[95] = t[117] ^ x[38];
  assign t[96] = t[118] ^ x[40];
  assign t[97] = t[119] ^ x[47];
  assign t[98] = t[120] ^ x[48];
  assign t[99] = t[121] ^ x[50];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39] & ~t[56]) | (~t[0] & t[39] & ~t[56]) | (~t[0] & ~t[39] & t[56]) | (t[0] & t[39] & t[56]);
endmodule

module R2ind99(x, y);
 input [52:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[101] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[102] = (t[129] & ~t[131] & ~t[132] & ~t[133] & ~t[134]) | (t[129] & ~t[130] & ~t[132] & ~t[133] & ~t[135]) | (t[129] & ~t[130] & ~t[131] & ~t[134] & ~t[135]) | (~t[129] & t[130] & t[131] & t[132] & ~t[135]) | (~t[129] & t[130] & t[133] & t[134] & ~t[135]) | (t[129] & ~t[131] & ~t[133] & t[135]) | (~t[129] & t[131] & t[133] & t[135]);
  assign t[103] = (t[129] & t[130] & ~t[131] & t[132] & ~t[133] & ~t[135]) | (t[129] & ~t[131] & ~t[132] & t[133] & ~t[134] & t[135]) | (~t[130] & t[131] & ~t[132] & ~t[133] & ~t[135]) | (~t[129] & t[131] & ~t[132] & ~t[133] & ~t[134]) | (~t[129] & ~t[130] & t[131] & ~t[134] & ~t[135]) | (~t[129] & t[131] & t[132] & ~t[133] & t[134]) | (t[131] & ~t[132] & t[134] & ~t[135]);
  assign t[104] = (t[136] & ~t[138] & ~t[139] & ~t[140] & ~t[141]) | (t[136] & ~t[137] & ~t[139] & ~t[140] & ~t[142]) | (t[136] & ~t[137] & ~t[138] & ~t[141] & ~t[142]) | (~t[136] & t[137] & t[138] & t[139] & ~t[142]) | (~t[136] & t[137] & t[140] & t[141] & ~t[142]) | (t[136] & ~t[138] & ~t[140] & t[142]) | (~t[136] & t[138] & t[140] & t[142]);
  assign t[105] = (t[136] & t[137] & ~t[138] & ~t[140] & t[141] & ~t[142]) | (t[136] & t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[142]) | (~t[136] & ~t[138] & ~t[139] & t[140] & ~t[141]) | (~t[136] & ~t[137] & ~t[139] & t[140] & ~t[142]) | (~t[136] & ~t[138] & t[139] & t[140] & t[141]) | (t[139] & t[140] & ~t[141] & ~t[142]);
  assign t[106] = (t[130] & ~t[131] & ~t[132] & ~t[133] & ~t[134]) | (~t[129] & t[130] & ~t[132] & ~t[133] & ~t[135]) | (~t[129] & t[130] & ~t[131] & ~t[134] & ~t[135]) | (t[129] & ~t[130] & t[131] & t[132] & ~t[135]) | (t[129] & ~t[130] & t[133] & t[134] & ~t[135]) | (t[130] & ~t[132] & ~t[134] & t[135]) | (~t[130] & t[132] & t[134] & t[135]);
  assign t[107] = (t[129] & t[130] & t[131] & ~t[132] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[132] & ~t[133] & t[134] & t[135]) | (~t[130] & ~t[131] & t[132] & ~t[133] & ~t[134]) | (~t[129] & ~t[131] & t[132] & ~t[134] & ~t[135]) | (~t[129] & ~t[130] & t[132] & ~t[133] & ~t[135]) | (~t[130] & t[131] & t[132] & t[133] & ~t[134]) | (~t[131] & t[132] & t[133] & ~t[135]);
  assign t[108] = (t[129] & t[130] & ~t[131] & ~t[133] & t[134] & ~t[135]) | (t[129] & t[131] & ~t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[131] & t[133] & ~t[134] & ~t[135]) | (~t[129] & ~t[131] & ~t[132] & t[133] & ~t[134]) | (~t[129] & ~t[130] & ~t[132] & t[133] & ~t[135]) | (~t[129] & ~t[131] & t[132] & t[133] & t[134]) | (t[132] & t[133] & ~t[134] & ~t[135]);
  assign t[109] = (t[129] & t[130] & ~t[132] & t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[131] & ~t[132] & ~t[133] & t[134]) | (~t[129] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[129] & ~t[130] & ~t[131] & t[134] & ~t[135]) | (~t[130] & t[131] & ~t[132] & t[133] & t[134]) | (t[131] & ~t[133] & t[134] & ~t[135]);
  assign t[10] = t[16] ^ t[14];
  assign t[110] = (t[143] & ~t[145] & ~t[146] & ~t[147] & ~t[148]) | (t[143] & ~t[144] & ~t[146] & ~t[147] & ~t[149]) | (t[143] & ~t[144] & ~t[145] & ~t[148] & ~t[149]) | (~t[143] & t[144] & t[145] & t[146] & ~t[149]) | (~t[143] & t[144] & t[147] & t[148] & ~t[149]) | (t[143] & ~t[145] & ~t[147] & t[149]) | (~t[143] & t[145] & t[147] & t[149]);
  assign t[111] = (t[143] & t[144] & ~t[145] & t[146] & ~t[147] & ~t[149]) | (t[143] & ~t[145] & ~t[146] & t[147] & ~t[148] & t[149]) | (~t[144] & t[145] & ~t[146] & ~t[147] & ~t[149]) | (~t[143] & t[145] & ~t[146] & ~t[147] & ~t[148]) | (~t[143] & ~t[144] & t[145] & ~t[148] & ~t[149]) | (~t[143] & t[145] & t[146] & ~t[147] & t[148]) | (t[145] & ~t[146] & t[148] & ~t[149]);
  assign t[112] = (t[144] & ~t[145] & ~t[146] & ~t[147] & ~t[148]) | (~t[143] & t[144] & ~t[146] & ~t[147] & ~t[149]) | (~t[143] & t[144] & ~t[145] & ~t[148] & ~t[149]) | (t[143] & ~t[144] & t[145] & t[146] & ~t[149]) | (t[143] & ~t[144] & t[147] & t[148] & ~t[149]) | (t[144] & ~t[146] & ~t[148] & t[149]) | (~t[144] & t[146] & t[148] & t[149]);
  assign t[113] = (t[143] & t[144] & t[145] & ~t[146] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[146] & ~t[147] & t[148] & t[149]) | (~t[144] & ~t[145] & t[146] & ~t[147] & ~t[148]) | (~t[143] & ~t[145] & t[146] & ~t[148] & ~t[149]) | (~t[143] & ~t[144] & t[146] & ~t[147] & ~t[149]) | (~t[144] & t[145] & t[146] & t[147] & ~t[148]) | (~t[145] & t[146] & t[147] & ~t[149]);
  assign t[114] = (t[143] & t[144] & ~t[145] & ~t[147] & t[148] & ~t[149]) | (t[143] & t[145] & ~t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[145] & t[147] & ~t[148] & ~t[149]) | (~t[143] & ~t[145] & ~t[146] & t[147] & ~t[148]) | (~t[143] & ~t[144] & ~t[146] & t[147] & ~t[149]) | (~t[143] & ~t[145] & t[146] & t[147] & t[148]) | (t[146] & t[147] & ~t[148] & ~t[149]);
  assign t[115] = (t[143] & t[144] & ~t[146] & t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[145] & ~t[146] & ~t[147] & t[148]) | (~t[143] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[143] & ~t[144] & ~t[145] & t[148] & ~t[149]) | (~t[144] & t[145] & ~t[146] & t[147] & t[148]) | (t[145] & ~t[147] & t[148] & ~t[149]);
  assign t[116] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[117] = (t[150] & ~t[152] & ~t[153] & ~t[154] & ~t[155]) | (t[150] & ~t[151] & ~t[153] & ~t[154] & ~t[156]) | (t[150] & ~t[151] & ~t[152] & ~t[155] & ~t[156]) | (~t[150] & t[151] & t[152] & t[153] & ~t[156]) | (~t[150] & t[151] & t[154] & t[155] & ~t[156]) | (t[150] & ~t[152] & ~t[154] & t[156]) | (~t[150] & t[152] & t[154] & t[156]);
  assign t[118] = (t[150] & t[151] & ~t[152] & ~t[154] & t[155] & ~t[156]) | (t[150] & t[152] & ~t[153] & ~t[154] & ~t[155] & t[156]) | (~t[151] & ~t[152] & t[154] & ~t[155] & ~t[156]) | (~t[150] & ~t[152] & ~t[153] & t[154] & ~t[155]) | (~t[150] & ~t[151] & ~t[153] & t[154] & ~t[156]) | (~t[150] & ~t[152] & t[153] & t[154] & t[155]) | (t[153] & t[154] & ~t[155] & ~t[156]);
  assign t[119] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[121] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[122] = t[157] ^ x[7];
  assign t[123] = t[158] ^ x[50];
  assign t[124] = t[159] ^ x[40];
  assign t[125] = t[160] ^ x[51];
  assign t[126] = t[161] ^ x[8];
  assign t[127] = t[162] ^ x[52];
  assign t[128] = t[163] ^ x[6];
  assign t[129] = t[164] ^ x[14];
  assign t[12] = ~(t[18] ^ t[67]);
  assign t[130] = t[165] ^ x[24];
  assign t[131] = t[166] ^ x[15];
  assign t[132] = t[167] ^ x[25];
  assign t[133] = t[168] ^ x[26];
  assign t[134] = t[169] ^ x[27];
  assign t[135] = t[170] ^ x[13];
  assign t[136] = t[171] ^ x[22];
  assign t[137] = t[172] ^ x[17];
  assign t[138] = t[173] ^ x[18];
  assign t[139] = t[174] ^ x[19];
  assign t[13] = t[19] ^ t[20];
  assign t[140] = t[175] ^ x[23];
  assign t[141] = t[176] ^ x[20];
  assign t[142] = t[177] ^ x[21];
  assign t[143] = t[178] ^ x[33];
  assign t[144] = t[179] ^ x[35];
  assign t[145] = t[180] ^ x[34];
  assign t[146] = t[181] ^ x[36];
  assign t[147] = t[182] ^ x[37];
  assign t[148] = t[183] ^ x[38];
  assign t[149] = t[184] ^ x[32];
  assign t[14] = ~(t[68]);
  assign t[150] = t[185] ^ x[47];
  assign t[151] = t[186] ^ x[42];
  assign t[152] = t[187] ^ x[43];
  assign t[153] = t[188] ^ x[44];
  assign t[154] = t[189] ^ x[48];
  assign t[155] = t[190] ^ x[45];
  assign t[156] = t[191] ^ x[46];
  assign t[157] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[158] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[159] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[15] = ~(t[66] ^ t[14]);
  assign t[160] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[161] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[162] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[163] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[164] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[165] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[166] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[167] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[168] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[169] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[16] = t[69] ^ t[68];
  assign t[170] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[171] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[172] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[173] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[174] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[175] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[176] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[177] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[178] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[179] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[180] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[181] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[182] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[183] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[184] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[185] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[186] = (x[41] & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0);
  assign t[187] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[188] = (x[41] & ~1'b0) | (~x[41] & 1'b0);
  assign t[189] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[18] = ~t[22];
  assign t[190] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[19] = t[66] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[66] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[68] ^ t[70];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[71] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[72]);
  assign t[32] = ~(t[71] ^ t[31]);
  assign t[33] = t[73] ^ t[72];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[71] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[71] ^ t[38];
  assign t[38] = t[72] ^ t[74];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44] ^ t[45]);
  assign t[43] = ~(t[46] ^ t[75]);
  assign t[44] = t[47] ^ t[9];
  assign t[45] = t[5] ^ t[48];
  assign t[46] = ~t[49];
  assign t[47] = t[16] ^ t[20];
  assign t[48] = t[66] ^ t[14];
  assign t[49] = ~(t[50] ^ t[76]);
  assign t[4] = ~(t[7] ^ t[65]);
  assign t[50] = ~t[51];
  assign t[51] = ~(t[52] ^ t[53]);
  assign t[52] = t[54] ^ t[27];
  assign t[53] = t[24] ^ t[55];
  assign t[54] = t[33] ^ t[36];
  assign t[55] = t[71] ^ t[31];
  assign t[56] = x[0] ? x[49] : t[57];
  assign t[57] = ~(t[58] ^ t[59]);
  assign t[58] = ~t[60];
  assign t[59] = ~(t[44]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[61] ^ t[77]);
  assign t[61] = ~t[62];
  assign t[62] = ~t[63];
  assign t[63] = ~t[64];
  assign t[64] = ~(t[52]);
  assign t[65] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[66] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[67] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[68] = (t[80] & ~t[85] & ~t[87]) | (~t[84] & t[85] & ~t[86]) | (~t[80] & ~t[85] & t[87]) | (t[84] & t[85] & t[86]);
  assign t[69] = (t[80] & ~t[86]) | (~t[80] & t[86]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[80] & ~t[85] & ~t[86]) | (~t[84] & t[85] & ~t[87]) | (~t[80] & ~t[85] & t[86]) | (t[84] & t[85] & t[87]);
  assign t[71] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[72] = (t[88] & ~t[91] & ~t[93]) | (~t[90] & t[91] & ~t[92]) | (~t[88] & ~t[91] & t[93]) | (t[90] & t[91] & t[92]);
  assign t[73] = (t[88] & ~t[92]) | (~t[88] & t[92]);
  assign t[74] = (t[88] & ~t[91] & ~t[92]) | (~t[90] & t[91] & ~t[93]) | (~t[88] & ~t[91] & t[92]) | (t[90] & t[91] & t[93]);
  assign t[75] = (t[78] & ~t[94]) | (~t[78] & t[94]);
  assign t[76] = (t[95] & ~t[96]) | (~t[95] & t[96]);
  assign t[77] = (t[78] & ~t[98] & ~t[79]) | (~t[97] & t[98] & ~t[99]) | (~t[78] & ~t[98] & t[79]) | (t[97] & t[98] & t[99]);
  assign t[78] = t[100] ^ x[7];
  assign t[79] = t[101] ^ x[8];
  assign t[7] = ~t[12];
  assign t[80] = t[102] ^ x[14];
  assign t[81] = t[103] ^ x[15];
  assign t[82] = t[104] ^ x[22];
  assign t[83] = t[105] ^ x[23];
  assign t[84] = t[106] ^ x[24];
  assign t[85] = t[107] ^ x[25];
  assign t[86] = t[108] ^ x[26];
  assign t[87] = t[109] ^ x[27];
  assign t[88] = t[110] ^ x[33];
  assign t[89] = t[111] ^ x[34];
  assign t[8] = t[66] & t[13];
  assign t[90] = t[112] ^ x[35];
  assign t[91] = t[113] ^ x[36];
  assign t[92] = t[114] ^ x[37];
  assign t[93] = t[115] ^ x[38];
  assign t[94] = t[116] ^ x[40];
  assign t[95] = t[117] ^ x[47];
  assign t[96] = t[118] ^ x[48];
  assign t[97] = t[119] ^ x[50];
  assign t[98] = t[120] ^ x[51];
  assign t[99] = t[121] ^ x[52];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39] & ~t[56]) | (~t[0] & t[39] & ~t[56]) | (~t[0] & ~t[39] & t[56]) | (t[0] & t[39] & t[56]);
endmodule

module R2ind100(x, y);
 input [43:0] x;
 output y;

 wire [154:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] ^ x[41];
  assign t[101] = t[129] ^ x[6];
  assign t[102] = t[130] ^ x[42];
  assign t[103] = t[131] ^ x[9];
  assign t[104] = t[132] ^ x[43];
  assign t[105] = t[133] ^ x[7];
  assign t[106] = t[134] ^ x[15];
  assign t[107] = t[135] ^ x[25];
  assign t[108] = t[136] ^ x[16];
  assign t[109] = t[137] ^ x[26];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[138] ^ x[27];
  assign t[111] = t[139] ^ x[28];
  assign t[112] = t[140] ^ x[14];
  assign t[113] = t[141] ^ x[23];
  assign t[114] = t[142] ^ x[18];
  assign t[115] = t[143] ^ x[19];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[24];
  assign t[118] = t[146] ^ x[21];
  assign t[119] = t[147] ^ x[22];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[148] ^ x[34];
  assign t[121] = t[149] ^ x[36];
  assign t[122] = t[150] ^ x[35];
  assign t[123] = t[151] ^ x[37];
  assign t[124] = t[152] ^ x[38];
  assign t[125] = t[153] ^ x[39];
  assign t[126] = t[154] ^ x[33];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = ~(t[18] ^ t[52]);
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[135] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[136] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[137] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[138] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[139] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[141] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[142] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[143] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[144] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[29] & ~x[30] & ~x[31]) | (~x[29] & x[30] & ~x[31]) | (~x[29] & ~x[30] & x[31]) | (x[29] & x[30] & x[31]);
  assign t[149] = (x[29] & ~x[30] & ~x[32]) | (~x[29] & x[30] & ~x[32]) | (~x[29] & ~x[30] & x[32]) | (x[29] & x[30] & x[32]);
  assign t[14] = ~(t[53]);
  assign t[150] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[151] = (x[29] & ~x[32]) | (~x[29] & x[32]);
  assign t[152] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[153] = (x[30] & ~x[32]) | (~x[30] & x[32]);
  assign t[154] = (x[31] & ~x[32]) | (~x[31] & x[32]);
  assign t[15] = ~(t[51] ^ t[14]);
  assign t[16] = t[54] ^ t[53];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[51] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[51] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[53] ^ t[55];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[56] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[57]);
  assign t[32] = ~(t[56] ^ t[31]);
  assign t[33] = t[58] ^ t[57];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[56] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[56] ^ t[38];
  assign t[38] = t[57] ^ t[59];
  assign t[39] = x[0] ? x[40] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44]);
  assign t[43] = ~(t[45] ^ t[60]);
  assign t[44] = t[23] ^ t[9];
  assign t[45] = ~t[46];
  assign t[46] = ~t[47];
  assign t[47] = ~t[48];
  assign t[48] = ~(t[49]);
  assign t[49] = t[38] ^ t[27];
  assign t[4] = ~(t[7] ^ t[50]);
  assign t[50] = (t[61] & ~t[62]) | (~t[61] & t[62]);
  assign t[51] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[52] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[53] = (t[63] & ~t[68] & ~t[70]) | (~t[67] & t[68] & ~t[69]) | (~t[63] & ~t[68] & t[70]) | (t[67] & t[68] & t[69]);
  assign t[54] = (t[63] & ~t[69]) | (~t[63] & t[69]);
  assign t[55] = (t[63] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[70]) | (~t[63] & ~t[68] & t[69]) | (t[67] & t[68] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[71] & ~t[74] & ~t[76]) | (~t[73] & t[74] & ~t[75]) | (~t[71] & ~t[74] & t[76]) | (t[73] & t[74] & t[75]);
  assign t[58] = (t[71] & ~t[75]) | (~t[71] & t[75]);
  assign t[59] = (t[71] & ~t[74] & ~t[75]) | (~t[73] & t[74] & ~t[76]) | (~t[71] & ~t[74] & t[75]) | (t[73] & t[74] & t[76]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[61] & ~t[78] & ~t[79]) | (~t[77] & t[78] & ~t[62]) | (~t[61] & ~t[78] & t[79]) | (t[77] & t[78] & t[62]);
  assign t[61] = t[80] ^ x[8];
  assign t[62] = t[81] ^ x[9];
  assign t[63] = t[82] ^ x[15];
  assign t[64] = t[83] ^ x[16];
  assign t[65] = t[84] ^ x[23];
  assign t[66] = t[85] ^ x[24];
  assign t[67] = t[86] ^ x[25];
  assign t[68] = t[87] ^ x[26];
  assign t[69] = t[88] ^ x[27];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[89] ^ x[28];
  assign t[71] = t[90] ^ x[34];
  assign t[72] = t[91] ^ x[35];
  assign t[73] = t[92] ^ x[36];
  assign t[74] = t[93] ^ x[37];
  assign t[75] = t[94] ^ x[38];
  assign t[76] = t[95] ^ x[39];
  assign t[77] = t[96] ^ x[41];
  assign t[78] = t[97] ^ x[42];
  assign t[79] = t[98] ^ x[43];
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[83] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[84] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[85] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[86] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[87] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[89] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[8] = t[51] & t[13];
  assign t[90] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[91] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[92] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[93] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[94] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[95] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[96] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[97] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[98] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[99] = t[127] ^ x[8];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind101(x, y);
 input [43:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[101] & t[102] & ~t[104] & t[105] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[104] & ~t[105] & t[106] & ~t[107]) | (~t[101] & ~t[102] & ~t[103] & t[106] & ~t[107]) | (~t[102] & t[103] & ~t[104] & t[105] & t[106]) | (t[103] & ~t[105] & t[106] & ~t[107]);
  assign t[101] = t[129] ^ x[8];
  assign t[102] = t[130] ^ x[41];
  assign t[103] = t[131] ^ x[6];
  assign t[104] = t[132] ^ x[42];
  assign t[105] = t[133] ^ x[9];
  assign t[106] = t[134] ^ x[43];
  assign t[107] = t[135] ^ x[7];
  assign t[108] = t[136] ^ x[15];
  assign t[109] = t[137] ^ x[25];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[138] ^ x[16];
  assign t[111] = t[139] ^ x[26];
  assign t[112] = t[140] ^ x[27];
  assign t[113] = t[141] ^ x[28];
  assign t[114] = t[142] ^ x[14];
  assign t[115] = t[143] ^ x[23];
  assign t[116] = t[144] ^ x[18];
  assign t[117] = t[145] ^ x[19];
  assign t[118] = t[146] ^ x[20];
  assign t[119] = t[147] ^ x[24];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[148] ^ x[21];
  assign t[121] = t[149] ^ x[22];
  assign t[122] = t[150] ^ x[34];
  assign t[123] = t[151] ^ x[36];
  assign t[124] = t[152] ^ x[35];
  assign t[125] = t[153] ^ x[37];
  assign t[126] = t[154] ^ x[38];
  assign t[127] = t[155] ^ x[39];
  assign t[128] = t[156] ^ x[33];
  assign t[129] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = ~(t[18] ^ t[54]);
  assign t[130] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[131] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[132] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[133] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[134] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[135] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[136] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[137] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[138] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[139] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[13] = t[19] ^ t[20];
  assign t[140] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[141] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[142] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[143] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[144] = (x[17] & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0);
  assign t[145] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[146] = (x[17] & ~1'b0) | (~x[17] & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[149] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = ~(t[55]);
  assign t[150] = (x[29] & ~x[30] & ~x[31]) | (~x[29] & x[30] & ~x[31]) | (~x[29] & ~x[30] & x[31]) | (x[29] & x[30] & x[31]);
  assign t[151] = (x[29] & ~x[30] & ~x[32]) | (~x[29] & x[30] & ~x[32]) | (~x[29] & ~x[30] & x[32]) | (x[29] & x[30] & x[32]);
  assign t[152] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[153] = (x[29] & ~x[32]) | (~x[29] & x[32]);
  assign t[154] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[155] = (x[30] & ~x[32]) | (~x[30] & x[32]);
  assign t[156] = (x[31] & ~x[32]) | (~x[31] & x[32]);
  assign t[15] = ~(t[53] ^ t[14]);
  assign t[16] = t[56] ^ t[55];
  assign t[17] = ~(t[21] ^ t[10]);
  assign t[18] = ~t[22];
  assign t[19] = t[53] ^ t[16];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[14] & t[21];
  assign t[21] = t[53] ^ t[23];
  assign t[22] = t[24] ^ t[25];
  assign t[23] = t[55] ^ t[57];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] & t[29];
  assign t[26] = t[58] & t[30];
  assign t[27] = t[31] & t[32];
  assign t[28] = t[33] ^ t[31];
  assign t[29] = t[34] ^ t[27];
  assign t[2] = ~t[4];
  assign t[30] = t[35] ^ t[36];
  assign t[31] = ~(t[59]);
  assign t[32] = ~(t[58] ^ t[31]);
  assign t[33] = t[60] ^ t[59];
  assign t[34] = ~(t[37] ^ t[28]);
  assign t[35] = t[58] ^ t[33];
  assign t[36] = t[31] & t[37];
  assign t[37] = t[58] ^ t[38];
  assign t[38] = t[59] ^ t[61];
  assign t[39] = x[0] ? x[40] : t[40];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44]);
  assign t[43] = ~(t[45] ^ t[62]);
  assign t[44] = t[46] ^ t[9];
  assign t[45] = ~t[47];
  assign t[46] = t[16] ^ t[20];
  assign t[47] = ~t[48];
  assign t[48] = ~t[49];
  assign t[49] = ~(t[50]);
  assign t[4] = ~(t[7] ^ t[52]);
  assign t[50] = t[51] ^ t[27];
  assign t[51] = t[33] ^ t[36];
  assign t[52] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[53] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[54] = (t[67] & ~t[68]) | (~t[67] & t[68]);
  assign t[55] = (t[65] & ~t[70] & ~t[72]) | (~t[69] & t[70] & ~t[71]) | (~t[65] & ~t[70] & t[72]) | (t[69] & t[70] & t[71]);
  assign t[56] = (t[65] & ~t[71]) | (~t[65] & t[71]);
  assign t[57] = (t[65] & ~t[70] & ~t[71]) | (~t[69] & t[70] & ~t[72]) | (~t[65] & ~t[70] & t[71]) | (t[69] & t[70] & t[72]);
  assign t[58] = (t[73] & ~t[74]) | (~t[73] & t[74]);
  assign t[59] = (t[73] & ~t[76] & ~t[78]) | (~t[75] & t[76] & ~t[77]) | (~t[73] & ~t[76] & t[78]) | (t[75] & t[76] & t[77]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[73] & ~t[77]) | (~t[73] & t[77]);
  assign t[61] = (t[73] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[73] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[62] = (t[63] & ~t[80] & ~t[64]) | (~t[79] & t[80] & ~t[81]) | (~t[63] & ~t[80] & t[64]) | (t[79] & t[80] & t[81]);
  assign t[63] = t[82] ^ x[8];
  assign t[64] = t[83] ^ x[9];
  assign t[65] = t[84] ^ x[15];
  assign t[66] = t[85] ^ x[16];
  assign t[67] = t[86] ^ x[23];
  assign t[68] = t[87] ^ x[24];
  assign t[69] = t[88] ^ x[25];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[89] ^ x[26];
  assign t[71] = t[90] ^ x[27];
  assign t[72] = t[91] ^ x[28];
  assign t[73] = t[92] ^ x[34];
  assign t[74] = t[93] ^ x[35];
  assign t[75] = t[94] ^ x[36];
  assign t[76] = t[95] ^ x[37];
  assign t[77] = t[96] ^ x[38];
  assign t[78] = t[97] ^ x[39];
  assign t[79] = t[98] ^ x[41];
  assign t[7] = ~t[12];
  assign t[80] = t[99] ^ x[42];
  assign t[81] = t[100] ^ x[43];
  assign t[82] = (t[101] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & ~t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[102] & ~t[103] & ~t[106] & ~t[107]) | (~t[101] & t[102] & t[103] & t[104] & ~t[107]) | (~t[101] & t[102] & t[105] & t[106] & ~t[107]) | (t[101] & ~t[103] & ~t[105] & t[107]) | (~t[101] & t[103] & t[105] & t[107]);
  assign t[83] = (t[101] & t[102] & ~t[103] & ~t[105] & t[106] & ~t[107]) | (t[101] & t[103] & ~t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & t[105] & ~t[106] & ~t[107]) | (~t[101] & ~t[103] & ~t[104] & t[105] & ~t[106]) | (~t[101] & ~t[102] & ~t[104] & t[105] & ~t[107]) | (~t[101] & ~t[103] & t[104] & t[105] & t[106]) | (t[104] & t[105] & ~t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[85] = (t[108] & t[109] & ~t[110] & t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[110] & ~t[111] & t[112] & ~t[113] & t[114]) | (~t[109] & t[110] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[109] & t[110] & ~t[113] & ~t[114]) | (~t[108] & t[110] & t[111] & ~t[112] & t[113]) | (t[110] & ~t[111] & t[113] & ~t[114]);
  assign t[86] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[87] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[88] = (t[109] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & t[109] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[109] & ~t[110] & ~t[113] & ~t[114]) | (t[108] & ~t[109] & t[110] & t[111] & ~t[114]) | (t[108] & ~t[109] & t[112] & t[113] & ~t[114]) | (t[109] & ~t[111] & ~t[113] & t[114]) | (~t[109] & t[111] & t[113] & t[114]);
  assign t[89] = (t[108] & t[109] & t[110] & ~t[111] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[111] & ~t[112] & t[113] & t[114]) | (~t[109] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[110] & t[111] & ~t[113] & ~t[114]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[114]) | (~t[109] & t[110] & t[111] & t[112] & ~t[113]) | (~t[110] & t[111] & t[112] & ~t[114]);
  assign t[8] = t[53] & t[13];
  assign t[90] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[91] = (t[108] & t[109] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[108] & ~t[109] & ~t[110] & t[113] & ~t[114]) | (~t[109] & t[110] & ~t[111] & t[112] & t[113]) | (t[110] & ~t[112] & t[113] & ~t[114]);
  assign t[92] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[93] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[94] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[95] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[96] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[97] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[98] = (t[102] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & t[102] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[102] & ~t[103] & ~t[106] & ~t[107]) | (t[101] & ~t[102] & t[103] & t[104] & ~t[107]) | (t[101] & ~t[102] & t[105] & t[106] & ~t[107]) | (t[102] & ~t[104] & ~t[106] & t[107]) | (~t[102] & t[104] & t[106] & t[107]);
  assign t[99] = (t[101] & t[102] & t[103] & ~t[104] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & ~t[104] & ~t[105] & t[106] & t[107]) | (~t[102] & ~t[103] & t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[103] & t[104] & ~t[106] & ~t[107]) | (~t[101] & ~t[102] & t[104] & ~t[105] & ~t[107]) | (~t[102] & t[103] & t[104] & t[105] & ~t[106]) | (~t[103] & t[104] & t[105] & ~t[107]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind102(x, y);
 input [43:0] x;
 output y;

 wire [156:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[101] & t[102] & ~t[104] & t[105] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & ~t[104] & ~t[105] & t[106]) | (~t[101] & ~t[104] & ~t[105] & t[106] & ~t[107]) | (~t[101] & ~t[102] & ~t[103] & t[106] & ~t[107]) | (~t[102] & t[103] & ~t[104] & t[105] & t[106]) | (t[103] & ~t[105] & t[106] & ~t[107]);
  assign t[101] = t[129] ^ x[7];
  assign t[102] = t[130] ^ x[40];
  assign t[103] = t[131] ^ x[8];
  assign t[104] = t[132] ^ x[41];
  assign t[105] = t[133] ^ x[42];
  assign t[106] = t[134] ^ x[43];
  assign t[107] = t[135] ^ x[6];
  assign t[108] = t[136] ^ x[14];
  assign t[109] = t[137] ^ x[25];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[138] ^ x[15];
  assign t[111] = t[139] ^ x[26];
  assign t[112] = t[140] ^ x[24];
  assign t[113] = t[141] ^ x[27];
  assign t[114] = t[142] ^ x[13];
  assign t[115] = t[143] ^ x[22];
  assign t[116] = t[144] ^ x[17];
  assign t[117] = t[145] ^ x[18];
  assign t[118] = t[146] ^ x[19];
  assign t[119] = t[147] ^ x[23];
  assign t[11] = t[51] ^ t[15];
  assign t[120] = t[148] ^ x[20];
  assign t[121] = t[149] ^ x[21];
  assign t[122] = t[150] ^ x[33];
  assign t[123] = t[151] ^ x[36];
  assign t[124] = t[152] ^ x[34];
  assign t[125] = t[153] ^ x[37];
  assign t[126] = t[154] ^ x[35];
  assign t[127] = t[155] ^ x[38];
  assign t[128] = t[156] ^ x[32];
  assign t[129] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = ~(t[18] ^ t[52]);
  assign t[130] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[131] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[132] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[133] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[134] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[135] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[136] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[137] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[138] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[139] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[13] = t[53] ^ t[54];
  assign t[140] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[141] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[142] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[143] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[144] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[145] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[146] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[149] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[14] = t[15] & t[19];
  assign t[150] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[151] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[152] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[153] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[154] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[155] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[156] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[15] = ~(t[54]);
  assign t[16] = ~(t[51] ^ t[15]);
  assign t[17] = t[51] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[51] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[54] ^ t[55];
  assign t[23] = t[51] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[56] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[57] ^ t[58];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[58]);
  assign t[33] = ~(t[56] ^ t[32]);
  assign t[34] = t[56] & t[36];
  assign t[35] = t[56] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[58] ^ t[59];
  assign t[38] = t[56] ^ t[30];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[44]);
  assign t[43] = ~(t[45] ^ t[60]);
  assign t[44] = t[22] ^ t[9];
  assign t[45] = ~t[46];
  assign t[46] = ~t[47];
  assign t[47] = ~t[48];
  assign t[48] = ~(t[49]);
  assign t[49] = t[37] ^ t[27];
  assign t[4] = ~(t[7] ^ t[50]);
  assign t[50] = (t[61] & ~t[62]) | (~t[61] & t[62]);
  assign t[51] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[52] = (t[65] & ~t[66]) | (~t[65] & t[66]);
  assign t[53] = (t[63] & ~t[67]) | (~t[63] & t[67]);
  assign t[54] = (t[63] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[67]) | (~t[63] & ~t[69] & t[70]) | (t[68] & t[69] & t[67]);
  assign t[55] = (t[63] & ~t[69] & ~t[67]) | (~t[68] & t[69] & ~t[70]) | (~t[63] & ~t[69] & t[67]) | (t[68] & t[69] & t[70]);
  assign t[56] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[57] = (t[71] & ~t[73]) | (~t[71] & t[73]);
  assign t[58] = (t[71] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[73]) | (~t[71] & ~t[75] & t[76]) | (t[74] & t[75] & t[73]);
  assign t[59] = (t[71] & ~t[75] & ~t[73]) | (~t[74] & t[75] & ~t[76]) | (~t[71] & ~t[75] & t[73]) | (t[74] & t[75] & t[76]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[61] & ~t[78] & ~t[80]) | (~t[77] & t[78] & ~t[79]) | (~t[61] & ~t[78] & t[80]) | (t[77] & t[78] & t[79]);
  assign t[61] = t[81] ^ x[7];
  assign t[62] = t[82] ^ x[8];
  assign t[63] = t[83] ^ x[14];
  assign t[64] = t[84] ^ x[15];
  assign t[65] = t[85] ^ x[22];
  assign t[66] = t[86] ^ x[23];
  assign t[67] = t[87] ^ x[24];
  assign t[68] = t[88] ^ x[25];
  assign t[69] = t[89] ^ x[26];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[33];
  assign t[72] = t[92] ^ x[34];
  assign t[73] = t[93] ^ x[35];
  assign t[74] = t[94] ^ x[36];
  assign t[75] = t[95] ^ x[37];
  assign t[76] = t[96] ^ x[38];
  assign t[77] = t[97] ^ x[40];
  assign t[78] = t[98] ^ x[41];
  assign t[79] = t[99] ^ x[42];
  assign t[7] = ~t[12];
  assign t[80] = t[100] ^ x[43];
  assign t[81] = (t[101] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (t[101] & ~t[102] & ~t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[102] & ~t[103] & ~t[106] & ~t[107]) | (~t[101] & t[102] & t[103] & t[104] & ~t[107]) | (~t[101] & t[102] & t[105] & t[106] & ~t[107]) | (t[101] & ~t[103] & ~t[105] & t[107]) | (~t[101] & t[103] & t[105] & t[107]);
  assign t[82] = (t[101] & t[102] & ~t[103] & t[104] & ~t[105] & ~t[107]) | (t[101] & ~t[103] & ~t[104] & t[105] & ~t[106] & t[107]) | (~t[102] & t[103] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[102] & t[103] & ~t[106] & ~t[107]) | (~t[101] & t[103] & t[104] & ~t[105] & t[106]) | (t[103] & ~t[104] & t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[84] = (t[108] & t[109] & ~t[110] & t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[110] & ~t[111] & t[112] & ~t[113] & t[114]) | (~t[109] & t[110] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[109] & t[110] & ~t[113] & ~t[114]) | (~t[108] & t[110] & t[111] & ~t[112] & t[113]) | (t[110] & ~t[111] & t[113] & ~t[114]);
  assign t[85] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[86] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[87] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[88] = (t[109] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & t[109] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[109] & ~t[110] & ~t[113] & ~t[114]) | (t[108] & ~t[109] & t[110] & t[111] & ~t[114]) | (t[108] & ~t[109] & t[112] & t[113] & ~t[114]) | (t[109] & ~t[111] & ~t[113] & t[114]) | (~t[109] & t[111] & t[113] & t[114]);
  assign t[89] = (t[108] & t[109] & t[110] & ~t[111] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[111] & ~t[112] & t[113] & t[114]) | (~t[109] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[110] & t[111] & ~t[113] & ~t[114]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[114]) | (~t[109] & t[110] & t[111] & t[112] & ~t[113]) | (~t[110] & t[111] & t[112] & ~t[114]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[108] & t[109] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[108] & ~t[109] & ~t[110] & t[113] & ~t[114]) | (~t[109] & t[110] & ~t[111] & t[112] & t[113]) | (t[110] & ~t[112] & t[113] & ~t[114]);
  assign t[91] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[92] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[93] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[94] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[95] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[96] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[97] = (t[102] & ~t[103] & ~t[104] & ~t[105] & ~t[106]) | (~t[101] & t[102] & ~t[104] & ~t[105] & ~t[107]) | (~t[101] & t[102] & ~t[103] & ~t[106] & ~t[107]) | (t[101] & ~t[102] & t[103] & t[104] & ~t[107]) | (t[101] & ~t[102] & t[105] & t[106] & ~t[107]) | (t[102] & ~t[104] & ~t[106] & t[107]) | (~t[102] & t[104] & t[106] & t[107]);
  assign t[98] = (t[101] & t[102] & t[103] & ~t[104] & ~t[106] & ~t[107]) | (t[102] & ~t[103] & ~t[104] & ~t[105] & t[106] & t[107]) | (~t[102] & ~t[103] & t[104] & ~t[105] & ~t[106]) | (~t[101] & ~t[103] & t[104] & ~t[106] & ~t[107]) | (~t[101] & ~t[102] & t[104] & ~t[105] & ~t[107]) | (~t[102] & t[103] & t[104] & t[105] & ~t[106]) | (~t[103] & t[104] & t[105] & ~t[107]);
  assign t[99] = (t[101] & t[102] & ~t[103] & ~t[105] & t[106] & ~t[107]) | (t[101] & t[103] & ~t[104] & ~t[105] & ~t[106] & t[107]) | (~t[102] & ~t[103] & t[105] & ~t[106] & ~t[107]) | (~t[101] & ~t[103] & ~t[104] & t[105] & ~t[106]) | (~t[101] & ~t[102] & ~t[104] & t[105] & ~t[107]) | (~t[101] & ~t[103] & t[104] & t[105] & t[106]) | (t[104] & t[105] & ~t[106] & ~t[107]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind103(x, y);
 input [43:0] x;
 output y;

 wire [154:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] ^ x[40];
  assign t[101] = t[129] ^ x[8];
  assign t[102] = t[130] ^ x[41];
  assign t[103] = t[131] ^ x[42];
  assign t[104] = t[132] ^ x[43];
  assign t[105] = t[133] ^ x[6];
  assign t[106] = t[134] ^ x[14];
  assign t[107] = t[135] ^ x[25];
  assign t[108] = t[136] ^ x[15];
  assign t[109] = t[137] ^ x[26];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[138] ^ x[24];
  assign t[111] = t[139] ^ x[27];
  assign t[112] = t[140] ^ x[13];
  assign t[113] = t[141] ^ x[22];
  assign t[114] = t[142] ^ x[17];
  assign t[115] = t[143] ^ x[18];
  assign t[116] = t[144] ^ x[19];
  assign t[117] = t[145] ^ x[23];
  assign t[118] = t[146] ^ x[20];
  assign t[119] = t[147] ^ x[21];
  assign t[11] = t[49] ^ t[15];
  assign t[120] = t[148] ^ x[33];
  assign t[121] = t[149] ^ x[36];
  assign t[122] = t[150] ^ x[34];
  assign t[123] = t[151] ^ x[37];
  assign t[124] = t[152] ^ x[35];
  assign t[125] = t[153] ^ x[38];
  assign t[126] = t[154] ^ x[32];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = ~(t[18] ^ t[50]);
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[135] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[136] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[137] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[138] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[139] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[13] = t[51] ^ t[52];
  assign t[140] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[141] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[142] = (x[16] & ~1'b0 & ~1'b0) | (~x[16] & 1'b0 & ~1'b0) | (~x[16] & ~1'b0 & 1'b0) | (x[16] & 1'b0 & 1'b0);
  assign t[143] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[144] = (x[16] & ~1'b0) | (~x[16] & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[148] = (x[28] & ~x[29] & ~x[30]) | (~x[28] & x[29] & ~x[30]) | (~x[28] & ~x[29] & x[30]) | (x[28] & x[29] & x[30]);
  assign t[149] = (x[28] & ~x[29] & ~x[31]) | (~x[28] & x[29] & ~x[31]) | (~x[28] & ~x[29] & x[31]) | (x[28] & x[29] & x[31]);
  assign t[14] = t[15] & t[19];
  assign t[150] = (x[28] & ~x[30]) | (~x[28] & x[30]);
  assign t[151] = (x[28] & ~x[31]) | (~x[28] & x[31]);
  assign t[152] = (x[29] & ~x[30]) | (~x[29] & x[30]);
  assign t[153] = (x[29] & ~x[31]) | (~x[29] & x[31]);
  assign t[154] = (x[30] & ~x[31]) | (~x[30] & x[31]);
  assign t[15] = ~(t[52]);
  assign t[16] = ~(t[49] ^ t[15]);
  assign t[17] = t[49] & t[20];
  assign t[18] = ~t[21];
  assign t[19] = t[49] ^ t[22];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[23] ^ t[14];
  assign t[21] = ~(t[24] ^ t[25]);
  assign t[22] = t[52] ^ t[53];
  assign t[23] = t[49] ^ t[13];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = t[28] ^ t[29];
  assign t[26] = t[30] ^ t[31];
  assign t[27] = t[32] & t[33];
  assign t[28] = t[34] ^ t[27];
  assign t[29] = t[54] ^ t[32];
  assign t[2] = ~t[4];
  assign t[30] = t[55] ^ t[56];
  assign t[31] = t[32] & t[35];
  assign t[32] = ~(t[56]);
  assign t[33] = ~(t[54] ^ t[32]);
  assign t[34] = t[54] & t[36];
  assign t[35] = t[54] ^ t[37];
  assign t[36] = t[38] ^ t[31];
  assign t[37] = t[56] ^ t[57];
  assign t[38] = t[54] ^ t[30];
  assign t[39] = x[0] ? x[39] : t[40];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[41] ^ t[42]);
  assign t[41] = ~t[43];
  assign t[42] = ~(t[5]);
  assign t[43] = ~(t[44] ^ t[58]);
  assign t[44] = ~t[45];
  assign t[45] = ~t[46];
  assign t[46] = ~t[47];
  assign t[47] = ~(t[24]);
  assign t[48] = (t[59] & ~t[60]) | (~t[59] & t[60]);
  assign t[49] = (t[61] & ~t[62]) | (~t[61] & t[62]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[51] = (t[61] & ~t[65]) | (~t[61] & t[65]);
  assign t[52] = (t[61] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[65]) | (~t[61] & ~t[67] & t[68]) | (t[66] & t[67] & t[65]);
  assign t[53] = (t[61] & ~t[67] & ~t[65]) | (~t[66] & t[67] & ~t[68]) | (~t[61] & ~t[67] & t[65]) | (t[66] & t[67] & t[68]);
  assign t[54] = (t[69] & ~t[70]) | (~t[69] & t[70]);
  assign t[55] = (t[69] & ~t[71]) | (~t[69] & t[71]);
  assign t[56] = (t[69] & ~t[73] & ~t[74]) | (~t[72] & t[73] & ~t[71]) | (~t[69] & ~t[73] & t[74]) | (t[72] & t[73] & t[71]);
  assign t[57] = (t[69] & ~t[73] & ~t[71]) | (~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[73] & t[71]) | (t[72] & t[73] & t[74]);
  assign t[58] = (t[59] & ~t[76] & ~t[77]) | (~t[75] & t[76] & ~t[78]) | (~t[59] & ~t[76] & t[77]) | (t[75] & t[76] & t[78]);
  assign t[59] = t[79] ^ x[7];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[80] ^ x[8];
  assign t[61] = t[81] ^ x[14];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[22];
  assign t[64] = t[84] ^ x[23];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[25];
  assign t[67] = t[87] ^ x[26];
  assign t[68] = t[88] ^ x[27];
  assign t[69] = t[89] ^ x[33];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[90] ^ x[34];
  assign t[71] = t[91] ^ x[35];
  assign t[72] = t[92] ^ x[36];
  assign t[73] = t[93] ^ x[37];
  assign t[74] = t[94] ^ x[38];
  assign t[75] = t[95] ^ x[40];
  assign t[76] = t[96] ^ x[41];
  assign t[77] = t[97] ^ x[42];
  assign t[78] = t[98] ^ x[43];
  assign t[79] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[82] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[83] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[84] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[85] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[86] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[87] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[91] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[92] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[93] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[94] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[95] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[96] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[97] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[98] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[99] = t[127] ^ x[7];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[39]) | (~t[0] & t[39]);
endmodule

module R2ind104(x, y);
 input [35:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[32];
  assign t[101] = t[122] ^ x[33];
  assign t[102] = t[123] ^ x[28];
  assign t[103] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[104] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[105] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[106] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[107] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[108] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[109] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[10] = ~(t[39]);
  assign t[110] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[111] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[112] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[113] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[114] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[115] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[116] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[117] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[118] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[119] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[11] = ~(t[41] ^ t[10]);
  assign t[120] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[121] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[122] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[123] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[12] = ~t[13];
  assign t[13] = ~(t[14]);
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[42] ^ t[43];
  assign t[16] = t[17] & t[18];
  assign t[17] = ~(t[42]);
  assign t[18] = ~(t[44] ^ t[17]);
  assign t[19] = x[0] ? x[35] : t[20];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[21] ^ t[22]);
  assign t[21] = ~t[23];
  assign t[22] = ~(t[24]);
  assign t[23] = ~(t[25] ^ t[45]);
  assign t[24] = t[26] ^ t[8];
  assign t[25] = ~t[27];
  assign t[26] = t[28] ^ t[29];
  assign t[27] = ~t[30];
  assign t[28] = t[46] ^ t[39];
  assign t[29] = t[10] & t[31];
  assign t[2] = ~t[4];
  assign t[30] = ~t[32];
  assign t[31] = t[41] ^ t[7];
  assign t[32] = ~(t[33]);
  assign t[33] = t[34] ^ t[16];
  assign t[34] = t[35] ^ t[36];
  assign t[35] = t[47] ^ t[42];
  assign t[36] = t[17] & t[37];
  assign t[37] = t[44] ^ t[15];
  assign t[38] = (t[48] & ~t[50] & ~t[52]) | (~t[49] & t[50] & ~t[51]) | (~t[48] & ~t[50] & t[52]) | (t[49] & t[50] & t[51]);
  assign t[39] = (t[53] & ~t[55] & ~t[57]) | (~t[54] & t[55] & ~t[56]) | (~t[53] & ~t[55] & t[57]) | (t[54] & t[55] & t[56]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[53] & ~t[55] & ~t[56]) | (~t[54] & t[55] & ~t[57]) | (~t[53] & ~t[55] & t[56]) | (t[54] & t[55] & t[57]);
  assign t[41] = (t[53] & ~t[58]) | (~t[53] & t[58]);
  assign t[42] = (t[59] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[59] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[43] = (t[59] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[59] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[44] = (t[59] & ~t[64]) | (~t[59] & t[64]);
  assign t[45] = (t[48] & ~t[50] & ~t[51]) | (~t[49] & t[50] & ~t[52]) | (~t[48] & ~t[50] & t[51]) | (t[49] & t[50] & t[52]);
  assign t[46] = (t[53] & ~t[56]) | (~t[53] & t[56]);
  assign t[47] = (t[59] & ~t[62]) | (~t[59] & t[62]);
  assign t[48] = t[65] ^ x[8];
  assign t[49] = t[66] ^ x[9];
  assign t[4] = ~(t[6] ^ t[38]);
  assign t[50] = t[67] ^ x[10];
  assign t[51] = t[68] ^ x[11];
  assign t[52] = t[69] ^ x[12];
  assign t[53] = t[70] ^ x[18];
  assign t[54] = t[71] ^ x[19];
  assign t[55] = t[72] ^ x[20];
  assign t[56] = t[73] ^ x[21];
  assign t[57] = t[74] ^ x[22];
  assign t[58] = t[75] ^ x[23];
  assign t[59] = t[76] ^ x[29];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[30];
  assign t[61] = t[78] ^ x[31];
  assign t[62] = t[79] ^ x[32];
  assign t[63] = t[80] ^ x[33];
  assign t[64] = t[81] ^ x[34];
  assign t[65] = (t[82] & ~t[84] & ~t[85] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & ~t[85] & ~t[86] & ~t[88]) | (t[82] & ~t[83] & ~t[84] & ~t[87] & ~t[88]) | (~t[82] & t[83] & t[84] & t[85] & ~t[88]) | (~t[82] & t[83] & t[86] & t[87] & ~t[88]) | (t[82] & ~t[84] & ~t[86] & t[88]) | (~t[82] & t[84] & t[86] & t[88]);
  assign t[66] = (t[83] & ~t[84] & ~t[85] & ~t[86] & ~t[87]) | (~t[82] & t[83] & ~t[85] & ~t[86] & ~t[88]) | (~t[82] & t[83] & ~t[84] & ~t[87] & ~t[88]) | (t[82] & ~t[83] & t[84] & t[85] & ~t[88]) | (t[82] & ~t[83] & t[86] & t[87] & ~t[88]) | (t[83] & ~t[85] & ~t[87] & t[88]) | (~t[83] & t[85] & t[87] & t[88]);
  assign t[67] = (t[82] & t[83] & t[84] & ~t[85] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[85] & ~t[86] & t[87] & t[88]) | (~t[83] & ~t[84] & t[85] & ~t[86] & ~t[87]) | (~t[82] & ~t[84] & t[85] & ~t[87] & ~t[88]) | (~t[82] & ~t[83] & t[85] & ~t[86] & ~t[88]) | (~t[83] & t[84] & t[85] & t[86] & ~t[87]) | (~t[84] & t[85] & t[86] & ~t[88]);
  assign t[68] = (t[82] & t[83] & ~t[84] & ~t[86] & t[87] & ~t[88]) | (t[82] & t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[88]) | (~t[82] & ~t[84] & ~t[85] & t[86] & ~t[87]) | (~t[82] & ~t[83] & ~t[85] & t[86] & ~t[88]) | (~t[82] & ~t[84] & t[85] & t[86] & t[87]) | (t[85] & t[86] & ~t[87] & ~t[88]);
  assign t[69] = (t[82] & t[83] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[82] & ~t[83] & ~t[84] & t[87] & ~t[88]) | (~t[83] & t[84] & ~t[85] & t[86] & t[87]) | (t[84] & ~t[86] & t[87] & ~t[88]);
  assign t[6] = ~t[9];
  assign t[70] = (t[89] & ~t[91] & ~t[92] & ~t[93] & ~t[94]) | (t[89] & ~t[90] & ~t[92] & ~t[93] & ~t[95]) | (t[89] & ~t[90] & ~t[91] & ~t[94] & ~t[95]) | (~t[89] & t[90] & t[91] & t[92] & ~t[95]) | (~t[89] & t[90] & t[93] & t[94] & ~t[95]) | (t[89] & ~t[91] & ~t[93] & t[95]) | (~t[89] & t[91] & t[93] & t[95]);
  assign t[71] = (t[90] & ~t[91] & ~t[92] & ~t[93] & ~t[94]) | (~t[89] & t[90] & ~t[92] & ~t[93] & ~t[95]) | (~t[89] & t[90] & ~t[91] & ~t[94] & ~t[95]) | (t[89] & ~t[90] & t[91] & t[92] & ~t[95]) | (t[89] & ~t[90] & t[93] & t[94] & ~t[95]) | (t[90] & ~t[92] & ~t[94] & t[95]) | (~t[90] & t[92] & t[94] & t[95]);
  assign t[72] = (t[89] & t[90] & t[91] & ~t[92] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[92] & ~t[93] & t[94] & t[95]) | (~t[90] & ~t[91] & t[92] & ~t[93] & ~t[94]) | (~t[89] & ~t[91] & t[92] & ~t[94] & ~t[95]) | (~t[89] & ~t[90] & t[92] & ~t[93] & ~t[95]) | (~t[90] & t[91] & t[92] & t[93] & ~t[94]) | (~t[91] & t[92] & t[93] & ~t[95]);
  assign t[73] = (t[89] & t[90] & ~t[91] & ~t[93] & t[94] & ~t[95]) | (t[89] & t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[95]) | (~t[89] & ~t[91] & ~t[92] & t[93] & ~t[94]) | (~t[89] & ~t[90] & ~t[92] & t[93] & ~t[95]) | (~t[89] & ~t[91] & t[92] & t[93] & t[94]) | (t[92] & t[93] & ~t[94] & ~t[95]);
  assign t[74] = (t[89] & t[90] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[91] & ~t[92] & ~t[93] & t[94]) | (~t[89] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[89] & ~t[90] & ~t[91] & t[94] & ~t[95]) | (~t[90] & t[91] & ~t[92] & t[93] & t[94]) | (t[91] & ~t[93] & t[94] & ~t[95]);
  assign t[75] = (t[89] & t[90] & ~t[91] & t[92] & ~t[93] & ~t[95]) | (t[89] & ~t[91] & ~t[92] & t[93] & ~t[94] & t[95]) | (~t[90] & t[91] & ~t[92] & ~t[93] & ~t[95]) | (~t[89] & t[91] & ~t[92] & ~t[93] & ~t[94]) | (~t[89] & ~t[90] & t[91] & ~t[94] & ~t[95]) | (~t[89] & t[91] & t[92] & ~t[93] & t[94]) | (t[91] & ~t[92] & t[94] & ~t[95]);
  assign t[76] = (t[96] & ~t[98] & ~t[99] & ~t[100] & ~t[101]) | (t[96] & ~t[97] & ~t[99] & ~t[100] & ~t[102]) | (t[96] & ~t[97] & ~t[98] & ~t[101] & ~t[102]) | (~t[96] & t[97] & t[98] & t[99] & ~t[102]) | (~t[96] & t[97] & t[100] & t[101] & ~t[102]) | (t[96] & ~t[98] & ~t[100] & t[102]) | (~t[96] & t[98] & t[100] & t[102]);
  assign t[77] = (t[97] & ~t[98] & ~t[99] & ~t[100] & ~t[101]) | (~t[96] & t[97] & ~t[99] & ~t[100] & ~t[102]) | (~t[96] & t[97] & ~t[98] & ~t[101] & ~t[102]) | (t[96] & ~t[97] & t[98] & t[99] & ~t[102]) | (t[96] & ~t[97] & t[100] & t[101] & ~t[102]) | (t[97] & ~t[99] & ~t[101] & t[102]) | (~t[97] & t[99] & t[101] & t[102]);
  assign t[78] = (t[96] & t[97] & t[98] & ~t[99] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[99] & ~t[100] & t[101] & t[102]) | (~t[97] & ~t[98] & t[99] & ~t[100] & ~t[101]) | (~t[96] & ~t[98] & t[99] & ~t[101] & ~t[102]) | (~t[96] & ~t[97] & t[99] & ~t[100] & ~t[102]) | (~t[97] & t[98] & t[99] & t[100] & ~t[101]) | (~t[98] & t[99] & t[100] & ~t[102]);
  assign t[79] = (t[96] & t[97] & ~t[98] & ~t[100] & t[101] & ~t[102]) | (t[96] & t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[102]) | (~t[96] & ~t[98] & ~t[99] & t[100] & ~t[101]) | (~t[96] & ~t[97] & ~t[99] & t[100] & ~t[102]) | (~t[96] & ~t[98] & t[99] & t[100] & t[101]) | (t[99] & t[100] & ~t[101] & ~t[102]);
  assign t[7] = t[39] ^ t[40];
  assign t[80] = (t[96] & t[97] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[98] & ~t[99] & ~t[100] & t[101]) | (~t[96] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[96] & ~t[97] & ~t[98] & t[101] & ~t[102]) | (~t[97] & t[98] & ~t[99] & t[100] & t[101]) | (t[98] & ~t[100] & t[101] & ~t[102]);
  assign t[81] = (t[96] & t[97] & ~t[98] & t[99] & ~t[100] & ~t[102]) | (t[96] & ~t[98] & ~t[99] & t[100] & ~t[101] & t[102]) | (~t[97] & t[98] & ~t[99] & ~t[100] & ~t[102]) | (~t[96] & t[98] & ~t[99] & ~t[100] & ~t[101]) | (~t[96] & ~t[97] & t[98] & ~t[101] & ~t[102]) | (~t[96] & t[98] & t[99] & ~t[100] & t[101]) | (t[98] & ~t[99] & t[101] & ~t[102]);
  assign t[82] = t[103] ^ x[8];
  assign t[83] = t[104] ^ x[9];
  assign t[84] = t[105] ^ x[6];
  assign t[85] = t[106] ^ x[10];
  assign t[86] = t[107] ^ x[11];
  assign t[87] = t[108] ^ x[12];
  assign t[88] = t[109] ^ x[7];
  assign t[89] = t[110] ^ x[18];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[19];
  assign t[91] = t[112] ^ x[23];
  assign t[92] = t[113] ^ x[20];
  assign t[93] = t[114] ^ x[21];
  assign t[94] = t[115] ^ x[22];
  assign t[95] = t[116] ^ x[17];
  assign t[96] = t[117] ^ x[29];
  assign t[97] = t[118] ^ x[30];
  assign t[98] = t[119] ^ x[34];
  assign t[99] = t[120] ^ x[31];
  assign t[9] = ~t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind105(x, y);
 input [36:0] x;
 output y;

 wire [149:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & t[123] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[123] & ~t[124] & ~t[127] & ~t[128]) | (t[122] & ~t[123] & t[124] & t[125] & ~t[128]) | (t[122] & ~t[123] & t[126] & t[127] & ~t[128]) | (t[123] & ~t[125] & ~t[127] & t[128]) | (~t[123] & t[125] & t[127] & t[128]);
  assign t[101] = (t[122] & t[123] & t[124] & ~t[125] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[125] & ~t[126] & t[127] & t[128]) | (~t[123] & ~t[124] & t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[124] & t[125] & ~t[127] & ~t[128]) | (~t[122] & ~t[123] & t[125] & ~t[126] & ~t[128]) | (~t[123] & t[124] & t[125] & t[126] & ~t[127]) | (~t[124] & t[125] & t[126] & ~t[128]);
  assign t[102] = (t[122] & t[123] & ~t[124] & ~t[126] & t[127] & ~t[128]) | (t[122] & t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[128]) | (~t[122] & ~t[124] & ~t[125] & t[126] & ~t[127]) | (~t[122] & ~t[123] & ~t[125] & t[126] & ~t[128]) | (~t[122] & ~t[124] & t[125] & t[126] & t[127]) | (t[125] & t[126] & ~t[127] & ~t[128]);
  assign t[103] = (t[122] & t[123] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[124] & ~t[125] & ~t[126] & t[127]) | (~t[122] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[122] & ~t[123] & ~t[124] & t[127] & ~t[128]) | (~t[123] & t[124] & ~t[125] & t[126] & t[127]) | (t[124] & ~t[126] & t[127] & ~t[128]);
  assign t[104] = (t[108] & t[109] & ~t[110] & t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[110] & ~t[111] & t[112] & ~t[113] & t[114]) | (~t[109] & t[110] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[109] & t[110] & ~t[113] & ~t[114]) | (~t[108] & t[110] & t[111] & ~t[112] & t[113]) | (t[110] & ~t[111] & t[113] & ~t[114]);
  assign t[105] = (t[109] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (~t[108] & t[109] & ~t[111] & ~t[112] & ~t[114]) | (~t[108] & t[109] & ~t[110] & ~t[113] & ~t[114]) | (t[108] & ~t[109] & t[110] & t[111] & ~t[114]) | (t[108] & ~t[109] & t[112] & t[113] & ~t[114]) | (t[109] & ~t[111] & ~t[113] & t[114]) | (~t[109] & t[111] & t[113] & t[114]);
  assign t[106] = (t[108] & t[109] & t[110] & ~t[111] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & ~t[111] & ~t[112] & t[113] & t[114]) | (~t[109] & ~t[110] & t[111] & ~t[112] & ~t[113]) | (~t[108] & ~t[110] & t[111] & ~t[113] & ~t[114]) | (~t[108] & ~t[109] & t[111] & ~t[112] & ~t[114]) | (~t[109] & t[110] & t[111] & t[112] & ~t[113]) | (~t[110] & t[111] & t[112] & ~t[114]);
  assign t[107] = (t[108] & t[109] & ~t[111] & t[112] & ~t[113] & ~t[114]) | (t[109] & ~t[110] & t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & ~t[111] & ~t[112] & t[113]) | (~t[108] & ~t[111] & ~t[112] & t[113] & ~t[114]) | (~t[108] & ~t[109] & ~t[110] & t[113] & ~t[114]) | (~t[109] & t[110] & ~t[111] & t[112] & t[113]) | (t[110] & ~t[112] & t[113] & ~t[114]);
  assign t[108] = t[129] ^ x[7];
  assign t[109] = t[130] ^ x[34];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[32];
  assign t[111] = t[132] ^ x[35];
  assign t[112] = t[133] ^ x[8];
  assign t[113] = t[134] ^ x[36];
  assign t[114] = t[135] ^ x[6];
  assign t[115] = t[136] ^ x[14];
  assign t[116] = t[137] ^ x[16];
  assign t[117] = t[138] ^ x[15];
  assign t[118] = t[139] ^ x[17];
  assign t[119] = t[140] ^ x[18];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[19];
  assign t[121] = t[142] ^ x[13];
  assign t[122] = t[143] ^ x[25];
  assign t[123] = t[144] ^ x[27];
  assign t[124] = t[145] ^ x[26];
  assign t[125] = t[146] ^ x[28];
  assign t[126] = t[147] ^ x[29];
  assign t[127] = t[148] ^ x[30];
  assign t[128] = t[149] ^ x[24];
  assign t[129] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[131] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[132] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[133] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[134] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[135] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[136] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[137] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[138] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[139] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[141] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[142] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[143] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[144] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[145] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[146] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[147] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[148] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[149] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[63]);
  assign t[15] = ~(t[62] ^ t[14]);
  assign t[16] = t[64] ^ t[63];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[62] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[62] ^ t[27];
  assign t[23] = t[65] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[63] ^ t[66];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[67]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[65] ^ t[29]);
  assign t[31] = t[68] ^ t[67];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[65] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[65] ^ t[36];
  assign t[36] = t[67] ^ t[69];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[70]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[62] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[61]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[65] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[57]);
  assign t[56] = ~(t[58] ^ t[71]);
  assign t[57] = t[27] ^ t[9];
  assign t[58] = ~t[59];
  assign t[59] = ~(t[60]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[36] ^ t[24];
  assign t[61] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[62] = (t[74] & ~t[75]) | (~t[74] & t[75]);
  assign t[63] = (t[74] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[74] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[64] = (t[74] & ~t[78]) | (~t[74] & t[78]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[74] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[74] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[67] = (t[80] & ~t[83] & ~t[85]) | (~t[82] & t[83] & ~t[84]) | (~t[80] & ~t[83] & t[85]) | (t[82] & t[83] & t[84]);
  assign t[68] = (t[80] & ~t[84]) | (~t[80] & t[84]);
  assign t[69] = (t[80] & ~t[83] & ~t[84]) | (~t[82] & t[83] & ~t[85]) | (~t[80] & ~t[83] & t[84]) | (t[82] & t[83] & t[85]);
  assign t[6] = t[10] & t[11];
  assign t[70] = (t[72] & ~t[86]) | (~t[72] & t[86]);
  assign t[71] = (t[72] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[73]) | (~t[72] & ~t[88] & t[89]) | (t[87] & t[88] & t[73]);
  assign t[72] = t[90] ^ x[7];
  assign t[73] = t[91] ^ x[8];
  assign t[74] = t[92] ^ x[14];
  assign t[75] = t[93] ^ x[15];
  assign t[76] = t[94] ^ x[16];
  assign t[77] = t[95] ^ x[17];
  assign t[78] = t[96] ^ x[18];
  assign t[79] = t[97] ^ x[19];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[25];
  assign t[81] = t[99] ^ x[26];
  assign t[82] = t[100] ^ x[27];
  assign t[83] = t[101] ^ x[28];
  assign t[84] = t[102] ^ x[29];
  assign t[85] = t[103] ^ x[30];
  assign t[86] = t[104] ^ x[32];
  assign t[87] = t[105] ^ x[34];
  assign t[88] = t[106] ^ x[35];
  assign t[89] = t[107] ^ x[36];
  assign t[8] = t[62] & t[13];
  assign t[90] = (t[108] & ~t[110] & ~t[111] & ~t[112] & ~t[113]) | (t[108] & ~t[109] & ~t[111] & ~t[112] & ~t[114]) | (t[108] & ~t[109] & ~t[110] & ~t[113] & ~t[114]) | (~t[108] & t[109] & t[110] & t[111] & ~t[114]) | (~t[108] & t[109] & t[112] & t[113] & ~t[114]) | (t[108] & ~t[110] & ~t[112] & t[114]) | (~t[108] & t[110] & t[112] & t[114]);
  assign t[91] = (t[108] & t[109] & ~t[110] & ~t[112] & t[113] & ~t[114]) | (t[108] & t[110] & ~t[111] & ~t[112] & ~t[113] & t[114]) | (~t[109] & ~t[110] & t[112] & ~t[113] & ~t[114]) | (~t[108] & ~t[110] & ~t[111] & t[112] & ~t[113]) | (~t[108] & ~t[109] & ~t[111] & t[112] & ~t[114]) | (~t[108] & ~t[110] & t[111] & t[112] & t[113]) | (t[111] & t[112] & ~t[113] & ~t[114]);
  assign t[92] = (t[115] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (t[115] & ~t[116] & ~t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[116] & ~t[117] & ~t[120] & ~t[121]) | (~t[115] & t[116] & t[117] & t[118] & ~t[121]) | (~t[115] & t[116] & t[119] & t[120] & ~t[121]) | (t[115] & ~t[117] & ~t[119] & t[121]) | (~t[115] & t[117] & t[119] & t[121]);
  assign t[93] = (t[115] & t[116] & ~t[117] & t[118] & ~t[119] & ~t[121]) | (t[115] & ~t[117] & ~t[118] & t[119] & ~t[120] & t[121]) | (~t[116] & t[117] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[116] & t[117] & ~t[120] & ~t[121]) | (~t[115] & t[117] & t[118] & ~t[119] & t[120]) | (t[117] & ~t[118] & t[120] & ~t[121]);
  assign t[94] = (t[116] & ~t[117] & ~t[118] & ~t[119] & ~t[120]) | (~t[115] & t[116] & ~t[118] & ~t[119] & ~t[121]) | (~t[115] & t[116] & ~t[117] & ~t[120] & ~t[121]) | (t[115] & ~t[116] & t[117] & t[118] & ~t[121]) | (t[115] & ~t[116] & t[119] & t[120] & ~t[121]) | (t[116] & ~t[118] & ~t[120] & t[121]) | (~t[116] & t[118] & t[120] & t[121]);
  assign t[95] = (t[115] & t[116] & t[117] & ~t[118] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & ~t[118] & ~t[119] & t[120] & t[121]) | (~t[116] & ~t[117] & t[118] & ~t[119] & ~t[120]) | (~t[115] & ~t[117] & t[118] & ~t[120] & ~t[121]) | (~t[115] & ~t[116] & t[118] & ~t[119] & ~t[121]) | (~t[116] & t[117] & t[118] & t[119] & ~t[120]) | (~t[117] & t[118] & t[119] & ~t[121]);
  assign t[96] = (t[115] & t[116] & ~t[117] & ~t[119] & t[120] & ~t[121]) | (t[115] & t[117] & ~t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & t[119] & ~t[120] & ~t[121]) | (~t[115] & ~t[117] & ~t[118] & t[119] & ~t[120]) | (~t[115] & ~t[116] & ~t[118] & t[119] & ~t[121]) | (~t[115] & ~t[117] & t[118] & t[119] & t[120]) | (t[118] & t[119] & ~t[120] & ~t[121]);
  assign t[97] = (t[115] & t[116] & ~t[118] & t[119] & ~t[120] & ~t[121]) | (t[116] & ~t[117] & t[118] & ~t[119] & ~t[120] & t[121]) | (~t[116] & ~t[117] & ~t[118] & ~t[119] & t[120]) | (~t[115] & ~t[118] & ~t[119] & t[120] & ~t[121]) | (~t[115] & ~t[116] & ~t[117] & t[120] & ~t[121]) | (~t[116] & t[117] & ~t[118] & t[119] & t[120]) | (t[117] & ~t[119] & t[120] & ~t[121]);
  assign t[98] = (t[122] & ~t[124] & ~t[125] & ~t[126] & ~t[127]) | (t[122] & ~t[123] & ~t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[123] & ~t[124] & ~t[127] & ~t[128]) | (~t[122] & t[123] & t[124] & t[125] & ~t[128]) | (~t[122] & t[123] & t[126] & t[127] & ~t[128]) | (t[122] & ~t[124] & ~t[126] & t[128]) | (~t[122] & t[124] & t[126] & t[128]);
  assign t[99] = (t[122] & t[123] & ~t[124] & t[125] & ~t[126] & ~t[128]) | (t[122] & ~t[124] & ~t[125] & t[126] & ~t[127] & t[128]) | (~t[123] & t[124] & ~t[125] & ~t[126] & ~t[128]) | (~t[122] & t[124] & ~t[125] & ~t[126] & ~t[127]) | (~t[122] & ~t[123] & t[124] & ~t[127] & ~t[128]) | (~t[122] & t[124] & t[125] & ~t[126] & t[127]) | (t[124] & ~t[125] & t[127] & ~t[128]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind106(x, y);
 input [36:0] x;
 output y;

 wire [147:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[101] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[102] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[103] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[104] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[105] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[106] = t[127] ^ x[7];
  assign t[107] = t[128] ^ x[34];
  assign t[108] = t[129] ^ x[32];
  assign t[109] = t[130] ^ x[35];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[8];
  assign t[111] = t[132] ^ x[36];
  assign t[112] = t[133] ^ x[6];
  assign t[113] = t[134] ^ x[14];
  assign t[114] = t[135] ^ x[16];
  assign t[115] = t[136] ^ x[15];
  assign t[116] = t[137] ^ x[17];
  assign t[117] = t[138] ^ x[18];
  assign t[118] = t[139] ^ x[19];
  assign t[119] = t[140] ^ x[13];
  assign t[11] = t[17] ^ t[9];
  assign t[120] = t[141] ^ x[25];
  assign t[121] = t[142] ^ x[27];
  assign t[122] = t[143] ^ x[26];
  assign t[123] = t[144] ^ x[28];
  assign t[124] = t[145] ^ x[29];
  assign t[125] = t[146] ^ x[30];
  assign t[126] = t[147] ^ x[24];
  assign t[127] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[128] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[129] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[131] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[132] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[133] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[134] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[135] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[136] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[137] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[138] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[139] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[13] = t[20] ^ t[21];
  assign t[140] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[141] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[142] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[143] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[144] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[145] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[146] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[147] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[14] = ~(t[61]);
  assign t[15] = ~(t[60] ^ t[14]);
  assign t[16] = t[62] ^ t[61];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[60] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[60] ^ t[27];
  assign t[23] = t[63] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[61] ^ t[64];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[65]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[63] ^ t[29]);
  assign t[31] = t[66] ^ t[65];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[63] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[63] ^ t[36];
  assign t[36] = t[65] ^ t[67];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42] ^ t[43]);
  assign t[41] = ~(t[44] ^ t[68]);
  assign t[42] = t[45] ^ t[9];
  assign t[43] = t[5] ^ t[46];
  assign t[44] = ~t[47];
  assign t[45] = t[16] ^ t[21];
  assign t[46] = t[60] ^ t[14];
  assign t[47] = ~(t[48] ^ t[49]);
  assign t[48] = t[50] ^ t[24];
  assign t[49] = t[18] ^ t[51];
  assign t[4] = ~(t[7] ^ t[59]);
  assign t[50] = t[31] ^ t[34];
  assign t[51] = t[63] ^ t[29];
  assign t[52] = x[0] ? x[33] : t[53];
  assign t[53] = ~(t[54] ^ t[55]);
  assign t[54] = ~t[56];
  assign t[55] = ~(t[42]);
  assign t[56] = ~(t[57] ^ t[69]);
  assign t[57] = ~t[58];
  assign t[58] = ~(t[48]);
  assign t[59] = (t[70] & ~t[71]) | (~t[70] & t[71]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = (t[72] & ~t[73]) | (~t[72] & t[73]);
  assign t[61] = (t[72] & ~t[75] & ~t[77]) | (~t[74] & t[75] & ~t[76]) | (~t[72] & ~t[75] & t[77]) | (t[74] & t[75] & t[76]);
  assign t[62] = (t[72] & ~t[76]) | (~t[72] & t[76]);
  assign t[63] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[64] = (t[72] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[77]) | (~t[72] & ~t[75] & t[76]) | (t[74] & t[75] & t[77]);
  assign t[65] = (t[78] & ~t[81] & ~t[83]) | (~t[80] & t[81] & ~t[82]) | (~t[78] & ~t[81] & t[83]) | (t[80] & t[81] & t[82]);
  assign t[66] = (t[78] & ~t[82]) | (~t[78] & t[82]);
  assign t[67] = (t[78] & ~t[81] & ~t[82]) | (~t[80] & t[81] & ~t[83]) | (~t[78] & ~t[81] & t[82]) | (t[80] & t[81] & t[83]);
  assign t[68] = (t[70] & ~t[84]) | (~t[70] & t[84]);
  assign t[69] = (t[70] & ~t[86] & ~t[71]) | (~t[85] & t[86] & ~t[87]) | (~t[70] & ~t[86] & t[71]) | (t[85] & t[86] & t[87]);
  assign t[6] = t[10] & t[11];
  assign t[70] = t[88] ^ x[7];
  assign t[71] = t[89] ^ x[8];
  assign t[72] = t[90] ^ x[14];
  assign t[73] = t[91] ^ x[15];
  assign t[74] = t[92] ^ x[16];
  assign t[75] = t[93] ^ x[17];
  assign t[76] = t[94] ^ x[18];
  assign t[77] = t[95] ^ x[19];
  assign t[78] = t[96] ^ x[25];
  assign t[79] = t[97] ^ x[26];
  assign t[7] = ~t[12];
  assign t[80] = t[98] ^ x[27];
  assign t[81] = t[99] ^ x[28];
  assign t[82] = t[100] ^ x[29];
  assign t[83] = t[101] ^ x[30];
  assign t[84] = t[102] ^ x[32];
  assign t[85] = t[103] ^ x[34];
  assign t[86] = t[104] ^ x[35];
  assign t[87] = t[105] ^ x[36];
  assign t[88] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[89] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[8] = t[60] & t[13];
  assign t[90] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[92] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[93] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[94] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[95] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[96] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[97] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[98] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[99] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37] & ~t[52]) | (~t[0] & t[37] & ~t[52]) | (~t[0] & ~t[37] & t[52]) | (t[0] & t[37] & t[52]);
endmodule

module R2ind107(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[19];
  assign t[102] = t[123] ^ x[20];
  assign t[103] = t[124] ^ x[14];
  assign t[104] = t[125] ^ x[26];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[27];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[30];
  assign t[109] = t[130] ^ x[31];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[25];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[119] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[121] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[122] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[123] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[124] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[125] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[126] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[127] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[128] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[129] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[131] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[48]);
  assign t[15] = ~(t[47] ^ t[14]);
  assign t[16] = t[49] ^ t[48];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[47] ^ t[27];
  assign t[23] = t[50] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[48] ^ t[51];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[52]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[50] ^ t[29]);
  assign t[31] = t[53] ^ t[52];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[50] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[50] ^ t[36];
  assign t[36] = t[52] ^ t[54];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[27] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[36] ^ t[24];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[61] & ~t[63]) | (~t[60] & t[61] & ~t[62]) | (~t[58] & ~t[61] & t[63]) | (t[60] & t[61] & t[62]);
  assign t[49] = (t[58] & ~t[62]) | (~t[58] & t[62]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[61] & ~t[62]) | (~t[60] & t[61] & ~t[63]) | (~t[58] & ~t[61] & t[62]) | (t[60] & t[61] & t[63]);
  assign t[52] = (t[64] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[64] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[53] = (t[64] & ~t[68]) | (~t[64] & t[68]);
  assign t[54] = (t[64] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[64] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[72]) | (~t[70] & t[71] & ~t[57]) | (~t[56] & ~t[71] & t[72]) | (t[70] & t[71] & t[57]);
  assign t[56] = t[73] ^ x[8];
  assign t[57] = t[74] ^ x[9];
  assign t[58] = t[75] ^ x[15];
  assign t[59] = t[76] ^ x[16];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[17];
  assign t[61] = t[78] ^ x[18];
  assign t[62] = t[79] ^ x[19];
  assign t[63] = t[80] ^ x[20];
  assign t[64] = t[81] ^ x[26];
  assign t[65] = t[82] ^ x[27];
  assign t[66] = t[83] ^ x[28];
  assign t[67] = t[84] ^ x[29];
  assign t[68] = t[85] ^ x[30];
  assign t[69] = t[86] ^ x[31];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[33];
  assign t[71] = t[88] ^ x[34];
  assign t[72] = t[89] ^ x[35];
  assign t[73] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[74] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[75] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[86] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[87] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[88] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[47] & t[13];
  assign t[90] = t[111] ^ x[8];
  assign t[91] = t[112] ^ x[33];
  assign t[92] = t[113] ^ x[6];
  assign t[93] = t[114] ^ x[34];
  assign t[94] = t[115] ^ x[9];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[7];
  assign t[97] = t[118] ^ x[15];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[16];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind108(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[19];
  assign t[104] = t[125] ^ x[20];
  assign t[105] = t[126] ^ x[14];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[16] ^ t[14];
  assign t[110] = t[131] ^ x[30];
  assign t[111] = t[132] ^ x[31];
  assign t[112] = t[133] ^ x[25];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[17] ^ t[9];
  assign t[120] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[121] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[122] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[123] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[126] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[127] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[128] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[129] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[12] = t[18] ^ t[19];
  assign t[130] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[132] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[133] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[13] = t[20] ^ t[21];
  assign t[14] = ~(t[50]);
  assign t[15] = ~(t[49] ^ t[14]);
  assign t[16] = t[51] ^ t[50];
  assign t[17] = ~(t[22] ^ t[10]);
  assign t[18] = t[23] ^ t[24];
  assign t[19] = t[25] & t[26];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[49] ^ t[16];
  assign t[21] = t[14] & t[22];
  assign t[22] = t[49] ^ t[27];
  assign t[23] = t[52] & t[28];
  assign t[24] = t[29] & t[30];
  assign t[25] = t[31] ^ t[29];
  assign t[26] = t[32] ^ t[24];
  assign t[27] = t[50] ^ t[53];
  assign t[28] = t[33] ^ t[34];
  assign t[29] = ~(t[54]);
  assign t[2] = ~t[4];
  assign t[30] = ~(t[52] ^ t[29]);
  assign t[31] = t[55] ^ t[54];
  assign t[32] = ~(t[35] ^ t[25]);
  assign t[33] = t[52] ^ t[31];
  assign t[34] = t[29] & t[35];
  assign t[35] = t[52] ^ t[36];
  assign t[36] = t[54] ^ t[56];
  assign t[37] = x[0] ? x[32] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = t[5] ^ t[6];
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[57]);
  assign t[42] = t[44] ^ t[9];
  assign t[43] = ~t[45];
  assign t[44] = t[16] ^ t[21];
  assign t[45] = ~(t[46]);
  assign t[46] = t[47] ^ t[24];
  assign t[47] = t[31] ^ t[34];
  assign t[48] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[49] = (t[60] & ~t[61]) | (~t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[48]);
  assign t[50] = (t[60] & ~t[63] & ~t[65]) | (~t[62] & t[63] & ~t[64]) | (~t[60] & ~t[63] & t[65]) | (t[62] & t[63] & t[64]);
  assign t[51] = (t[60] & ~t[64]) | (~t[60] & t[64]);
  assign t[52] = (t[66] & ~t[67]) | (~t[66] & t[67]);
  assign t[53] = (t[60] & ~t[63] & ~t[64]) | (~t[62] & t[63] & ~t[65]) | (~t[60] & ~t[63] & t[64]) | (t[62] & t[63] & t[65]);
  assign t[54] = (t[66] & ~t[69] & ~t[71]) | (~t[68] & t[69] & ~t[70]) | (~t[66] & ~t[69] & t[71]) | (t[68] & t[69] & t[70]);
  assign t[55] = (t[66] & ~t[70]) | (~t[66] & t[70]);
  assign t[56] = (t[66] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[66] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[57] = (t[58] & ~t[73] & ~t[59]) | (~t[72] & t[73] & ~t[74]) | (~t[58] & ~t[73] & t[59]) | (t[72] & t[73] & t[74]);
  assign t[58] = t[75] ^ x[8];
  assign t[59] = t[76] ^ x[9];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[77] ^ x[15];
  assign t[61] = t[78] ^ x[16];
  assign t[62] = t[79] ^ x[17];
  assign t[63] = t[80] ^ x[18];
  assign t[64] = t[81] ^ x[19];
  assign t[65] = t[82] ^ x[20];
  assign t[66] = t[83] ^ x[26];
  assign t[67] = t[84] ^ x[27];
  assign t[68] = t[85] ^ x[28];
  assign t[69] = t[86] ^ x[29];
  assign t[6] = t[10] & t[11];
  assign t[70] = t[87] ^ x[30];
  assign t[71] = t[88] ^ x[31];
  assign t[72] = t[89] ^ x[33];
  assign t[73] = t[90] ^ x[34];
  assign t[74] = t[91] ^ x[35];
  assign t[75] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[76] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[77] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[82] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[88] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[89] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[8] = t[49] & t[13];
  assign t[90] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[6];
  assign t[95] = t[116] ^ x[34];
  assign t[96] = t[117] ^ x[9];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[7];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind109(x, y);
 input [35:0] x;
 output y;

 wire [133:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[17];
  assign t[101] = t[122] ^ x[15];
  assign t[102] = t[123] ^ x[18];
  assign t[103] = t[124] ^ x[16];
  assign t[104] = t[125] ^ x[19];
  assign t[105] = t[126] ^ x[13];
  assign t[106] = t[127] ^ x[25];
  assign t[107] = t[128] ^ x[28];
  assign t[108] = t[129] ^ x[26];
  assign t[109] = t[130] ^ x[29];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[27];
  assign t[111] = t[132] ^ x[30];
  assign t[112] = t[133] ^ x[24];
  assign t[113] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[114] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[115] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[116] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[117] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[118] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[119] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[11] = t[47] ^ t[15];
  assign t[120] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[121] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[122] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[123] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[124] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[125] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[126] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[127] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[128] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[129] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[131] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[132] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[133] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[48] ^ t[49];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[49]);
  assign t[16] = ~(t[47] ^ t[15]);
  assign t[17] = t[47] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[47] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[50] ^ t[30];
  assign t[26] = t[49] ^ t[51];
  assign t[27] = t[47] ^ t[13];
  assign t[28] = t[52] ^ t[53];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[53]);
  assign t[31] = ~(t[50] ^ t[30]);
  assign t[32] = t[50] & t[34];
  assign t[33] = t[50] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[53] ^ t[54];
  assign t[36] = t[50] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[42]);
  assign t[41] = ~(t[43] ^ t[55]);
  assign t[42] = t[26] ^ t[9];
  assign t[43] = ~t[44];
  assign t[44] = ~(t[45]);
  assign t[45] = t[35] ^ t[23];
  assign t[46] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[47] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[48] = (t[58] & ~t[60]) | (~t[58] & t[60]);
  assign t[49] = (t[58] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[60]) | (~t[58] & ~t[62] & t[63]) | (t[61] & t[62] & t[60]);
  assign t[4] = ~(t[7] ^ t[46]);
  assign t[50] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[51] = (t[58] & ~t[62] & ~t[60]) | (~t[61] & t[62] & ~t[63]) | (~t[58] & ~t[62] & t[60]) | (t[61] & t[62] & t[63]);
  assign t[52] = (t[64] & ~t[66]) | (~t[64] & t[66]);
  assign t[53] = (t[64] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[66]) | (~t[64] & ~t[68] & t[69]) | (t[67] & t[68] & t[66]);
  assign t[54] = (t[64] & ~t[68] & ~t[66]) | (~t[67] & t[68] & ~t[69]) | (~t[64] & ~t[68] & t[66]) | (t[67] & t[68] & t[69]);
  assign t[55] = (t[56] & ~t[71] & ~t[73]) | (~t[70] & t[71] & ~t[72]) | (~t[56] & ~t[71] & t[73]) | (t[70] & t[71] & t[72]);
  assign t[56] = t[74] ^ x[7];
  assign t[57] = t[75] ^ x[8];
  assign t[58] = t[76] ^ x[14];
  assign t[59] = t[77] ^ x[15];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[16];
  assign t[61] = t[79] ^ x[17];
  assign t[62] = t[80] ^ x[18];
  assign t[63] = t[81] ^ x[19];
  assign t[64] = t[82] ^ x[25];
  assign t[65] = t[83] ^ x[26];
  assign t[66] = t[84] ^ x[27];
  assign t[67] = t[85] ^ x[28];
  assign t[68] = t[86] ^ x[29];
  assign t[69] = t[87] ^ x[30];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[32];
  assign t[71] = t[89] ^ x[33];
  assign t[72] = t[90] ^ x[34];
  assign t[73] = t[91] ^ x[35];
  assign t[74] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[76] = (t[99] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[100] & ~t[101] & ~t[104] & ~t[105]) | (~t[99] & t[100] & t[101] & t[102] & ~t[105]) | (~t[99] & t[100] & t[103] & t[104] & ~t[105]) | (t[99] & ~t[101] & ~t[103] & t[105]) | (~t[99] & t[101] & t[103] & t[105]);
  assign t[77] = (t[99] & t[100] & ~t[101] & t[102] & ~t[103] & ~t[105]) | (t[99] & ~t[101] & ~t[102] & t[103] & ~t[104] & t[105]) | (~t[100] & t[101] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[100] & t[101] & ~t[104] & ~t[105]) | (~t[99] & t[101] & t[102] & ~t[103] & t[104]) | (t[101] & ~t[102] & t[104] & ~t[105]);
  assign t[78] = (t[99] & t[100] & ~t[101] & ~t[103] & t[104] & ~t[105]) | (t[99] & t[101] & ~t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & t[103] & ~t[104] & ~t[105]) | (~t[99] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[99] & ~t[100] & ~t[102] & t[103] & ~t[105]) | (~t[99] & ~t[101] & t[102] & t[103] & t[104]) | (t[102] & t[103] & ~t[104] & ~t[105]);
  assign t[79] = (t[100] & ~t[101] & ~t[102] & ~t[103] & ~t[104]) | (~t[99] & t[100] & ~t[102] & ~t[103] & ~t[105]) | (~t[99] & t[100] & ~t[101] & ~t[104] & ~t[105]) | (t[99] & ~t[100] & t[101] & t[102] & ~t[105]) | (t[99] & ~t[100] & t[103] & t[104] & ~t[105]) | (t[100] & ~t[102] & ~t[104] & t[105]) | (~t[100] & t[102] & t[104] & t[105]);
  assign t[7] = ~t[12];
  assign t[80] = (t[99] & t[100] & t[101] & ~t[102] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & ~t[102] & ~t[103] & t[104] & t[105]) | (~t[100] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (~t[99] & ~t[101] & t[102] & ~t[104] & ~t[105]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[105]) | (~t[100] & t[101] & t[102] & t[103] & ~t[104]) | (~t[101] & t[102] & t[103] & ~t[105]);
  assign t[81] = (t[99] & t[100] & ~t[102] & t[103] & ~t[104] & ~t[105]) | (t[100] & ~t[101] & t[102] & ~t[103] & ~t[104] & t[105]) | (~t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[102] & ~t[103] & t[104] & ~t[105]) | (~t[99] & ~t[100] & ~t[101] & t[104] & ~t[105]) | (~t[100] & t[101] & ~t[102] & t[103] & t[104]) | (t[101] & ~t[103] & t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[83] = (t[106] & t[107] & ~t[108] & t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[108] & ~t[109] & t[110] & ~t[111] & t[112]) | (~t[107] & t[108] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[107] & t[108] & ~t[111] & ~t[112]) | (~t[106] & t[108] & t[109] & ~t[110] & t[111]) | (t[108] & ~t[109] & t[111] & ~t[112]);
  assign t[84] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[85] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[86] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[89] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[91] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[92] = t[113] ^ x[7];
  assign t[93] = t[114] ^ x[32];
  assign t[94] = t[115] ^ x[8];
  assign t[95] = t[116] ^ x[33];
  assign t[96] = t[117] ^ x[34];
  assign t[97] = t[118] ^ x[35];
  assign t[98] = t[119] ^ x[6];
  assign t[99] = t[120] ^ x[14];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind110(x, y);
 input [35:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[121] ^ x[18];
  assign t[101] = t[122] ^ x[16];
  assign t[102] = t[123] ^ x[19];
  assign t[103] = t[124] ^ x[13];
  assign t[104] = t[125] ^ x[25];
  assign t[105] = t[126] ^ x[28];
  assign t[106] = t[127] ^ x[26];
  assign t[107] = t[128] ^ x[29];
  assign t[108] = t[129] ^ x[27];
  assign t[109] = t[130] ^ x[30];
  assign t[10] = t[17] ^ t[9];
  assign t[110] = t[131] ^ x[24];
  assign t[111] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[112] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[113] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[114] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[115] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[116] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[117] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[118] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[119] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[11] = t[45] ^ t[15];
  assign t[120] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[121] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[122] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[123] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[124] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[125] = (x[20] & ~x[21] & ~x[22]) | (~x[20] & x[21] & ~x[22]) | (~x[20] & ~x[21] & x[22]) | (x[20] & x[21] & x[22]);
  assign t[126] = (x[20] & ~x[21] & ~x[23]) | (~x[20] & x[21] & ~x[23]) | (~x[20] & ~x[21] & x[23]) | (x[20] & x[21] & x[23]);
  assign t[127] = (x[20] & ~x[22]) | (~x[20] & x[22]);
  assign t[128] = (x[20] & ~x[23]) | (~x[20] & x[23]);
  assign t[129] = (x[21] & ~x[22]) | (~x[21] & x[22]);
  assign t[12] = ~(t[18] ^ t[19]);
  assign t[130] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[131] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[13] = t[46] ^ t[47];
  assign t[14] = t[15] & t[20];
  assign t[15] = ~(t[47]);
  assign t[16] = ~(t[45] ^ t[15]);
  assign t[17] = t[45] & t[21];
  assign t[18] = t[22] ^ t[23];
  assign t[19] = t[24] ^ t[25];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[45] ^ t[26];
  assign t[21] = t[27] ^ t[14];
  assign t[22] = t[28] ^ t[29];
  assign t[23] = t[30] & t[31];
  assign t[24] = t[32] ^ t[23];
  assign t[25] = t[48] ^ t[30];
  assign t[26] = t[47] ^ t[49];
  assign t[27] = t[45] ^ t[13];
  assign t[28] = t[50] ^ t[51];
  assign t[29] = t[30] & t[33];
  assign t[2] = ~t[4];
  assign t[30] = ~(t[51]);
  assign t[31] = ~(t[48] ^ t[30]);
  assign t[32] = t[48] & t[34];
  assign t[33] = t[48] ^ t[35];
  assign t[34] = t[36] ^ t[29];
  assign t[35] = t[51] ^ t[52];
  assign t[36] = t[48] ^ t[28];
  assign t[37] = x[0] ? x[31] : t[38];
  assign t[38] = ~(t[39] ^ t[40]);
  assign t[39] = ~t[41];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[5]);
  assign t[41] = ~(t[42] ^ t[53]);
  assign t[42] = ~t[43];
  assign t[43] = ~(t[18]);
  assign t[44] = (t[54] & ~t[55]) | (~t[54] & t[55]);
  assign t[45] = (t[56] & ~t[57]) | (~t[56] & t[57]);
  assign t[46] = (t[56] & ~t[58]) | (~t[56] & t[58]);
  assign t[47] = (t[56] & ~t[60] & ~t[61]) | (~t[59] & t[60] & ~t[58]) | (~t[56] & ~t[60] & t[61]) | (t[59] & t[60] & t[58]);
  assign t[48] = (t[62] & ~t[63]) | (~t[62] & t[63]);
  assign t[49] = (t[56] & ~t[60] & ~t[58]) | (~t[59] & t[60] & ~t[61]) | (~t[56] & ~t[60] & t[58]) | (t[59] & t[60] & t[61]);
  assign t[4] = ~(t[7] ^ t[44]);
  assign t[50] = (t[62] & ~t[64]) | (~t[62] & t[64]);
  assign t[51] = (t[62] & ~t[66] & ~t[67]) | (~t[65] & t[66] & ~t[64]) | (~t[62] & ~t[66] & t[67]) | (t[65] & t[66] & t[64]);
  assign t[52] = (t[62] & ~t[66] & ~t[64]) | (~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[66] & t[64]) | (t[65] & t[66] & t[67]);
  assign t[53] = (t[54] & ~t[69] & ~t[70]) | (~t[68] & t[69] & ~t[71]) | (~t[54] & ~t[69] & t[70]) | (t[68] & t[69] & t[71]);
  assign t[54] = t[72] ^ x[7];
  assign t[55] = t[73] ^ x[8];
  assign t[56] = t[74] ^ x[14];
  assign t[57] = t[75] ^ x[15];
  assign t[58] = t[76] ^ x[16];
  assign t[59] = t[77] ^ x[17];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[78] ^ x[18];
  assign t[61] = t[79] ^ x[19];
  assign t[62] = t[80] ^ x[25];
  assign t[63] = t[81] ^ x[26];
  assign t[64] = t[82] ^ x[27];
  assign t[65] = t[83] ^ x[28];
  assign t[66] = t[84] ^ x[29];
  assign t[67] = t[85] ^ x[30];
  assign t[68] = t[86] ^ x[32];
  assign t[69] = t[87] ^ x[33];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[88] ^ x[34];
  assign t[71] = t[89] ^ x[35];
  assign t[72] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[73] = (t[90] & t[91] & ~t[92] & t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[92] & ~t[93] & t[94] & ~t[95] & t[96]) | (~t[91] & t[92] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[91] & t[92] & ~t[95] & ~t[96]) | (~t[90] & t[92] & t[93] & ~t[94] & t[95]) | (t[92] & ~t[93] & t[95] & ~t[96]);
  assign t[74] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[75] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[76] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[77] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[78] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[79] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[7] = ~t[12];
  assign t[80] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[81] = (t[104] & t[105] & ~t[106] & t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[106] & ~t[107] & t[108] & ~t[109] & t[110]) | (~t[105] & t[106] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[105] & t[106] & ~t[109] & ~t[110]) | (~t[104] & t[106] & t[107] & ~t[108] & t[109]) | (t[106] & ~t[107] & t[109] & ~t[110]);
  assign t[82] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[83] = (t[105] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (~t[104] & t[105] & ~t[107] & ~t[108] & ~t[110]) | (~t[104] & t[105] & ~t[106] & ~t[109] & ~t[110]) | (t[104] & ~t[105] & t[106] & t[107] & ~t[110]) | (t[104] & ~t[105] & t[108] & t[109] & ~t[110]) | (t[105] & ~t[107] & ~t[109] & t[110]) | (~t[105] & t[107] & t[109] & t[110]);
  assign t[84] = (t[104] & t[105] & t[106] & ~t[107] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[107] & ~t[108] & t[109] & t[110]) | (~t[105] & ~t[106] & t[107] & ~t[108] & ~t[109]) | (~t[104] & ~t[106] & t[107] & ~t[109] & ~t[110]) | (~t[104] & ~t[105] & t[107] & ~t[108] & ~t[110]) | (~t[105] & t[106] & t[107] & t[108] & ~t[109]) | (~t[106] & t[107] & t[108] & ~t[110]);
  assign t[85] = (t[104] & t[105] & ~t[107] & t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & ~t[107] & ~t[108] & t[109]) | (~t[104] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[104] & ~t[105] & ~t[106] & t[109] & ~t[110]) | (~t[105] & t[106] & ~t[107] & t[108] & t[109]) | (t[106] & ~t[108] & t[109] & ~t[110]);
  assign t[86] = (t[91] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (~t[90] & t[91] & ~t[93] & ~t[94] & ~t[96]) | (~t[90] & t[91] & ~t[92] & ~t[95] & ~t[96]) | (t[90] & ~t[91] & t[92] & t[93] & ~t[96]) | (t[90] & ~t[91] & t[94] & t[95] & ~t[96]) | (t[91] & ~t[93] & ~t[95] & t[96]) | (~t[91] & t[93] & t[95] & t[96]);
  assign t[87] = (t[90] & t[91] & t[92] & ~t[93] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[93] & ~t[94] & t[95] & t[96]) | (~t[91] & ~t[92] & t[93] & ~t[94] & ~t[95]) | (~t[90] & ~t[92] & t[93] & ~t[95] & ~t[96]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[96]) | (~t[91] & t[92] & t[93] & t[94] & ~t[95]) | (~t[92] & t[93] & t[94] & ~t[96]);
  assign t[88] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[89] = (t[90] & t[91] & ~t[93] & t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[90] & ~t[91] & ~t[92] & t[95] & ~t[96]) | (~t[91] & t[92] & ~t[93] & t[94] & t[95]) | (t[92] & ~t[94] & t[95] & ~t[96]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[111] ^ x[7];
  assign t[91] = t[112] ^ x[32];
  assign t[92] = t[113] ^ x[8];
  assign t[93] = t[114] ^ x[33];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[35];
  assign t[96] = t[117] ^ x[6];
  assign t[97] = t[118] ^ x[14];
  assign t[98] = t[119] ^ x[17];
  assign t[99] = t[120] ^ x[15];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[37]) | (~t[0] & t[37]);
endmodule

module R2ind111(x, y);
 input [35:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[101] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[102] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[103] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[104] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[105] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[106] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[107] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[108] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[109] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[10] = ~(t[35]);
  assign t[110] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[111] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[112] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[113] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[114] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[115] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[116] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[117] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[118] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[119] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[11] = ~(t[37] ^ t[10]);
  assign t[12] = t[13] ^ t[14];
  assign t[13] = t[38] ^ t[39];
  assign t[14] = t[15] & t[16];
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[40] ^ t[15]);
  assign t[17] = x[0] ? x[35] : t[18];
  assign t[18] = ~(t[19] ^ t[20]);
  assign t[19] = ~t[21];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[22]);
  assign t[21] = ~(t[23] ^ t[41]);
  assign t[22] = t[24] ^ t[8];
  assign t[23] = ~t[25];
  assign t[24] = t[26] ^ t[27];
  assign t[25] = ~(t[28]);
  assign t[26] = t[42] ^ t[35];
  assign t[27] = t[10] & t[29];
  assign t[28] = t[30] ^ t[14];
  assign t[29] = t[37] ^ t[7];
  assign t[2] = ~t[4];
  assign t[30] = t[31] ^ t[32];
  assign t[31] = t[43] ^ t[38];
  assign t[32] = t[15] & t[33];
  assign t[33] = t[40] ^ t[13];
  assign t[34] = (t[44] & ~t[46] & ~t[48]) | (~t[45] & t[46] & ~t[47]) | (~t[44] & ~t[46] & t[48]) | (t[45] & t[46] & t[47]);
  assign t[35] = (t[49] & ~t[51] & ~t[53]) | (~t[50] & t[51] & ~t[52]) | (~t[49] & ~t[51] & t[53]) | (t[50] & t[51] & t[52]);
  assign t[36] = (t[49] & ~t[51] & ~t[52]) | (~t[50] & t[51] & ~t[53]) | (~t[49] & ~t[51] & t[52]) | (t[50] & t[51] & t[53]);
  assign t[37] = (t[49] & ~t[54]) | (~t[49] & t[54]);
  assign t[38] = (t[55] & ~t[57] & ~t[59]) | (~t[56] & t[57] & ~t[58]) | (~t[55] & ~t[57] & t[59]) | (t[56] & t[57] & t[58]);
  assign t[39] = (t[55] & ~t[57] & ~t[58]) | (~t[56] & t[57] & ~t[59]) | (~t[55] & ~t[57] & t[58]) | (t[56] & t[57] & t[59]);
  assign t[3] = ~(t[5]);
  assign t[40] = (t[55] & ~t[60]) | (~t[55] & t[60]);
  assign t[41] = (t[44] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[44] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[42] = (t[49] & ~t[52]) | (~t[49] & t[52]);
  assign t[43] = (t[55] & ~t[58]) | (~t[55] & t[58]);
  assign t[44] = t[61] ^ x[8];
  assign t[45] = t[62] ^ x[9];
  assign t[46] = t[63] ^ x[10];
  assign t[47] = t[64] ^ x[11];
  assign t[48] = t[65] ^ x[12];
  assign t[49] = t[66] ^ x[18];
  assign t[4] = ~(t[6] ^ t[34]);
  assign t[50] = t[67] ^ x[19];
  assign t[51] = t[68] ^ x[20];
  assign t[52] = t[69] ^ x[21];
  assign t[53] = t[70] ^ x[22];
  assign t[54] = t[71] ^ x[23];
  assign t[55] = t[72] ^ x[29];
  assign t[56] = t[73] ^ x[30];
  assign t[57] = t[74] ^ x[31];
  assign t[58] = t[75] ^ x[32];
  assign t[59] = t[76] ^ x[33];
  assign t[5] = t[7] ^ t[8];
  assign t[60] = t[77] ^ x[34];
  assign t[61] = (t[78] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (t[78] & ~t[79] & ~t[81] & ~t[82] & ~t[84]) | (t[78] & ~t[79] & ~t[80] & ~t[83] & ~t[84]) | (~t[78] & t[79] & t[80] & t[81] & ~t[84]) | (~t[78] & t[79] & t[82] & t[83] & ~t[84]) | (t[78] & ~t[80] & ~t[82] & t[84]) | (~t[78] & t[80] & t[82] & t[84]);
  assign t[62] = (t[79] & ~t[80] & ~t[81] & ~t[82] & ~t[83]) | (~t[78] & t[79] & ~t[81] & ~t[82] & ~t[84]) | (~t[78] & t[79] & ~t[80] & ~t[83] & ~t[84]) | (t[78] & ~t[79] & t[80] & t[81] & ~t[84]) | (t[78] & ~t[79] & t[82] & t[83] & ~t[84]) | (t[79] & ~t[81] & ~t[83] & t[84]) | (~t[79] & t[81] & t[83] & t[84]);
  assign t[63] = (t[78] & t[79] & t[80] & ~t[81] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & ~t[81] & ~t[82] & t[83] & t[84]) | (~t[79] & ~t[80] & t[81] & ~t[82] & ~t[83]) | (~t[78] & ~t[80] & t[81] & ~t[83] & ~t[84]) | (~t[78] & ~t[79] & t[81] & ~t[82] & ~t[84]) | (~t[79] & t[80] & t[81] & t[82] & ~t[83]) | (~t[80] & t[81] & t[82] & ~t[84]);
  assign t[64] = (t[78] & t[79] & ~t[80] & ~t[82] & t[83] & ~t[84]) | (t[78] & t[80] & ~t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & t[82] & ~t[83] & ~t[84]) | (~t[78] & ~t[80] & ~t[81] & t[82] & ~t[83]) | (~t[78] & ~t[79] & ~t[81] & t[82] & ~t[84]) | (~t[78] & ~t[80] & t[81] & t[82] & t[83]) | (t[81] & t[82] & ~t[83] & ~t[84]);
  assign t[65] = (t[78] & t[79] & ~t[81] & t[82] & ~t[83] & ~t[84]) | (t[79] & ~t[80] & t[81] & ~t[82] & ~t[83] & t[84]) | (~t[79] & ~t[80] & ~t[81] & ~t[82] & t[83]) | (~t[78] & ~t[81] & ~t[82] & t[83] & ~t[84]) | (~t[78] & ~t[79] & ~t[80] & t[83] & ~t[84]) | (~t[79] & t[80] & ~t[81] & t[82] & t[83]) | (t[80] & ~t[82] & t[83] & ~t[84]);
  assign t[66] = (t[85] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[86] & ~t[87] & ~t[90] & ~t[91]) | (~t[85] & t[86] & t[87] & t[88] & ~t[91]) | (~t[85] & t[86] & t[89] & t[90] & ~t[91]) | (t[85] & ~t[87] & ~t[89] & t[91]) | (~t[85] & t[87] & t[89] & t[91]);
  assign t[67] = (t[86] & ~t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & t[86] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[86] & ~t[87] & ~t[90] & ~t[91]) | (t[85] & ~t[86] & t[87] & t[88] & ~t[91]) | (t[85] & ~t[86] & t[89] & t[90] & ~t[91]) | (t[86] & ~t[88] & ~t[90] & t[91]) | (~t[86] & t[88] & t[90] & t[91]);
  assign t[68] = (t[85] & t[86] & t[87] & ~t[88] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & ~t[88] & ~t[89] & t[90] & t[91]) | (~t[86] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[87] & t[88] & ~t[90] & ~t[91]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[91]) | (~t[86] & t[87] & t[88] & t[89] & ~t[90]) | (~t[87] & t[88] & t[89] & ~t[91]);
  assign t[69] = (t[85] & t[86] & ~t[87] & ~t[89] & t[90] & ~t[91]) | (t[85] & t[87] & ~t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & t[89] & ~t[90] & ~t[91]) | (~t[85] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[85] & ~t[86] & ~t[88] & t[89] & ~t[91]) | (~t[85] & ~t[87] & t[88] & t[89] & t[90]) | (t[88] & t[89] & ~t[90] & ~t[91]);
  assign t[6] = ~t[9];
  assign t[70] = (t[85] & t[86] & ~t[88] & t[89] & ~t[90] & ~t[91]) | (t[86] & ~t[87] & t[88] & ~t[89] & ~t[90] & t[91]) | (~t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[88] & ~t[89] & t[90] & ~t[91]) | (~t[85] & ~t[86] & ~t[87] & t[90] & ~t[91]) | (~t[86] & t[87] & ~t[88] & t[89] & t[90]) | (t[87] & ~t[89] & t[90] & ~t[91]);
  assign t[71] = (t[85] & t[86] & ~t[87] & t[88] & ~t[89] & ~t[91]) | (t[85] & ~t[87] & ~t[88] & t[89] & ~t[90] & t[91]) | (~t[86] & t[87] & ~t[88] & ~t[89] & ~t[91]) | (~t[85] & t[87] & ~t[88] & ~t[89] & ~t[90]) | (~t[85] & ~t[86] & t[87] & ~t[90] & ~t[91]) | (~t[85] & t[87] & t[88] & ~t[89] & t[90]) | (t[87] & ~t[88] & t[90] & ~t[91]);
  assign t[72] = (t[92] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (t[92] & ~t[93] & ~t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[93] & ~t[94] & ~t[97] & ~t[98]) | (~t[92] & t[93] & t[94] & t[95] & ~t[98]) | (~t[92] & t[93] & t[96] & t[97] & ~t[98]) | (t[92] & ~t[94] & ~t[96] & t[98]) | (~t[92] & t[94] & t[96] & t[98]);
  assign t[73] = (t[93] & ~t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & t[93] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[93] & ~t[94] & ~t[97] & ~t[98]) | (t[92] & ~t[93] & t[94] & t[95] & ~t[98]) | (t[92] & ~t[93] & t[96] & t[97] & ~t[98]) | (t[93] & ~t[95] & ~t[97] & t[98]) | (~t[93] & t[95] & t[97] & t[98]);
  assign t[74] = (t[92] & t[93] & t[94] & ~t[95] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & ~t[95] & ~t[96] & t[97] & t[98]) | (~t[93] & ~t[94] & t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[94] & t[95] & ~t[97] & ~t[98]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[98]) | (~t[93] & t[94] & t[95] & t[96] & ~t[97]) | (~t[94] & t[95] & t[96] & ~t[98]);
  assign t[75] = (t[92] & t[93] & ~t[94] & ~t[96] & t[97] & ~t[98]) | (t[92] & t[94] & ~t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & t[96] & ~t[97] & ~t[98]) | (~t[92] & ~t[94] & ~t[95] & t[96] & ~t[97]) | (~t[92] & ~t[93] & ~t[95] & t[96] & ~t[98]) | (~t[92] & ~t[94] & t[95] & t[96] & t[97]) | (t[95] & t[96] & ~t[97] & ~t[98]);
  assign t[76] = (t[92] & t[93] & ~t[95] & t[96] & ~t[97] & ~t[98]) | (t[93] & ~t[94] & t[95] & ~t[96] & ~t[97] & t[98]) | (~t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[95] & ~t[96] & t[97] & ~t[98]) | (~t[92] & ~t[93] & ~t[94] & t[97] & ~t[98]) | (~t[93] & t[94] & ~t[95] & t[96] & t[97]) | (t[94] & ~t[96] & t[97] & ~t[98]);
  assign t[77] = (t[92] & t[93] & ~t[94] & t[95] & ~t[96] & ~t[98]) | (t[92] & ~t[94] & ~t[95] & t[96] & ~t[97] & t[98]) | (~t[93] & t[94] & ~t[95] & ~t[96] & ~t[98]) | (~t[92] & t[94] & ~t[95] & ~t[96] & ~t[97]) | (~t[92] & ~t[93] & t[94] & ~t[97] & ~t[98]) | (~t[92] & t[94] & t[95] & ~t[96] & t[97]) | (t[94] & ~t[95] & t[97] & ~t[98]);
  assign t[78] = t[99] ^ x[8];
  assign t[79] = t[100] ^ x[9];
  assign t[7] = t[35] ^ t[36];
  assign t[80] = t[101] ^ x[6];
  assign t[81] = t[102] ^ x[10];
  assign t[82] = t[103] ^ x[11];
  assign t[83] = t[104] ^ x[12];
  assign t[84] = t[105] ^ x[7];
  assign t[85] = t[106] ^ x[18];
  assign t[86] = t[107] ^ x[19];
  assign t[87] = t[108] ^ x[23];
  assign t[88] = t[109] ^ x[20];
  assign t[89] = t[110] ^ x[21];
  assign t[8] = t[10] & t[11];
  assign t[90] = t[111] ^ x[22];
  assign t[91] = t[112] ^ x[17];
  assign t[92] = t[113] ^ x[29];
  assign t[93] = t[114] ^ x[30];
  assign t[94] = t[115] ^ x[34];
  assign t[95] = t[116] ^ x[31];
  assign t[96] = t[117] ^ x[32];
  assign t[97] = t[118] ^ x[33];
  assign t[98] = t[119] ^ x[28];
  assign t[99] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[9] = ~(t[12]);
  assign y = (t[0] & ~t[17]) | (~t[0] & t[17]);
endmodule

module R2ind112(x, y);
 input [25:0] x;
 output y;

 wire [90:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[34]);
  assign t[12] = ~(t[33] ^ t[11]);
  assign t[13] = t[35] ^ t[34];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[33] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[33] ^ t[18];
  assign t[18] = t[34] ^ t[36];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[32]);
  assign t[20] = ~(t[21] ^ t[37]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[33] ^ t[11];
  assign t[27] = x[0] ? x[22] : t[28];
  assign t[28] = ~(t[29] ^ t[38]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[31]);
  assign t[31] = t[18] ^ t[7];
  assign t[32] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[33] = (t[41] & ~t[42]) | (~t[41] & t[42]);
  assign t[34] = (t[41] & ~t[44] & ~t[46]) | (~t[43] & t[44] & ~t[45]) | (~t[41] & ~t[44] & t[46]) | (t[43] & t[44] & t[45]);
  assign t[35] = (t[41] & ~t[45]) | (~t[41] & t[45]);
  assign t[36] = (t[41] & ~t[44] & ~t[45]) | (~t[43] & t[44] & ~t[46]) | (~t[41] & ~t[44] & t[45]) | (t[43] & t[44] & t[46]);
  assign t[37] = (t[39] & ~t[47]) | (~t[39] & t[47]);
  assign t[38] = (t[39] & ~t[49] & ~t[50]) | (~t[48] & t[49] & ~t[40]) | (~t[39] & ~t[49] & t[50]) | (t[48] & t[49] & t[40]);
  assign t[39] = t[51] ^ x[7];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[52] ^ x[8];
  assign t[41] = t[53] ^ x[14];
  assign t[42] = t[54] ^ x[15];
  assign t[43] = t[55] ^ x[16];
  assign t[44] = t[56] ^ x[17];
  assign t[45] = t[57] ^ x[18];
  assign t[46] = t[58] ^ x[19];
  assign t[47] = t[59] ^ x[21];
  assign t[48] = t[60] ^ x[23];
  assign t[49] = t[61] ^ x[24];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[62] ^ x[25];
  assign t[51] = (t[63] & ~t[65] & ~t[66] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & ~t[66] & ~t[67] & ~t[69]) | (t[63] & ~t[64] & ~t[65] & ~t[68] & ~t[69]) | (~t[63] & t[64] & t[65] & t[66] & ~t[69]) | (~t[63] & t[64] & t[67] & t[68] & ~t[69]) | (t[63] & ~t[65] & ~t[67] & t[69]) | (~t[63] & t[65] & t[67] & t[69]);
  assign t[52] = (t[63] & t[64] & ~t[65] & ~t[67] & t[68] & ~t[69]) | (t[63] & t[65] & ~t[66] & ~t[67] & ~t[68] & t[69]) | (~t[64] & ~t[65] & t[67] & ~t[68] & ~t[69]) | (~t[63] & ~t[65] & ~t[66] & t[67] & ~t[68]) | (~t[63] & ~t[64] & ~t[66] & t[67] & ~t[69]) | (~t[63] & ~t[65] & t[66] & t[67] & t[68]) | (t[66] & t[67] & ~t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[72] & ~t[73] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & ~t[73] & ~t[74] & ~t[76]) | (t[70] & ~t[71] & ~t[72] & ~t[75] & ~t[76]) | (~t[70] & t[71] & t[72] & t[73] & ~t[76]) | (~t[70] & t[71] & t[74] & t[75] & ~t[76]) | (t[70] & ~t[72] & ~t[74] & t[76]) | (~t[70] & t[72] & t[74] & t[76]);
  assign t[54] = (t[70] & t[71] & ~t[72] & t[73] & ~t[74] & ~t[76]) | (t[70] & ~t[72] & ~t[73] & t[74] & ~t[75] & t[76]) | (~t[71] & t[72] & ~t[73] & ~t[74] & ~t[76]) | (~t[70] & t[72] & ~t[73] & ~t[74] & ~t[75]) | (~t[70] & ~t[71] & t[72] & ~t[75] & ~t[76]) | (~t[70] & t[72] & t[73] & ~t[74] & t[75]) | (t[72] & ~t[73] & t[75] & ~t[76]);
  assign t[55] = (t[71] & ~t[72] & ~t[73] & ~t[74] & ~t[75]) | (~t[70] & t[71] & ~t[73] & ~t[74] & ~t[76]) | (~t[70] & t[71] & ~t[72] & ~t[75] & ~t[76]) | (t[70] & ~t[71] & t[72] & t[73] & ~t[76]) | (t[70] & ~t[71] & t[74] & t[75] & ~t[76]) | (t[71] & ~t[73] & ~t[75] & t[76]) | (~t[71] & t[73] & t[75] & t[76]);
  assign t[56] = (t[70] & t[71] & t[72] & ~t[73] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[73] & ~t[74] & t[75] & t[76]) | (~t[71] & ~t[72] & t[73] & ~t[74] & ~t[75]) | (~t[70] & ~t[72] & t[73] & ~t[75] & ~t[76]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[76]) | (~t[71] & t[72] & t[73] & t[74] & ~t[75]) | (~t[72] & t[73] & t[74] & ~t[76]);
  assign t[57] = (t[70] & t[71] & ~t[72] & ~t[74] & t[75] & ~t[76]) | (t[70] & t[72] & ~t[73] & ~t[74] & ~t[75] & t[76]) | (~t[71] & ~t[72] & t[74] & ~t[75] & ~t[76]) | (~t[70] & ~t[72] & ~t[73] & t[74] & ~t[75]) | (~t[70] & ~t[71] & ~t[73] & t[74] & ~t[76]) | (~t[70] & ~t[72] & t[73] & t[74] & t[75]) | (t[73] & t[74] & ~t[75] & ~t[76]);
  assign t[58] = (t[70] & t[71] & ~t[73] & t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & t[73] & ~t[74] & ~t[75] & t[76]) | (~t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[70] & ~t[71] & ~t[72] & t[75] & ~t[76]) | (~t[71] & t[72] & ~t[73] & t[74] & t[75]) | (t[72] & ~t[74] & t[75] & ~t[76]);
  assign t[59] = (t[63] & t[64] & ~t[65] & t[66] & ~t[67] & ~t[69]) | (t[63] & ~t[65] & ~t[66] & t[67] & ~t[68] & t[69]) | (~t[64] & t[65] & ~t[66] & ~t[67] & ~t[69]) | (~t[63] & t[65] & ~t[66] & ~t[67] & ~t[68]) | (~t[63] & ~t[64] & t[65] & ~t[68] & ~t[69]) | (~t[63] & t[65] & t[66] & ~t[67] & t[68]) | (t[65] & ~t[66] & t[68] & ~t[69]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[64] & ~t[65] & ~t[66] & ~t[67] & ~t[68]) | (~t[63] & t[64] & ~t[66] & ~t[67] & ~t[69]) | (~t[63] & t[64] & ~t[65] & ~t[68] & ~t[69]) | (t[63] & ~t[64] & t[65] & t[66] & ~t[69]) | (t[63] & ~t[64] & t[67] & t[68] & ~t[69]) | (t[64] & ~t[66] & ~t[68] & t[69]) | (~t[64] & t[66] & t[68] & t[69]);
  assign t[61] = (t[63] & t[64] & t[65] & ~t[66] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[66] & ~t[67] & t[68] & t[69]) | (~t[64] & ~t[65] & t[66] & ~t[67] & ~t[68]) | (~t[63] & ~t[65] & t[66] & ~t[68] & ~t[69]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[69]) | (~t[64] & t[65] & t[66] & t[67] & ~t[68]) | (~t[65] & t[66] & t[67] & ~t[69]);
  assign t[62] = (t[63] & t[64] & ~t[66] & t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & t[66] & ~t[67] & ~t[68] & t[69]) | (~t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[63] & ~t[64] & ~t[65] & t[68] & ~t[69]) | (~t[64] & t[65] & ~t[66] & t[67] & t[68]) | (t[65] & ~t[67] & t[68] & ~t[69]);
  assign t[63] = t[77] ^ x[7];
  assign t[64] = t[78] ^ x[23];
  assign t[65] = t[79] ^ x[21];
  assign t[66] = t[80] ^ x[24];
  assign t[67] = t[81] ^ x[8];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[33] & t[10];
  assign t[70] = t[84] ^ x[14];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[15];
  assign t[73] = t[87] ^ x[17];
  assign t[74] = t[88] ^ x[18];
  assign t[75] = t[89] ^ x[19];
  assign t[76] = t[90] ^ x[13];
  assign t[77] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[78] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[79] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[81] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[82] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[83] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[84] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[85] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[86] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[87] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[88] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[89] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[8] = t[13] ^ t[11];
  assign t[90] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27]) | (~t[0] & t[19] & ~t[27]) | (~t[0] & ~t[19] & t[27]) | (t[0] & t[19] & t[27]);
endmodule

module R2ind113(x, y);
 input [25:0] x;
 output y;

 wire [89:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[32] ^ t[11]);
  assign t[13] = t[34] ^ t[33];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[32] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[32] ^ t[18];
  assign t[18] = t[33] ^ t[35];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[31]);
  assign t[20] = ~(t[21] ^ t[36]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[32] ^ t[11];
  assign t[27] = x[0] ? x[22] : t[28];
  assign t[28] = ~(t[29] ^ t[37]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[23]);
  assign t[31] = (t[38] & ~t[39]) | (~t[38] & t[39]);
  assign t[32] = (t[40] & ~t[41]) | (~t[40] & t[41]);
  assign t[33] = (t[40] & ~t[43] & ~t[45]) | (~t[42] & t[43] & ~t[44]) | (~t[40] & ~t[43] & t[45]) | (t[42] & t[43] & t[44]);
  assign t[34] = (t[40] & ~t[44]) | (~t[40] & t[44]);
  assign t[35] = (t[40] & ~t[43] & ~t[44]) | (~t[42] & t[43] & ~t[45]) | (~t[40] & ~t[43] & t[44]) | (t[42] & t[43] & t[45]);
  assign t[36] = (t[38] & ~t[46]) | (~t[38] & t[46]);
  assign t[37] = (t[38] & ~t[48] & ~t[39]) | (~t[47] & t[48] & ~t[49]) | (~t[38] & ~t[48] & t[39]) | (t[47] & t[48] & t[49]);
  assign t[38] = t[50] ^ x[7];
  assign t[39] = t[51] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[52] ^ x[14];
  assign t[41] = t[53] ^ x[15];
  assign t[42] = t[54] ^ x[16];
  assign t[43] = t[55] ^ x[17];
  assign t[44] = t[56] ^ x[18];
  assign t[45] = t[57] ^ x[19];
  assign t[46] = t[58] ^ x[21];
  assign t[47] = t[59] ^ x[23];
  assign t[48] = t[60] ^ x[24];
  assign t[49] = t[61] ^ x[25];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[51] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[53] = (t[69] & t[70] & ~t[71] & t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[71] & ~t[72] & t[73] & ~t[74] & t[75]) | (~t[70] & t[71] & ~t[72] & ~t[73] & ~t[75]) | (~t[69] & t[71] & ~t[72] & ~t[73] & ~t[74]) | (~t[69] & ~t[70] & t[71] & ~t[74] & ~t[75]) | (~t[69] & t[71] & t[72] & ~t[73] & t[74]) | (t[71] & ~t[72] & t[74] & ~t[75]);
  assign t[54] = (t[70] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (~t[69] & t[70] & ~t[72] & ~t[73] & ~t[75]) | (~t[69] & t[70] & ~t[71] & ~t[74] & ~t[75]) | (t[69] & ~t[70] & t[71] & t[72] & ~t[75]) | (t[69] & ~t[70] & t[73] & t[74] & ~t[75]) | (t[70] & ~t[72] & ~t[74] & t[75]) | (~t[70] & t[72] & t[74] & t[75]);
  assign t[55] = (t[69] & t[70] & t[71] & ~t[72] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & ~t[72] & ~t[73] & t[74] & t[75]) | (~t[70] & ~t[71] & t[72] & ~t[73] & ~t[74]) | (~t[69] & ~t[71] & t[72] & ~t[74] & ~t[75]) | (~t[69] & ~t[70] & t[72] & ~t[73] & ~t[75]) | (~t[70] & t[71] & t[72] & t[73] & ~t[74]) | (~t[71] & t[72] & t[73] & ~t[75]);
  assign t[56] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[57] = (t[69] & t[70] & ~t[72] & t[73] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & ~t[72] & ~t[73] & t[74]) | (~t[69] & ~t[72] & ~t[73] & t[74] & ~t[75]) | (~t[69] & ~t[70] & ~t[71] & t[74] & ~t[75]) | (~t[70] & t[71] & ~t[72] & t[73] & t[74]) | (t[71] & ~t[73] & t[74] & ~t[75]);
  assign t[58] = (t[62] & t[63] & ~t[64] & t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[64] & ~t[65] & t[66] & ~t[67] & t[68]) | (~t[63] & t[64] & ~t[65] & ~t[66] & ~t[68]) | (~t[62] & t[64] & ~t[65] & ~t[66] & ~t[67]) | (~t[62] & ~t[63] & t[64] & ~t[67] & ~t[68]) | (~t[62] & t[64] & t[65] & ~t[66] & t[67]) | (t[64] & ~t[65] & t[67] & ~t[68]);
  assign t[59] = (t[63] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (~t[62] & t[63] & ~t[65] & ~t[66] & ~t[68]) | (~t[62] & t[63] & ~t[64] & ~t[67] & ~t[68]) | (t[62] & ~t[63] & t[64] & t[65] & ~t[68]) | (t[62] & ~t[63] & t[66] & t[67] & ~t[68]) | (t[63] & ~t[65] & ~t[67] & t[68]) | (~t[63] & t[65] & t[67] & t[68]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[62] & t[63] & t[64] & ~t[65] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & ~t[65] & ~t[66] & t[67] & t[68]) | (~t[63] & ~t[64] & t[65] & ~t[66] & ~t[67]) | (~t[62] & ~t[64] & t[65] & ~t[67] & ~t[68]) | (~t[62] & ~t[63] & t[65] & ~t[66] & ~t[68]) | (~t[63] & t[64] & t[65] & t[66] & ~t[67]) | (~t[64] & t[65] & t[66] & ~t[68]);
  assign t[61] = (t[62] & t[63] & ~t[65] & t[66] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[65] & ~t[66] & t[67] & ~t[68]) | (~t[62] & ~t[63] & ~t[64] & t[67] & ~t[68]) | (~t[63] & t[64] & ~t[65] & t[66] & t[67]) | (t[64] & ~t[66] & t[67] & ~t[68]);
  assign t[62] = t[76] ^ x[7];
  assign t[63] = t[77] ^ x[23];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[24];
  assign t[66] = t[80] ^ x[8];
  assign t[67] = t[81] ^ x[25];
  assign t[68] = t[82] ^ x[6];
  assign t[69] = t[83] ^ x[14];
  assign t[6] = t[32] & t[10];
  assign t[70] = t[84] ^ x[16];
  assign t[71] = t[85] ^ x[15];
  assign t[72] = t[86] ^ x[17];
  assign t[73] = t[87] ^ x[18];
  assign t[74] = t[88] ^ x[19];
  assign t[75] = t[89] ^ x[13];
  assign t[76] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[77] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[78] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[79] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[81] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[82] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[83] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[84] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[85] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[86] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[87] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[88] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[89] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27]) | (~t[0] & t[19] & ~t[27]) | (~t[0] & ~t[19] & t[27]) | (t[0] & t[19] & t[27]);
endmodule

module R2ind114(x, y);
 input [24:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[25] ^ t[11]);
  assign t[13] = t[27] ^ t[26];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[25] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[25] ^ t[18];
  assign t[18] = t[26] ^ t[28];
  assign t[19] = x[0] ? x[21] : t[20];
  assign t[1] = ~(t[2] ^ t[24]);
  assign t[20] = ~(t[21] ^ t[29]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[18] ^ t[7];
  assign t[24] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[25] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[26] = (t[32] & ~t[35] & ~t[37]) | (~t[34] & t[35] & ~t[36]) | (~t[32] & ~t[35] & t[37]) | (t[34] & t[35] & t[36]);
  assign t[27] = (t[32] & ~t[36]) | (~t[32] & t[36]);
  assign t[28] = (t[32] & ~t[35] & ~t[36]) | (~t[34] & t[35] & ~t[37]) | (~t[32] & ~t[35] & t[36]) | (t[34] & t[35] & t[37]);
  assign t[29] = (t[30] & ~t[39] & ~t[40]) | (~t[38] & t[39] & ~t[31]) | (~t[30] & ~t[39] & t[40]) | (t[38] & t[39] & t[31]);
  assign t[2] = ~t[3];
  assign t[30] = t[41] ^ x[8];
  assign t[31] = t[42] ^ x[9];
  assign t[32] = t[43] ^ x[15];
  assign t[33] = t[44] ^ x[16];
  assign t[34] = t[45] ^ x[17];
  assign t[35] = t[46] ^ x[18];
  assign t[36] = t[47] ^ x[19];
  assign t[37] = t[48] ^ x[20];
  assign t[38] = t[49] ^ x[22];
  assign t[39] = t[50] ^ x[23];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[51] ^ x[24];
  assign t[41] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[42] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[43] = (t[59] & ~t[61] & ~t[62] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & ~t[62] & ~t[63] & ~t[65]) | (t[59] & ~t[60] & ~t[61] & ~t[64] & ~t[65]) | (~t[59] & t[60] & t[61] & t[62] & ~t[65]) | (~t[59] & t[60] & t[63] & t[64] & ~t[65]) | (t[59] & ~t[61] & ~t[63] & t[65]) | (~t[59] & t[61] & t[63] & t[65]);
  assign t[44] = (t[59] & t[60] & ~t[61] & t[62] & ~t[63] & ~t[65]) | (t[59] & ~t[61] & ~t[62] & t[63] & ~t[64] & t[65]) | (~t[60] & t[61] & ~t[62] & ~t[63] & ~t[65]) | (~t[59] & t[61] & ~t[62] & ~t[63] & ~t[64]) | (~t[59] & ~t[60] & t[61] & ~t[64] & ~t[65]) | (~t[59] & t[61] & t[62] & ~t[63] & t[64]) | (t[61] & ~t[62] & t[64] & ~t[65]);
  assign t[45] = (t[60] & ~t[61] & ~t[62] & ~t[63] & ~t[64]) | (~t[59] & t[60] & ~t[62] & ~t[63] & ~t[65]) | (~t[59] & t[60] & ~t[61] & ~t[64] & ~t[65]) | (t[59] & ~t[60] & t[61] & t[62] & ~t[65]) | (t[59] & ~t[60] & t[63] & t[64] & ~t[65]) | (t[60] & ~t[62] & ~t[64] & t[65]) | (~t[60] & t[62] & t[64] & t[65]);
  assign t[46] = (t[59] & t[60] & t[61] & ~t[62] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[62] & ~t[63] & t[64] & t[65]) | (~t[60] & ~t[61] & t[62] & ~t[63] & ~t[64]) | (~t[59] & ~t[61] & t[62] & ~t[64] & ~t[65]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[65]) | (~t[60] & t[61] & t[62] & t[63] & ~t[64]) | (~t[61] & t[62] & t[63] & ~t[65]);
  assign t[47] = (t[59] & t[60] & ~t[61] & ~t[63] & t[64] & ~t[65]) | (t[59] & t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[65]) | (~t[59] & ~t[61] & ~t[62] & t[63] & ~t[64]) | (~t[59] & ~t[60] & ~t[62] & t[63] & ~t[65]) | (~t[59] & ~t[61] & t[62] & t[63] & t[64]) | (t[62] & t[63] & ~t[64] & ~t[65]);
  assign t[48] = (t[59] & t[60] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[59] & ~t[60] & ~t[61] & t[64] & ~t[65]) | (~t[60] & t[61] & ~t[62] & t[63] & t[64]) | (t[61] & ~t[63] & t[64] & ~t[65]);
  assign t[49] = (t[53] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (~t[52] & t[53] & ~t[55] & ~t[56] & ~t[58]) | (~t[52] & t[53] & ~t[54] & ~t[57] & ~t[58]) | (t[52] & ~t[53] & t[54] & t[55] & ~t[58]) | (t[52] & ~t[53] & t[56] & t[57] & ~t[58]) | (t[53] & ~t[55] & ~t[57] & t[58]) | (~t[53] & t[55] & t[57] & t[58]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[52] & t[53] & t[54] & ~t[55] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[55] & ~t[56] & t[57] & t[58]) | (~t[53] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (~t[52] & ~t[54] & t[55] & ~t[57] & ~t[58]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[58]) | (~t[53] & t[54] & t[55] & t[56] & ~t[57]) | (~t[54] & t[55] & t[56] & ~t[58]);
  assign t[51] = (t[52] & t[53] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[52] & ~t[53] & ~t[54] & t[57] & ~t[58]) | (~t[53] & t[54] & ~t[55] & t[56] & t[57]) | (t[54] & ~t[56] & t[57] & ~t[58]);
  assign t[52] = t[66] ^ x[8];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[6];
  assign t[55] = t[69] ^ x[23];
  assign t[56] = t[70] ^ x[9];
  assign t[57] = t[71] ^ x[24];
  assign t[58] = t[72] ^ x[7];
  assign t[59] = t[73] ^ x[15];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[16];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[19];
  assign t[64] = t[78] ^ x[20];
  assign t[65] = t[79] ^ x[14];
  assign t[66] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[67] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[68] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[69] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[6] = t[25] & t[10];
  assign t[70] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[71] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[72] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[73] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[74] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[75] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[76] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[77] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[78] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[79] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind115(x, y);
 input [24:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[26] ^ t[11]);
  assign t[13] = t[28] ^ t[27];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[26] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[26] ^ t[18];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = x[0] ? x[21] : t[20];
  assign t[1] = ~(t[2] ^ t[25]);
  assign t[20] = ~(t[21] ^ t[30]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[24] ^ t[7];
  assign t[24] = t[13] ^ t[16];
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[27] = (t[33] & ~t[36] & ~t[38]) | (~t[35] & t[36] & ~t[37]) | (~t[33] & ~t[36] & t[38]) | (t[35] & t[36] & t[37]);
  assign t[28] = (t[33] & ~t[37]) | (~t[33] & t[37]);
  assign t[29] = (t[33] & ~t[36] & ~t[37]) | (~t[35] & t[36] & ~t[38]) | (~t[33] & ~t[36] & t[37]) | (t[35] & t[36] & t[38]);
  assign t[2] = ~t[3];
  assign t[30] = (t[31] & ~t[40] & ~t[32]) | (~t[39] & t[40] & ~t[41]) | (~t[31] & ~t[40] & t[32]) | (t[39] & t[40] & t[41]);
  assign t[31] = t[42] ^ x[8];
  assign t[32] = t[43] ^ x[9];
  assign t[33] = t[44] ^ x[15];
  assign t[34] = t[45] ^ x[16];
  assign t[35] = t[46] ^ x[17];
  assign t[36] = t[47] ^ x[18];
  assign t[37] = t[48] ^ x[19];
  assign t[38] = t[49] ^ x[20];
  assign t[39] = t[50] ^ x[22];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[51] ^ x[23];
  assign t[41] = t[52] ^ x[24];
  assign t[42] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[43] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[45] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[51] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[8];
  assign t[54] = t[68] ^ x[22];
  assign t[55] = t[69] ^ x[6];
  assign t[56] = t[70] ^ x[23];
  assign t[57] = t[71] ^ x[9];
  assign t[58] = t[72] ^ x[24];
  assign t[59] = t[73] ^ x[7];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[74] ^ x[15];
  assign t[61] = t[75] ^ x[17];
  assign t[62] = t[76] ^ x[16];
  assign t[63] = t[77] ^ x[18];
  assign t[64] = t[78] ^ x[19];
  assign t[65] = t[79] ^ x[20];
  assign t[66] = t[80] ^ x[14];
  assign t[67] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[68] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[69] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[6] = t[26] & t[10];
  assign t[70] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[71] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[72] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[73] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[74] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[75] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[76] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[77] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[78] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[79] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind116(x, y);
 input [24:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[25] ^ t[12]);
  assign t[14] = t[25] & t[16];
  assign t[15] = t[25] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[27] ^ t[28];
  assign t[18] = t[25] ^ t[10];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[24]);
  assign t[20] = ~(t[21] ^ t[29]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[17] ^ t[7];
  assign t[24] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[25] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[26] = (t[32] & ~t[34]) | (~t[32] & t[34]);
  assign t[27] = (t[32] & ~t[36] & ~t[37]) | (~t[35] & t[36] & ~t[34]) | (~t[32] & ~t[36] & t[37]) | (t[35] & t[36] & t[34]);
  assign t[28] = (t[32] & ~t[36] & ~t[34]) | (~t[35] & t[36] & ~t[37]) | (~t[32] & ~t[36] & t[34]) | (t[35] & t[36] & t[37]);
  assign t[29] = (t[30] & ~t[39] & ~t[41]) | (~t[38] & t[39] & ~t[40]) | (~t[30] & ~t[39] & t[41]) | (t[38] & t[39] & t[40]);
  assign t[2] = ~t[3];
  assign t[30] = t[42] ^ x[7];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[18];
  assign t[37] = t[49] ^ x[19];
  assign t[38] = t[50] ^ x[21];
  assign t[39] = t[51] ^ x[22];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[52] ^ x[23];
  assign t[41] = t[53] ^ x[24];
  assign t[42] = (t[54] & ~t[56] & ~t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[57] & ~t[58] & ~t[60]) | (t[54] & ~t[55] & ~t[56] & ~t[59] & ~t[60]) | (~t[54] & t[55] & t[56] & t[57] & ~t[60]) | (~t[54] & t[55] & t[58] & t[59] & ~t[60]) | (t[54] & ~t[56] & ~t[58] & t[60]) | (~t[54] & t[56] & t[58] & t[60]);
  assign t[43] = (t[54] & t[55] & ~t[56] & t[57] & ~t[58] & ~t[60]) | (t[54] & ~t[56] & ~t[57] & t[58] & ~t[59] & t[60]) | (~t[55] & t[56] & ~t[57] & ~t[58] & ~t[60]) | (~t[54] & t[56] & ~t[57] & ~t[58] & ~t[59]) | (~t[54] & ~t[55] & t[56] & ~t[59] & ~t[60]) | (~t[54] & t[56] & t[57] & ~t[58] & t[59]) | (t[56] & ~t[57] & t[59] & ~t[60]);
  assign t[44] = (t[61] & ~t[63] & ~t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[64] & ~t[65] & ~t[67]) | (t[61] & ~t[62] & ~t[63] & ~t[66] & ~t[67]) | (~t[61] & t[62] & t[63] & t[64] & ~t[67]) | (~t[61] & t[62] & t[65] & t[66] & ~t[67]) | (t[61] & ~t[63] & ~t[65] & t[67]) | (~t[61] & t[63] & t[65] & t[67]);
  assign t[45] = (t[61] & t[62] & ~t[63] & t[64] & ~t[65] & ~t[67]) | (t[61] & ~t[63] & ~t[64] & t[65] & ~t[66] & t[67]) | (~t[62] & t[63] & ~t[64] & ~t[65] & ~t[67]) | (~t[61] & t[63] & ~t[64] & ~t[65] & ~t[66]) | (~t[61] & ~t[62] & t[63] & ~t[66] & ~t[67]) | (~t[61] & t[63] & t[64] & ~t[65] & t[66]) | (t[63] & ~t[64] & t[66] & ~t[67]);
  assign t[46] = (t[61] & t[62] & ~t[63] & ~t[65] & t[66] & ~t[67]) | (t[61] & t[63] & ~t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[63] & t[65] & ~t[66] & ~t[67]) | (~t[61] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[61] & ~t[62] & ~t[64] & t[65] & ~t[67]) | (~t[61] & ~t[63] & t[64] & t[65] & t[66]) | (t[64] & t[65] & ~t[66] & ~t[67]);
  assign t[47] = (t[62] & ~t[63] & ~t[64] & ~t[65] & ~t[66]) | (~t[61] & t[62] & ~t[64] & ~t[65] & ~t[67]) | (~t[61] & t[62] & ~t[63] & ~t[66] & ~t[67]) | (t[61] & ~t[62] & t[63] & t[64] & ~t[67]) | (t[61] & ~t[62] & t[65] & t[66] & ~t[67]) | (t[62] & ~t[64] & ~t[66] & t[67]) | (~t[62] & t[64] & t[66] & t[67]);
  assign t[48] = (t[61] & t[62] & t[63] & ~t[64] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[64] & ~t[65] & t[66] & t[67]) | (~t[62] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (~t[61] & ~t[63] & t[64] & ~t[66] & ~t[67]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[67]) | (~t[62] & t[63] & t[64] & t[65] & ~t[66]) | (~t[63] & t[64] & t[65] & ~t[67]);
  assign t[49] = (t[61] & t[62] & ~t[64] & t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[61] & ~t[62] & ~t[63] & t[66] & ~t[67]) | (~t[62] & t[63] & ~t[64] & t[65] & t[66]) | (t[63] & ~t[65] & t[66] & ~t[67]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[55] & ~t[56] & ~t[57] & ~t[58] & ~t[59]) | (~t[54] & t[55] & ~t[57] & ~t[58] & ~t[60]) | (~t[54] & t[55] & ~t[56] & ~t[59] & ~t[60]) | (t[54] & ~t[55] & t[56] & t[57] & ~t[60]) | (t[54] & ~t[55] & t[58] & t[59] & ~t[60]) | (t[55] & ~t[57] & ~t[59] & t[60]) | (~t[55] & t[57] & t[59] & t[60]);
  assign t[51] = (t[54] & t[55] & t[56] & ~t[57] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[57] & ~t[58] & t[59] & t[60]) | (~t[55] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (~t[54] & ~t[56] & t[57] & ~t[59] & ~t[60]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[60]) | (~t[55] & t[56] & t[57] & t[58] & ~t[59]) | (~t[56] & t[57] & t[58] & ~t[60]);
  assign t[52] = (t[54] & t[55] & ~t[56] & ~t[58] & t[59] & ~t[60]) | (t[54] & t[56] & ~t[57] & ~t[58] & ~t[59] & t[60]) | (~t[55] & ~t[56] & t[58] & ~t[59] & ~t[60]) | (~t[54] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[54] & ~t[55] & ~t[57] & t[58] & ~t[60]) | (~t[54] & ~t[56] & t[57] & t[58] & t[59]) | (t[57] & t[58] & ~t[59] & ~t[60]);
  assign t[53] = (t[54] & t[55] & ~t[57] & t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & t[57] & ~t[58] & ~t[59] & t[60]) | (~t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[54] & ~t[55] & ~t[56] & t[59] & ~t[60]) | (~t[55] & t[56] & ~t[57] & t[58] & t[59]) | (t[56] & ~t[58] & t[59] & ~t[60]);
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[8];
  assign t[57] = t[71] ^ x[22];
  assign t[58] = t[72] ^ x[23];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[74] ^ x[6];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[17];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[16];
  assign t[66] = t[80] ^ x[19];
  assign t[67] = t[81] ^ x[13];
  assign t[68] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[69] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[71] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[72] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[73] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[74] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[75] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[76] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[77] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[78] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[79] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[7] = t[12] & t[13];
  assign t[80] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[81] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[25] ^ t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind117(x, y);
 input [24:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[25] ^ t[26];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[26]);
  assign t[13] = ~(t[24] ^ t[12]);
  assign t[14] = t[24] & t[16];
  assign t[15] = t[24] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[26] ^ t[27];
  assign t[18] = t[24] ^ t[10];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[23]);
  assign t[20] = ~(t[21] ^ t[28]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[4]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[25] = (t[31] & ~t[33]) | (~t[31] & t[33]);
  assign t[26] = (t[31] & ~t[35] & ~t[36]) | (~t[34] & t[35] & ~t[33]) | (~t[31] & ~t[35] & t[36]) | (t[34] & t[35] & t[33]);
  assign t[27] = (t[31] & ~t[35] & ~t[33]) | (~t[34] & t[35] & ~t[36]) | (~t[31] & ~t[35] & t[33]) | (t[34] & t[35] & t[36]);
  assign t[28] = (t[29] & ~t[38] & ~t[39]) | (~t[37] & t[38] & ~t[40]) | (~t[29] & ~t[38] & t[39]) | (t[37] & t[38] & t[40]);
  assign t[29] = t[41] ^ x[7];
  assign t[2] = ~t[3];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[14];
  assign t[32] = t[44] ^ x[15];
  assign t[33] = t[45] ^ x[16];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = t[48] ^ x[19];
  assign t[37] = t[49] ^ x[21];
  assign t[38] = t[50] ^ x[22];
  assign t[39] = t[51] ^ x[23];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[52] ^ x[24];
  assign t[41] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[42] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[44] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[45] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[7];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[8];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[23];
  assign t[58] = t[72] ^ x[24];
  assign t[59] = t[73] ^ x[6];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[74] ^ x[14];
  assign t[61] = t[75] ^ x[17];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[18];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = t[79] ^ x[19];
  assign t[66] = t[80] ^ x[13];
  assign t[67] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[68] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[69] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[71] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[72] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[73] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[74] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[75] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[76] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[77] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[78] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[79] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[7] = t[12] & t[13];
  assign t[80] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[24] ^ t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind118(x, y);
 input [24:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[11] ^ t[22]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[6];
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[19];
  assign t[16] = t[7] & t[17];
  assign t[17] = t[21] ^ t[5];
  assign t[18] = (t[24] & ~t[26] & ~t[28]) | (~t[25] & t[26] & ~t[27]) | (~t[24] & ~t[26] & t[28]) | (t[25] & t[26] & t[27]);
  assign t[19] = (t[29] & ~t[31] & ~t[33]) | (~t[30] & t[31] & ~t[32]) | (~t[29] & ~t[31] & t[33]) | (t[30] & t[31] & t[32]);
  assign t[1] = ~(t[2] ^ t[18]);
  assign t[20] = (t[29] & ~t[31] & ~t[32]) | (~t[30] & t[31] & ~t[33]) | (~t[29] & ~t[31] & t[32]) | (t[30] & t[31] & t[33]);
  assign t[21] = (t[29] & ~t[34]) | (~t[29] & t[34]);
  assign t[22] = (t[24] & ~t[26] & ~t[27]) | (~t[25] & t[26] & ~t[28]) | (~t[24] & ~t[26] & t[27]) | (t[25] & t[26] & t[28]);
  assign t[23] = (t[29] & ~t[32]) | (~t[29] & t[32]);
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[9];
  assign t[26] = t[37] ^ x[10];
  assign t[27] = t[38] ^ x[11];
  assign t[28] = t[39] ^ x[12];
  assign t[29] = t[40] ^ x[18];
  assign t[2] = ~t[3];
  assign t[30] = t[41] ^ x[19];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[23];
  assign t[35] = (t[46] & ~t[48] & ~t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[49] & ~t[50] & ~t[52]) | (t[46] & ~t[47] & ~t[48] & ~t[51] & ~t[52]) | (~t[46] & t[47] & t[48] & t[49] & ~t[52]) | (~t[46] & t[47] & t[50] & t[51] & ~t[52]) | (t[46] & ~t[48] & ~t[50] & t[52]) | (~t[46] & t[48] & t[50] & t[52]);
  assign t[36] = (t[47] & ~t[48] & ~t[49] & ~t[50] & ~t[51]) | (~t[46] & t[47] & ~t[49] & ~t[50] & ~t[52]) | (~t[46] & t[47] & ~t[48] & ~t[51] & ~t[52]) | (t[46] & ~t[47] & t[48] & t[49] & ~t[52]) | (t[46] & ~t[47] & t[50] & t[51] & ~t[52]) | (t[47] & ~t[49] & ~t[51] & t[52]) | (~t[47] & t[49] & t[51] & t[52]);
  assign t[37] = (t[46] & t[47] & t[48] & ~t[49] & ~t[51] & ~t[52]) | (t[47] & ~t[48] & ~t[49] & ~t[50] & t[51] & t[52]) | (~t[47] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (~t[46] & ~t[48] & t[49] & ~t[51] & ~t[52]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[52]) | (~t[47] & t[48] & t[49] & t[50] & ~t[51]) | (~t[48] & t[49] & t[50] & ~t[52]);
  assign t[38] = (t[46] & t[47] & ~t[48] & ~t[50] & t[51] & ~t[52]) | (t[46] & t[48] & ~t[49] & ~t[50] & ~t[51] & t[52]) | (~t[47] & ~t[48] & t[50] & ~t[51] & ~t[52]) | (~t[46] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[46] & ~t[47] & ~t[49] & t[50] & ~t[52]) | (~t[46] & ~t[48] & t[49] & t[50] & t[51]) | (t[49] & t[50] & ~t[51] & ~t[52]);
  assign t[39] = (t[46] & t[47] & ~t[49] & t[50] & ~t[51] & ~t[52]) | (t[47] & ~t[48] & t[49] & ~t[50] & ~t[51] & t[52]) | (~t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[49] & ~t[50] & t[51] & ~t[52]) | (~t[46] & ~t[47] & ~t[48] & t[51] & ~t[52]) | (~t[47] & t[48] & ~t[49] & t[50] & t[51]) | (t[48] & ~t[50] & t[51] & ~t[52]);
  assign t[3] = ~(t[4]);
  assign t[40] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[41] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[42] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[43] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[44] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[45] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[6];
  assign t[49] = t[63] ^ x[10];
  assign t[4] = t[5] ^ t[6];
  assign t[50] = t[64] ^ x[11];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[7];
  assign t[53] = t[67] ^ x[18];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[23];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = t[19] ^ t[20];
  assign t[60] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[61] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[62] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[63] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[64] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[65] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[66] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[67] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = t[7] & t[8];
  assign t[70] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[71] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[72] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[73] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[7] = ~(t[19]);
  assign t[8] = ~(t[21] ^ t[7]);
  assign t[9] = x[0] ? x[24] : t[10];
  assign y = (t[0] & ~t[9]) | (~t[0] & t[9]);
endmodule

module R2ind119(x, y);
 input [25:0] x;
 output y;

 wire [90:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[34]);
  assign t[12] = ~(t[33] ^ t[11]);
  assign t[13] = t[35] ^ t[34];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[33] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[33] ^ t[18];
  assign t[18] = t[34] ^ t[36];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[32]);
  assign t[20] = ~(t[21] ^ t[37]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[33] ^ t[11];
  assign t[27] = x[0] ? x[22] : t[28];
  assign t[28] = ~(t[29] ^ t[38]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[31]);
  assign t[31] = t[18] ^ t[7];
  assign t[32] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[33] = (t[41] & ~t[42]) | (~t[41] & t[42]);
  assign t[34] = (t[41] & ~t[44] & ~t[46]) | (~t[43] & t[44] & ~t[45]) | (~t[41] & ~t[44] & t[46]) | (t[43] & t[44] & t[45]);
  assign t[35] = (t[41] & ~t[45]) | (~t[41] & t[45]);
  assign t[36] = (t[41] & ~t[44] & ~t[45]) | (~t[43] & t[44] & ~t[46]) | (~t[41] & ~t[44] & t[45]) | (t[43] & t[44] & t[46]);
  assign t[37] = (t[39] & ~t[47]) | (~t[39] & t[47]);
  assign t[38] = (t[39] & ~t[49] & ~t[50]) | (~t[48] & t[49] & ~t[40]) | (~t[39] & ~t[49] & t[50]) | (t[48] & t[49] & t[40]);
  assign t[39] = t[51] ^ x[7];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[52] ^ x[8];
  assign t[41] = t[53] ^ x[14];
  assign t[42] = t[54] ^ x[15];
  assign t[43] = t[55] ^ x[16];
  assign t[44] = t[56] ^ x[17];
  assign t[45] = t[57] ^ x[18];
  assign t[46] = t[58] ^ x[19];
  assign t[47] = t[59] ^ x[21];
  assign t[48] = t[60] ^ x[23];
  assign t[49] = t[61] ^ x[24];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[62] ^ x[25];
  assign t[51] = (t[63] & ~t[65] & ~t[66] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & ~t[66] & ~t[67] & ~t[69]) | (t[63] & ~t[64] & ~t[65] & ~t[68] & ~t[69]) | (~t[63] & t[64] & t[65] & t[66] & ~t[69]) | (~t[63] & t[64] & t[67] & t[68] & ~t[69]) | (t[63] & ~t[65] & ~t[67] & t[69]) | (~t[63] & t[65] & t[67] & t[69]);
  assign t[52] = (t[63] & t[64] & ~t[65] & ~t[67] & t[68] & ~t[69]) | (t[63] & t[65] & ~t[66] & ~t[67] & ~t[68] & t[69]) | (~t[64] & ~t[65] & t[67] & ~t[68] & ~t[69]) | (~t[63] & ~t[65] & ~t[66] & t[67] & ~t[68]) | (~t[63] & ~t[64] & ~t[66] & t[67] & ~t[69]) | (~t[63] & ~t[65] & t[66] & t[67] & t[68]) | (t[66] & t[67] & ~t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[72] & ~t[73] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & ~t[73] & ~t[74] & ~t[76]) | (t[70] & ~t[71] & ~t[72] & ~t[75] & ~t[76]) | (~t[70] & t[71] & t[72] & t[73] & ~t[76]) | (~t[70] & t[71] & t[74] & t[75] & ~t[76]) | (t[70] & ~t[72] & ~t[74] & t[76]) | (~t[70] & t[72] & t[74] & t[76]);
  assign t[54] = (t[70] & t[71] & ~t[72] & t[73] & ~t[74] & ~t[76]) | (t[70] & ~t[72] & ~t[73] & t[74] & ~t[75] & t[76]) | (~t[71] & t[72] & ~t[73] & ~t[74] & ~t[76]) | (~t[70] & t[72] & ~t[73] & ~t[74] & ~t[75]) | (~t[70] & ~t[71] & t[72] & ~t[75] & ~t[76]) | (~t[70] & t[72] & t[73] & ~t[74] & t[75]) | (t[72] & ~t[73] & t[75] & ~t[76]);
  assign t[55] = (t[71] & ~t[72] & ~t[73] & ~t[74] & ~t[75]) | (~t[70] & t[71] & ~t[73] & ~t[74] & ~t[76]) | (~t[70] & t[71] & ~t[72] & ~t[75] & ~t[76]) | (t[70] & ~t[71] & t[72] & t[73] & ~t[76]) | (t[70] & ~t[71] & t[74] & t[75] & ~t[76]) | (t[71] & ~t[73] & ~t[75] & t[76]) | (~t[71] & t[73] & t[75] & t[76]);
  assign t[56] = (t[70] & t[71] & t[72] & ~t[73] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[73] & ~t[74] & t[75] & t[76]) | (~t[71] & ~t[72] & t[73] & ~t[74] & ~t[75]) | (~t[70] & ~t[72] & t[73] & ~t[75] & ~t[76]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[76]) | (~t[71] & t[72] & t[73] & t[74] & ~t[75]) | (~t[72] & t[73] & t[74] & ~t[76]);
  assign t[57] = (t[70] & t[71] & ~t[72] & ~t[74] & t[75] & ~t[76]) | (t[70] & t[72] & ~t[73] & ~t[74] & ~t[75] & t[76]) | (~t[71] & ~t[72] & t[74] & ~t[75] & ~t[76]) | (~t[70] & ~t[72] & ~t[73] & t[74] & ~t[75]) | (~t[70] & ~t[71] & ~t[73] & t[74] & ~t[76]) | (~t[70] & ~t[72] & t[73] & t[74] & t[75]) | (t[73] & t[74] & ~t[75] & ~t[76]);
  assign t[58] = (t[70] & t[71] & ~t[73] & t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & t[73] & ~t[74] & ~t[75] & t[76]) | (~t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[70] & ~t[71] & ~t[72] & t[75] & ~t[76]) | (~t[71] & t[72] & ~t[73] & t[74] & t[75]) | (t[72] & ~t[74] & t[75] & ~t[76]);
  assign t[59] = (t[63] & t[64] & ~t[65] & t[66] & ~t[67] & ~t[69]) | (t[63] & ~t[65] & ~t[66] & t[67] & ~t[68] & t[69]) | (~t[64] & t[65] & ~t[66] & ~t[67] & ~t[69]) | (~t[63] & t[65] & ~t[66] & ~t[67] & ~t[68]) | (~t[63] & ~t[64] & t[65] & ~t[68] & ~t[69]) | (~t[63] & t[65] & t[66] & ~t[67] & t[68]) | (t[65] & ~t[66] & t[68] & ~t[69]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[64] & ~t[65] & ~t[66] & ~t[67] & ~t[68]) | (~t[63] & t[64] & ~t[66] & ~t[67] & ~t[69]) | (~t[63] & t[64] & ~t[65] & ~t[68] & ~t[69]) | (t[63] & ~t[64] & t[65] & t[66] & ~t[69]) | (t[63] & ~t[64] & t[67] & t[68] & ~t[69]) | (t[64] & ~t[66] & ~t[68] & t[69]) | (~t[64] & t[66] & t[68] & t[69]);
  assign t[61] = (t[63] & t[64] & t[65] & ~t[66] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[66] & ~t[67] & t[68] & t[69]) | (~t[64] & ~t[65] & t[66] & ~t[67] & ~t[68]) | (~t[63] & ~t[65] & t[66] & ~t[68] & ~t[69]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[69]) | (~t[64] & t[65] & t[66] & t[67] & ~t[68]) | (~t[65] & t[66] & t[67] & ~t[69]);
  assign t[62] = (t[63] & t[64] & ~t[66] & t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & t[66] & ~t[67] & ~t[68] & t[69]) | (~t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[63] & ~t[64] & ~t[65] & t[68] & ~t[69]) | (~t[64] & t[65] & ~t[66] & t[67] & t[68]) | (t[65] & ~t[67] & t[68] & ~t[69]);
  assign t[63] = t[77] ^ x[7];
  assign t[64] = t[78] ^ x[23];
  assign t[65] = t[79] ^ x[21];
  assign t[66] = t[80] ^ x[24];
  assign t[67] = t[81] ^ x[8];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[33] & t[10];
  assign t[70] = t[84] ^ x[14];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[15];
  assign t[73] = t[87] ^ x[17];
  assign t[74] = t[88] ^ x[18];
  assign t[75] = t[89] ^ x[19];
  assign t[76] = t[90] ^ x[13];
  assign t[77] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[78] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[79] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[81] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[82] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[83] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[84] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[85] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[86] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[87] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[88] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[89] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[8] = t[13] ^ t[11];
  assign t[90] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27]) | (~t[0] & t[19] & ~t[27]) | (~t[0] & ~t[19] & t[27]) | (t[0] & t[19] & t[27]);
endmodule

module R2ind120(x, y);
 input [25:0] x;
 output y;

 wire [89:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[32] ^ t[11]);
  assign t[13] = t[34] ^ t[33];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[32] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[32] ^ t[18];
  assign t[18] = t[33] ^ t[35];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[31]);
  assign t[20] = ~(t[21] ^ t[36]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[32] ^ t[11];
  assign t[27] = x[0] ? x[22] : t[28];
  assign t[28] = ~(t[29] ^ t[37]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[23]);
  assign t[31] = (t[38] & ~t[39]) | (~t[38] & t[39]);
  assign t[32] = (t[40] & ~t[41]) | (~t[40] & t[41]);
  assign t[33] = (t[40] & ~t[43] & ~t[45]) | (~t[42] & t[43] & ~t[44]) | (~t[40] & ~t[43] & t[45]) | (t[42] & t[43] & t[44]);
  assign t[34] = (t[40] & ~t[44]) | (~t[40] & t[44]);
  assign t[35] = (t[40] & ~t[43] & ~t[44]) | (~t[42] & t[43] & ~t[45]) | (~t[40] & ~t[43] & t[44]) | (t[42] & t[43] & t[45]);
  assign t[36] = (t[38] & ~t[46]) | (~t[38] & t[46]);
  assign t[37] = (t[38] & ~t[48] & ~t[39]) | (~t[47] & t[48] & ~t[49]) | (~t[38] & ~t[48] & t[39]) | (t[47] & t[48] & t[49]);
  assign t[38] = t[50] ^ x[7];
  assign t[39] = t[51] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[52] ^ x[14];
  assign t[41] = t[53] ^ x[15];
  assign t[42] = t[54] ^ x[16];
  assign t[43] = t[55] ^ x[17];
  assign t[44] = t[56] ^ x[18];
  assign t[45] = t[57] ^ x[19];
  assign t[46] = t[58] ^ x[21];
  assign t[47] = t[59] ^ x[23];
  assign t[48] = t[60] ^ x[24];
  assign t[49] = t[61] ^ x[25];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[51] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[53] = (t[69] & t[70] & ~t[71] & t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[71] & ~t[72] & t[73] & ~t[74] & t[75]) | (~t[70] & t[71] & ~t[72] & ~t[73] & ~t[75]) | (~t[69] & t[71] & ~t[72] & ~t[73] & ~t[74]) | (~t[69] & ~t[70] & t[71] & ~t[74] & ~t[75]) | (~t[69] & t[71] & t[72] & ~t[73] & t[74]) | (t[71] & ~t[72] & t[74] & ~t[75]);
  assign t[54] = (t[70] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (~t[69] & t[70] & ~t[72] & ~t[73] & ~t[75]) | (~t[69] & t[70] & ~t[71] & ~t[74] & ~t[75]) | (t[69] & ~t[70] & t[71] & t[72] & ~t[75]) | (t[69] & ~t[70] & t[73] & t[74] & ~t[75]) | (t[70] & ~t[72] & ~t[74] & t[75]) | (~t[70] & t[72] & t[74] & t[75]);
  assign t[55] = (t[69] & t[70] & t[71] & ~t[72] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & ~t[72] & ~t[73] & t[74] & t[75]) | (~t[70] & ~t[71] & t[72] & ~t[73] & ~t[74]) | (~t[69] & ~t[71] & t[72] & ~t[74] & ~t[75]) | (~t[69] & ~t[70] & t[72] & ~t[73] & ~t[75]) | (~t[70] & t[71] & t[72] & t[73] & ~t[74]) | (~t[71] & t[72] & t[73] & ~t[75]);
  assign t[56] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[57] = (t[69] & t[70] & ~t[72] & t[73] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & ~t[72] & ~t[73] & t[74]) | (~t[69] & ~t[72] & ~t[73] & t[74] & ~t[75]) | (~t[69] & ~t[70] & ~t[71] & t[74] & ~t[75]) | (~t[70] & t[71] & ~t[72] & t[73] & t[74]) | (t[71] & ~t[73] & t[74] & ~t[75]);
  assign t[58] = (t[62] & t[63] & ~t[64] & t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[64] & ~t[65] & t[66] & ~t[67] & t[68]) | (~t[63] & t[64] & ~t[65] & ~t[66] & ~t[68]) | (~t[62] & t[64] & ~t[65] & ~t[66] & ~t[67]) | (~t[62] & ~t[63] & t[64] & ~t[67] & ~t[68]) | (~t[62] & t[64] & t[65] & ~t[66] & t[67]) | (t[64] & ~t[65] & t[67] & ~t[68]);
  assign t[59] = (t[63] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (~t[62] & t[63] & ~t[65] & ~t[66] & ~t[68]) | (~t[62] & t[63] & ~t[64] & ~t[67] & ~t[68]) | (t[62] & ~t[63] & t[64] & t[65] & ~t[68]) | (t[62] & ~t[63] & t[66] & t[67] & ~t[68]) | (t[63] & ~t[65] & ~t[67] & t[68]) | (~t[63] & t[65] & t[67] & t[68]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[62] & t[63] & t[64] & ~t[65] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & ~t[65] & ~t[66] & t[67] & t[68]) | (~t[63] & ~t[64] & t[65] & ~t[66] & ~t[67]) | (~t[62] & ~t[64] & t[65] & ~t[67] & ~t[68]) | (~t[62] & ~t[63] & t[65] & ~t[66] & ~t[68]) | (~t[63] & t[64] & t[65] & t[66] & ~t[67]) | (~t[64] & t[65] & t[66] & ~t[68]);
  assign t[61] = (t[62] & t[63] & ~t[65] & t[66] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[65] & ~t[66] & t[67] & ~t[68]) | (~t[62] & ~t[63] & ~t[64] & t[67] & ~t[68]) | (~t[63] & t[64] & ~t[65] & t[66] & t[67]) | (t[64] & ~t[66] & t[67] & ~t[68]);
  assign t[62] = t[76] ^ x[7];
  assign t[63] = t[77] ^ x[23];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[24];
  assign t[66] = t[80] ^ x[8];
  assign t[67] = t[81] ^ x[25];
  assign t[68] = t[82] ^ x[6];
  assign t[69] = t[83] ^ x[14];
  assign t[6] = t[32] & t[10];
  assign t[70] = t[84] ^ x[16];
  assign t[71] = t[85] ^ x[15];
  assign t[72] = t[86] ^ x[17];
  assign t[73] = t[87] ^ x[18];
  assign t[74] = t[88] ^ x[19];
  assign t[75] = t[89] ^ x[13];
  assign t[76] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[77] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[78] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[79] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[81] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[82] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[83] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[84] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[85] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[86] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[87] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[88] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[89] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27]) | (~t[0] & t[19] & ~t[27]) | (~t[0] & ~t[19] & t[27]) | (t[0] & t[19] & t[27]);
endmodule

module R2ind121(x, y);
 input [24:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[25] ^ t[11]);
  assign t[13] = t[27] ^ t[26];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[25] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[25] ^ t[18];
  assign t[18] = t[26] ^ t[28];
  assign t[19] = x[0] ? x[21] : t[20];
  assign t[1] = ~(t[2] ^ t[24]);
  assign t[20] = ~(t[21] ^ t[29]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[18] ^ t[7];
  assign t[24] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[25] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[26] = (t[32] & ~t[35] & ~t[37]) | (~t[34] & t[35] & ~t[36]) | (~t[32] & ~t[35] & t[37]) | (t[34] & t[35] & t[36]);
  assign t[27] = (t[32] & ~t[36]) | (~t[32] & t[36]);
  assign t[28] = (t[32] & ~t[35] & ~t[36]) | (~t[34] & t[35] & ~t[37]) | (~t[32] & ~t[35] & t[36]) | (t[34] & t[35] & t[37]);
  assign t[29] = (t[30] & ~t[39] & ~t[40]) | (~t[38] & t[39] & ~t[31]) | (~t[30] & ~t[39] & t[40]) | (t[38] & t[39] & t[31]);
  assign t[2] = ~t[3];
  assign t[30] = t[41] ^ x[8];
  assign t[31] = t[42] ^ x[9];
  assign t[32] = t[43] ^ x[15];
  assign t[33] = t[44] ^ x[16];
  assign t[34] = t[45] ^ x[17];
  assign t[35] = t[46] ^ x[18];
  assign t[36] = t[47] ^ x[19];
  assign t[37] = t[48] ^ x[20];
  assign t[38] = t[49] ^ x[22];
  assign t[39] = t[50] ^ x[23];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[51] ^ x[24];
  assign t[41] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[42] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[43] = (t[59] & ~t[61] & ~t[62] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & ~t[62] & ~t[63] & ~t[65]) | (t[59] & ~t[60] & ~t[61] & ~t[64] & ~t[65]) | (~t[59] & t[60] & t[61] & t[62] & ~t[65]) | (~t[59] & t[60] & t[63] & t[64] & ~t[65]) | (t[59] & ~t[61] & ~t[63] & t[65]) | (~t[59] & t[61] & t[63] & t[65]);
  assign t[44] = (t[59] & t[60] & ~t[61] & t[62] & ~t[63] & ~t[65]) | (t[59] & ~t[61] & ~t[62] & t[63] & ~t[64] & t[65]) | (~t[60] & t[61] & ~t[62] & ~t[63] & ~t[65]) | (~t[59] & t[61] & ~t[62] & ~t[63] & ~t[64]) | (~t[59] & ~t[60] & t[61] & ~t[64] & ~t[65]) | (~t[59] & t[61] & t[62] & ~t[63] & t[64]) | (t[61] & ~t[62] & t[64] & ~t[65]);
  assign t[45] = (t[60] & ~t[61] & ~t[62] & ~t[63] & ~t[64]) | (~t[59] & t[60] & ~t[62] & ~t[63] & ~t[65]) | (~t[59] & t[60] & ~t[61] & ~t[64] & ~t[65]) | (t[59] & ~t[60] & t[61] & t[62] & ~t[65]) | (t[59] & ~t[60] & t[63] & t[64] & ~t[65]) | (t[60] & ~t[62] & ~t[64] & t[65]) | (~t[60] & t[62] & t[64] & t[65]);
  assign t[46] = (t[59] & t[60] & t[61] & ~t[62] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[62] & ~t[63] & t[64] & t[65]) | (~t[60] & ~t[61] & t[62] & ~t[63] & ~t[64]) | (~t[59] & ~t[61] & t[62] & ~t[64] & ~t[65]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[65]) | (~t[60] & t[61] & t[62] & t[63] & ~t[64]) | (~t[61] & t[62] & t[63] & ~t[65]);
  assign t[47] = (t[59] & t[60] & ~t[61] & ~t[63] & t[64] & ~t[65]) | (t[59] & t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[65]) | (~t[59] & ~t[61] & ~t[62] & t[63] & ~t[64]) | (~t[59] & ~t[60] & ~t[62] & t[63] & ~t[65]) | (~t[59] & ~t[61] & t[62] & t[63] & t[64]) | (t[62] & t[63] & ~t[64] & ~t[65]);
  assign t[48] = (t[59] & t[60] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[59] & ~t[60] & ~t[61] & t[64] & ~t[65]) | (~t[60] & t[61] & ~t[62] & t[63] & t[64]) | (t[61] & ~t[63] & t[64] & ~t[65]);
  assign t[49] = (t[53] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (~t[52] & t[53] & ~t[55] & ~t[56] & ~t[58]) | (~t[52] & t[53] & ~t[54] & ~t[57] & ~t[58]) | (t[52] & ~t[53] & t[54] & t[55] & ~t[58]) | (t[52] & ~t[53] & t[56] & t[57] & ~t[58]) | (t[53] & ~t[55] & ~t[57] & t[58]) | (~t[53] & t[55] & t[57] & t[58]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[52] & t[53] & t[54] & ~t[55] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[55] & ~t[56] & t[57] & t[58]) | (~t[53] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (~t[52] & ~t[54] & t[55] & ~t[57] & ~t[58]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[58]) | (~t[53] & t[54] & t[55] & t[56] & ~t[57]) | (~t[54] & t[55] & t[56] & ~t[58]);
  assign t[51] = (t[52] & t[53] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[52] & ~t[53] & ~t[54] & t[57] & ~t[58]) | (~t[53] & t[54] & ~t[55] & t[56] & t[57]) | (t[54] & ~t[56] & t[57] & ~t[58]);
  assign t[52] = t[66] ^ x[8];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[6];
  assign t[55] = t[69] ^ x[23];
  assign t[56] = t[70] ^ x[9];
  assign t[57] = t[71] ^ x[24];
  assign t[58] = t[72] ^ x[7];
  assign t[59] = t[73] ^ x[15];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[16];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[19];
  assign t[64] = t[78] ^ x[20];
  assign t[65] = t[79] ^ x[14];
  assign t[66] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[67] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[68] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[69] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[6] = t[25] & t[10];
  assign t[70] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[71] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[72] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[73] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[74] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[75] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[76] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[77] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[78] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[79] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind122(x, y);
 input [24:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[26] ^ t[11]);
  assign t[13] = t[28] ^ t[27];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[26] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[26] ^ t[18];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = x[0] ? x[21] : t[20];
  assign t[1] = ~(t[2] ^ t[25]);
  assign t[20] = ~(t[21] ^ t[30]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[24] ^ t[7];
  assign t[24] = t[13] ^ t[16];
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[27] = (t[33] & ~t[36] & ~t[38]) | (~t[35] & t[36] & ~t[37]) | (~t[33] & ~t[36] & t[38]) | (t[35] & t[36] & t[37]);
  assign t[28] = (t[33] & ~t[37]) | (~t[33] & t[37]);
  assign t[29] = (t[33] & ~t[36] & ~t[37]) | (~t[35] & t[36] & ~t[38]) | (~t[33] & ~t[36] & t[37]) | (t[35] & t[36] & t[38]);
  assign t[2] = ~t[3];
  assign t[30] = (t[31] & ~t[40] & ~t[32]) | (~t[39] & t[40] & ~t[41]) | (~t[31] & ~t[40] & t[32]) | (t[39] & t[40] & t[41]);
  assign t[31] = t[42] ^ x[8];
  assign t[32] = t[43] ^ x[9];
  assign t[33] = t[44] ^ x[15];
  assign t[34] = t[45] ^ x[16];
  assign t[35] = t[46] ^ x[17];
  assign t[36] = t[47] ^ x[18];
  assign t[37] = t[48] ^ x[19];
  assign t[38] = t[49] ^ x[20];
  assign t[39] = t[50] ^ x[22];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[51] ^ x[23];
  assign t[41] = t[52] ^ x[24];
  assign t[42] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[43] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[45] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[51] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[8];
  assign t[54] = t[68] ^ x[22];
  assign t[55] = t[69] ^ x[6];
  assign t[56] = t[70] ^ x[23];
  assign t[57] = t[71] ^ x[9];
  assign t[58] = t[72] ^ x[24];
  assign t[59] = t[73] ^ x[7];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[74] ^ x[15];
  assign t[61] = t[75] ^ x[17];
  assign t[62] = t[76] ^ x[16];
  assign t[63] = t[77] ^ x[18];
  assign t[64] = t[78] ^ x[19];
  assign t[65] = t[79] ^ x[20];
  assign t[66] = t[80] ^ x[14];
  assign t[67] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[68] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[69] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[6] = t[26] & t[10];
  assign t[70] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[71] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[72] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[73] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[74] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[75] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[76] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[77] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[78] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[79] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind123(x, y);
 input [24:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[25] ^ t[12]);
  assign t[14] = t[25] & t[16];
  assign t[15] = t[25] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[27] ^ t[28];
  assign t[18] = t[25] ^ t[10];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[24]);
  assign t[20] = ~(t[21] ^ t[29]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[17] ^ t[7];
  assign t[24] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[25] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[26] = (t[32] & ~t[34]) | (~t[32] & t[34]);
  assign t[27] = (t[32] & ~t[36] & ~t[37]) | (~t[35] & t[36] & ~t[34]) | (~t[32] & ~t[36] & t[37]) | (t[35] & t[36] & t[34]);
  assign t[28] = (t[32] & ~t[36] & ~t[34]) | (~t[35] & t[36] & ~t[37]) | (~t[32] & ~t[36] & t[34]) | (t[35] & t[36] & t[37]);
  assign t[29] = (t[30] & ~t[39] & ~t[41]) | (~t[38] & t[39] & ~t[40]) | (~t[30] & ~t[39] & t[41]) | (t[38] & t[39] & t[40]);
  assign t[2] = ~t[3];
  assign t[30] = t[42] ^ x[7];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[18];
  assign t[37] = t[49] ^ x[19];
  assign t[38] = t[50] ^ x[21];
  assign t[39] = t[51] ^ x[22];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[52] ^ x[23];
  assign t[41] = t[53] ^ x[24];
  assign t[42] = (t[54] & ~t[56] & ~t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[57] & ~t[58] & ~t[60]) | (t[54] & ~t[55] & ~t[56] & ~t[59] & ~t[60]) | (~t[54] & t[55] & t[56] & t[57] & ~t[60]) | (~t[54] & t[55] & t[58] & t[59] & ~t[60]) | (t[54] & ~t[56] & ~t[58] & t[60]) | (~t[54] & t[56] & t[58] & t[60]);
  assign t[43] = (t[54] & t[55] & ~t[56] & t[57] & ~t[58] & ~t[60]) | (t[54] & ~t[56] & ~t[57] & t[58] & ~t[59] & t[60]) | (~t[55] & t[56] & ~t[57] & ~t[58] & ~t[60]) | (~t[54] & t[56] & ~t[57] & ~t[58] & ~t[59]) | (~t[54] & ~t[55] & t[56] & ~t[59] & ~t[60]) | (~t[54] & t[56] & t[57] & ~t[58] & t[59]) | (t[56] & ~t[57] & t[59] & ~t[60]);
  assign t[44] = (t[61] & ~t[63] & ~t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[64] & ~t[65] & ~t[67]) | (t[61] & ~t[62] & ~t[63] & ~t[66] & ~t[67]) | (~t[61] & t[62] & t[63] & t[64] & ~t[67]) | (~t[61] & t[62] & t[65] & t[66] & ~t[67]) | (t[61] & ~t[63] & ~t[65] & t[67]) | (~t[61] & t[63] & t[65] & t[67]);
  assign t[45] = (t[61] & t[62] & ~t[63] & t[64] & ~t[65] & ~t[67]) | (t[61] & ~t[63] & ~t[64] & t[65] & ~t[66] & t[67]) | (~t[62] & t[63] & ~t[64] & ~t[65] & ~t[67]) | (~t[61] & t[63] & ~t[64] & ~t[65] & ~t[66]) | (~t[61] & ~t[62] & t[63] & ~t[66] & ~t[67]) | (~t[61] & t[63] & t[64] & ~t[65] & t[66]) | (t[63] & ~t[64] & t[66] & ~t[67]);
  assign t[46] = (t[61] & t[62] & ~t[63] & ~t[65] & t[66] & ~t[67]) | (t[61] & t[63] & ~t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[63] & t[65] & ~t[66] & ~t[67]) | (~t[61] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[61] & ~t[62] & ~t[64] & t[65] & ~t[67]) | (~t[61] & ~t[63] & t[64] & t[65] & t[66]) | (t[64] & t[65] & ~t[66] & ~t[67]);
  assign t[47] = (t[62] & ~t[63] & ~t[64] & ~t[65] & ~t[66]) | (~t[61] & t[62] & ~t[64] & ~t[65] & ~t[67]) | (~t[61] & t[62] & ~t[63] & ~t[66] & ~t[67]) | (t[61] & ~t[62] & t[63] & t[64] & ~t[67]) | (t[61] & ~t[62] & t[65] & t[66] & ~t[67]) | (t[62] & ~t[64] & ~t[66] & t[67]) | (~t[62] & t[64] & t[66] & t[67]);
  assign t[48] = (t[61] & t[62] & t[63] & ~t[64] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[64] & ~t[65] & t[66] & t[67]) | (~t[62] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (~t[61] & ~t[63] & t[64] & ~t[66] & ~t[67]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[67]) | (~t[62] & t[63] & t[64] & t[65] & ~t[66]) | (~t[63] & t[64] & t[65] & ~t[67]);
  assign t[49] = (t[61] & t[62] & ~t[64] & t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[61] & ~t[62] & ~t[63] & t[66] & ~t[67]) | (~t[62] & t[63] & ~t[64] & t[65] & t[66]) | (t[63] & ~t[65] & t[66] & ~t[67]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[55] & ~t[56] & ~t[57] & ~t[58] & ~t[59]) | (~t[54] & t[55] & ~t[57] & ~t[58] & ~t[60]) | (~t[54] & t[55] & ~t[56] & ~t[59] & ~t[60]) | (t[54] & ~t[55] & t[56] & t[57] & ~t[60]) | (t[54] & ~t[55] & t[58] & t[59] & ~t[60]) | (t[55] & ~t[57] & ~t[59] & t[60]) | (~t[55] & t[57] & t[59] & t[60]);
  assign t[51] = (t[54] & t[55] & t[56] & ~t[57] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[57] & ~t[58] & t[59] & t[60]) | (~t[55] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (~t[54] & ~t[56] & t[57] & ~t[59] & ~t[60]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[60]) | (~t[55] & t[56] & t[57] & t[58] & ~t[59]) | (~t[56] & t[57] & t[58] & ~t[60]);
  assign t[52] = (t[54] & t[55] & ~t[56] & ~t[58] & t[59] & ~t[60]) | (t[54] & t[56] & ~t[57] & ~t[58] & ~t[59] & t[60]) | (~t[55] & ~t[56] & t[58] & ~t[59] & ~t[60]) | (~t[54] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[54] & ~t[55] & ~t[57] & t[58] & ~t[60]) | (~t[54] & ~t[56] & t[57] & t[58] & t[59]) | (t[57] & t[58] & ~t[59] & ~t[60]);
  assign t[53] = (t[54] & t[55] & ~t[57] & t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & t[57] & ~t[58] & ~t[59] & t[60]) | (~t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[54] & ~t[55] & ~t[56] & t[59] & ~t[60]) | (~t[55] & t[56] & ~t[57] & t[58] & t[59]) | (t[56] & ~t[58] & t[59] & ~t[60]);
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[8];
  assign t[57] = t[71] ^ x[22];
  assign t[58] = t[72] ^ x[23];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[74] ^ x[6];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[17];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[16];
  assign t[66] = t[80] ^ x[19];
  assign t[67] = t[81] ^ x[13];
  assign t[68] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[69] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[71] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[72] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[73] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[74] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[75] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[76] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[77] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[78] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[79] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[7] = t[12] & t[13];
  assign t[80] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[81] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[25] ^ t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind124(x, y);
 input [24:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[25] ^ t[26];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[26]);
  assign t[13] = ~(t[24] ^ t[12]);
  assign t[14] = t[24] & t[16];
  assign t[15] = t[24] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[26] ^ t[27];
  assign t[18] = t[24] ^ t[10];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[23]);
  assign t[20] = ~(t[21] ^ t[28]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[4]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[25] = (t[31] & ~t[33]) | (~t[31] & t[33]);
  assign t[26] = (t[31] & ~t[35] & ~t[36]) | (~t[34] & t[35] & ~t[33]) | (~t[31] & ~t[35] & t[36]) | (t[34] & t[35] & t[33]);
  assign t[27] = (t[31] & ~t[35] & ~t[33]) | (~t[34] & t[35] & ~t[36]) | (~t[31] & ~t[35] & t[33]) | (t[34] & t[35] & t[36]);
  assign t[28] = (t[29] & ~t[38] & ~t[39]) | (~t[37] & t[38] & ~t[40]) | (~t[29] & ~t[38] & t[39]) | (t[37] & t[38] & t[40]);
  assign t[29] = t[41] ^ x[7];
  assign t[2] = ~t[3];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[14];
  assign t[32] = t[44] ^ x[15];
  assign t[33] = t[45] ^ x[16];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = t[48] ^ x[19];
  assign t[37] = t[49] ^ x[21];
  assign t[38] = t[50] ^ x[22];
  assign t[39] = t[51] ^ x[23];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[52] ^ x[24];
  assign t[41] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[42] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[44] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[45] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[7];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[8];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[23];
  assign t[58] = t[72] ^ x[24];
  assign t[59] = t[73] ^ x[6];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[74] ^ x[14];
  assign t[61] = t[75] ^ x[17];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[18];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = t[79] ^ x[19];
  assign t[66] = t[80] ^ x[13];
  assign t[67] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[68] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[69] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[71] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[72] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[73] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[74] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[75] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[76] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[77] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[78] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[79] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[7] = t[12] & t[13];
  assign t[80] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[24] ^ t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind125(x, y);
 input [24:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[11] ^ t[22]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[6];
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[19];
  assign t[16] = t[7] & t[17];
  assign t[17] = t[21] ^ t[5];
  assign t[18] = (t[24] & ~t[26] & ~t[28]) | (~t[25] & t[26] & ~t[27]) | (~t[24] & ~t[26] & t[28]) | (t[25] & t[26] & t[27]);
  assign t[19] = (t[29] & ~t[31] & ~t[33]) | (~t[30] & t[31] & ~t[32]) | (~t[29] & ~t[31] & t[33]) | (t[30] & t[31] & t[32]);
  assign t[1] = ~(t[2] ^ t[18]);
  assign t[20] = (t[29] & ~t[31] & ~t[32]) | (~t[30] & t[31] & ~t[33]) | (~t[29] & ~t[31] & t[32]) | (t[30] & t[31] & t[33]);
  assign t[21] = (t[29] & ~t[34]) | (~t[29] & t[34]);
  assign t[22] = (t[24] & ~t[26] & ~t[27]) | (~t[25] & t[26] & ~t[28]) | (~t[24] & ~t[26] & t[27]) | (t[25] & t[26] & t[28]);
  assign t[23] = (t[29] & ~t[32]) | (~t[29] & t[32]);
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[9];
  assign t[26] = t[37] ^ x[10];
  assign t[27] = t[38] ^ x[11];
  assign t[28] = t[39] ^ x[12];
  assign t[29] = t[40] ^ x[18];
  assign t[2] = ~t[3];
  assign t[30] = t[41] ^ x[19];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[23];
  assign t[35] = (t[46] & ~t[48] & ~t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[49] & ~t[50] & ~t[52]) | (t[46] & ~t[47] & ~t[48] & ~t[51] & ~t[52]) | (~t[46] & t[47] & t[48] & t[49] & ~t[52]) | (~t[46] & t[47] & t[50] & t[51] & ~t[52]) | (t[46] & ~t[48] & ~t[50] & t[52]) | (~t[46] & t[48] & t[50] & t[52]);
  assign t[36] = (t[47] & ~t[48] & ~t[49] & ~t[50] & ~t[51]) | (~t[46] & t[47] & ~t[49] & ~t[50] & ~t[52]) | (~t[46] & t[47] & ~t[48] & ~t[51] & ~t[52]) | (t[46] & ~t[47] & t[48] & t[49] & ~t[52]) | (t[46] & ~t[47] & t[50] & t[51] & ~t[52]) | (t[47] & ~t[49] & ~t[51] & t[52]) | (~t[47] & t[49] & t[51] & t[52]);
  assign t[37] = (t[46] & t[47] & t[48] & ~t[49] & ~t[51] & ~t[52]) | (t[47] & ~t[48] & ~t[49] & ~t[50] & t[51] & t[52]) | (~t[47] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (~t[46] & ~t[48] & t[49] & ~t[51] & ~t[52]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[52]) | (~t[47] & t[48] & t[49] & t[50] & ~t[51]) | (~t[48] & t[49] & t[50] & ~t[52]);
  assign t[38] = (t[46] & t[47] & ~t[48] & ~t[50] & t[51] & ~t[52]) | (t[46] & t[48] & ~t[49] & ~t[50] & ~t[51] & t[52]) | (~t[47] & ~t[48] & t[50] & ~t[51] & ~t[52]) | (~t[46] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[46] & ~t[47] & ~t[49] & t[50] & ~t[52]) | (~t[46] & ~t[48] & t[49] & t[50] & t[51]) | (t[49] & t[50] & ~t[51] & ~t[52]);
  assign t[39] = (t[46] & t[47] & ~t[49] & t[50] & ~t[51] & ~t[52]) | (t[47] & ~t[48] & t[49] & ~t[50] & ~t[51] & t[52]) | (~t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[49] & ~t[50] & t[51] & ~t[52]) | (~t[46] & ~t[47] & ~t[48] & t[51] & ~t[52]) | (~t[47] & t[48] & ~t[49] & t[50] & t[51]) | (t[48] & ~t[50] & t[51] & ~t[52]);
  assign t[3] = ~(t[4]);
  assign t[40] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[41] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[42] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[43] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[44] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[45] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[6];
  assign t[49] = t[63] ^ x[10];
  assign t[4] = t[5] ^ t[6];
  assign t[50] = t[64] ^ x[11];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[7];
  assign t[53] = t[67] ^ x[18];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[23];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = t[19] ^ t[20];
  assign t[60] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[61] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[62] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[63] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[64] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[65] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[66] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[67] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = t[7] & t[8];
  assign t[70] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[71] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[72] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[73] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[7] = ~(t[19]);
  assign t[8] = ~(t[21] ^ t[7]);
  assign t[9] = x[0] ? x[24] : t[10];
  assign y = (t[0] & ~t[9]) | (~t[0] & t[9]);
endmodule

module R2ind126(x, y);
 input [25:0] x;
 output y;

 wire [90:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[34]);
  assign t[12] = ~(t[33] ^ t[11]);
  assign t[13] = t[35] ^ t[34];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[33] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[33] ^ t[18];
  assign t[18] = t[34] ^ t[36];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[32]);
  assign t[20] = ~(t[21] ^ t[37]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[33] ^ t[11];
  assign t[27] = x[0] ? x[22] : t[28];
  assign t[28] = ~(t[29] ^ t[38]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[31]);
  assign t[31] = t[18] ^ t[7];
  assign t[32] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[33] = (t[41] & ~t[42]) | (~t[41] & t[42]);
  assign t[34] = (t[41] & ~t[44] & ~t[46]) | (~t[43] & t[44] & ~t[45]) | (~t[41] & ~t[44] & t[46]) | (t[43] & t[44] & t[45]);
  assign t[35] = (t[41] & ~t[45]) | (~t[41] & t[45]);
  assign t[36] = (t[41] & ~t[44] & ~t[45]) | (~t[43] & t[44] & ~t[46]) | (~t[41] & ~t[44] & t[45]) | (t[43] & t[44] & t[46]);
  assign t[37] = (t[39] & ~t[47]) | (~t[39] & t[47]);
  assign t[38] = (t[39] & ~t[49] & ~t[50]) | (~t[48] & t[49] & ~t[40]) | (~t[39] & ~t[49] & t[50]) | (t[48] & t[49] & t[40]);
  assign t[39] = t[51] ^ x[7];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[52] ^ x[8];
  assign t[41] = t[53] ^ x[14];
  assign t[42] = t[54] ^ x[15];
  assign t[43] = t[55] ^ x[16];
  assign t[44] = t[56] ^ x[17];
  assign t[45] = t[57] ^ x[18];
  assign t[46] = t[58] ^ x[19];
  assign t[47] = t[59] ^ x[21];
  assign t[48] = t[60] ^ x[23];
  assign t[49] = t[61] ^ x[24];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = t[62] ^ x[25];
  assign t[51] = (t[63] & ~t[65] & ~t[66] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & ~t[66] & ~t[67] & ~t[69]) | (t[63] & ~t[64] & ~t[65] & ~t[68] & ~t[69]) | (~t[63] & t[64] & t[65] & t[66] & ~t[69]) | (~t[63] & t[64] & t[67] & t[68] & ~t[69]) | (t[63] & ~t[65] & ~t[67] & t[69]) | (~t[63] & t[65] & t[67] & t[69]);
  assign t[52] = (t[63] & t[64] & ~t[65] & ~t[67] & t[68] & ~t[69]) | (t[63] & t[65] & ~t[66] & ~t[67] & ~t[68] & t[69]) | (~t[64] & ~t[65] & t[67] & ~t[68] & ~t[69]) | (~t[63] & ~t[65] & ~t[66] & t[67] & ~t[68]) | (~t[63] & ~t[64] & ~t[66] & t[67] & ~t[69]) | (~t[63] & ~t[65] & t[66] & t[67] & t[68]) | (t[66] & t[67] & ~t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[72] & ~t[73] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & ~t[73] & ~t[74] & ~t[76]) | (t[70] & ~t[71] & ~t[72] & ~t[75] & ~t[76]) | (~t[70] & t[71] & t[72] & t[73] & ~t[76]) | (~t[70] & t[71] & t[74] & t[75] & ~t[76]) | (t[70] & ~t[72] & ~t[74] & t[76]) | (~t[70] & t[72] & t[74] & t[76]);
  assign t[54] = (t[70] & t[71] & ~t[72] & t[73] & ~t[74] & ~t[76]) | (t[70] & ~t[72] & ~t[73] & t[74] & ~t[75] & t[76]) | (~t[71] & t[72] & ~t[73] & ~t[74] & ~t[76]) | (~t[70] & t[72] & ~t[73] & ~t[74] & ~t[75]) | (~t[70] & ~t[71] & t[72] & ~t[75] & ~t[76]) | (~t[70] & t[72] & t[73] & ~t[74] & t[75]) | (t[72] & ~t[73] & t[75] & ~t[76]);
  assign t[55] = (t[71] & ~t[72] & ~t[73] & ~t[74] & ~t[75]) | (~t[70] & t[71] & ~t[73] & ~t[74] & ~t[76]) | (~t[70] & t[71] & ~t[72] & ~t[75] & ~t[76]) | (t[70] & ~t[71] & t[72] & t[73] & ~t[76]) | (t[70] & ~t[71] & t[74] & t[75] & ~t[76]) | (t[71] & ~t[73] & ~t[75] & t[76]) | (~t[71] & t[73] & t[75] & t[76]);
  assign t[56] = (t[70] & t[71] & t[72] & ~t[73] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & ~t[73] & ~t[74] & t[75] & t[76]) | (~t[71] & ~t[72] & t[73] & ~t[74] & ~t[75]) | (~t[70] & ~t[72] & t[73] & ~t[75] & ~t[76]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[76]) | (~t[71] & t[72] & t[73] & t[74] & ~t[75]) | (~t[72] & t[73] & t[74] & ~t[76]);
  assign t[57] = (t[70] & t[71] & ~t[72] & ~t[74] & t[75] & ~t[76]) | (t[70] & t[72] & ~t[73] & ~t[74] & ~t[75] & t[76]) | (~t[71] & ~t[72] & t[74] & ~t[75] & ~t[76]) | (~t[70] & ~t[72] & ~t[73] & t[74] & ~t[75]) | (~t[70] & ~t[71] & ~t[73] & t[74] & ~t[76]) | (~t[70] & ~t[72] & t[73] & t[74] & t[75]) | (t[73] & t[74] & ~t[75] & ~t[76]);
  assign t[58] = (t[70] & t[71] & ~t[73] & t[74] & ~t[75] & ~t[76]) | (t[71] & ~t[72] & t[73] & ~t[74] & ~t[75] & t[76]) | (~t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[73] & ~t[74] & t[75] & ~t[76]) | (~t[70] & ~t[71] & ~t[72] & t[75] & ~t[76]) | (~t[71] & t[72] & ~t[73] & t[74] & t[75]) | (t[72] & ~t[74] & t[75] & ~t[76]);
  assign t[59] = (t[63] & t[64] & ~t[65] & t[66] & ~t[67] & ~t[69]) | (t[63] & ~t[65] & ~t[66] & t[67] & ~t[68] & t[69]) | (~t[64] & t[65] & ~t[66] & ~t[67] & ~t[69]) | (~t[63] & t[65] & ~t[66] & ~t[67] & ~t[68]) | (~t[63] & ~t[64] & t[65] & ~t[68] & ~t[69]) | (~t[63] & t[65] & t[66] & ~t[67] & t[68]) | (t[65] & ~t[66] & t[68] & ~t[69]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[64] & ~t[65] & ~t[66] & ~t[67] & ~t[68]) | (~t[63] & t[64] & ~t[66] & ~t[67] & ~t[69]) | (~t[63] & t[64] & ~t[65] & ~t[68] & ~t[69]) | (t[63] & ~t[64] & t[65] & t[66] & ~t[69]) | (t[63] & ~t[64] & t[67] & t[68] & ~t[69]) | (t[64] & ~t[66] & ~t[68] & t[69]) | (~t[64] & t[66] & t[68] & t[69]);
  assign t[61] = (t[63] & t[64] & t[65] & ~t[66] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & ~t[66] & ~t[67] & t[68] & t[69]) | (~t[64] & ~t[65] & t[66] & ~t[67] & ~t[68]) | (~t[63] & ~t[65] & t[66] & ~t[68] & ~t[69]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[69]) | (~t[64] & t[65] & t[66] & t[67] & ~t[68]) | (~t[65] & t[66] & t[67] & ~t[69]);
  assign t[62] = (t[63] & t[64] & ~t[66] & t[67] & ~t[68] & ~t[69]) | (t[64] & ~t[65] & t[66] & ~t[67] & ~t[68] & t[69]) | (~t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[66] & ~t[67] & t[68] & ~t[69]) | (~t[63] & ~t[64] & ~t[65] & t[68] & ~t[69]) | (~t[64] & t[65] & ~t[66] & t[67] & t[68]) | (t[65] & ~t[67] & t[68] & ~t[69]);
  assign t[63] = t[77] ^ x[7];
  assign t[64] = t[78] ^ x[23];
  assign t[65] = t[79] ^ x[21];
  assign t[66] = t[80] ^ x[24];
  assign t[67] = t[81] ^ x[8];
  assign t[68] = t[82] ^ x[25];
  assign t[69] = t[83] ^ x[6];
  assign t[6] = t[33] & t[10];
  assign t[70] = t[84] ^ x[14];
  assign t[71] = t[85] ^ x[16];
  assign t[72] = t[86] ^ x[15];
  assign t[73] = t[87] ^ x[17];
  assign t[74] = t[88] ^ x[18];
  assign t[75] = t[89] ^ x[19];
  assign t[76] = t[90] ^ x[13];
  assign t[77] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[78] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[79] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[81] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[82] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[83] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[84] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[85] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[86] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[87] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[88] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[89] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[8] = t[13] ^ t[11];
  assign t[90] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27]) | (~t[0] & t[19] & ~t[27]) | (~t[0] & ~t[19] & t[27]) | (t[0] & t[19] & t[27]);
endmodule

module R2ind127(x, y);
 input [25:0] x;
 output y;

 wire [89:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[33]);
  assign t[12] = ~(t[32] ^ t[11]);
  assign t[13] = t[34] ^ t[33];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[32] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[32] ^ t[18];
  assign t[18] = t[33] ^ t[35];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[31]);
  assign t[20] = ~(t[21] ^ t[36]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23] ^ t[24]);
  assign t[23] = t[25] ^ t[7];
  assign t[24] = t[4] ^ t[26];
  assign t[25] = t[13] ^ t[16];
  assign t[26] = t[32] ^ t[11];
  assign t[27] = x[0] ? x[22] : t[28];
  assign t[28] = ~(t[29] ^ t[37]);
  assign t[29] = ~t[30];
  assign t[2] = ~t[3];
  assign t[30] = ~(t[23]);
  assign t[31] = (t[38] & ~t[39]) | (~t[38] & t[39]);
  assign t[32] = (t[40] & ~t[41]) | (~t[40] & t[41]);
  assign t[33] = (t[40] & ~t[43] & ~t[45]) | (~t[42] & t[43] & ~t[44]) | (~t[40] & ~t[43] & t[45]) | (t[42] & t[43] & t[44]);
  assign t[34] = (t[40] & ~t[44]) | (~t[40] & t[44]);
  assign t[35] = (t[40] & ~t[43] & ~t[44]) | (~t[42] & t[43] & ~t[45]) | (~t[40] & ~t[43] & t[44]) | (t[42] & t[43] & t[45]);
  assign t[36] = (t[38] & ~t[46]) | (~t[38] & t[46]);
  assign t[37] = (t[38] & ~t[48] & ~t[39]) | (~t[47] & t[48] & ~t[49]) | (~t[38] & ~t[48] & t[39]) | (t[47] & t[48] & t[49]);
  assign t[38] = t[50] ^ x[7];
  assign t[39] = t[51] ^ x[8];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[52] ^ x[14];
  assign t[41] = t[53] ^ x[15];
  assign t[42] = t[54] ^ x[16];
  assign t[43] = t[55] ^ x[17];
  assign t[44] = t[56] ^ x[18];
  assign t[45] = t[57] ^ x[19];
  assign t[46] = t[58] ^ x[21];
  assign t[47] = t[59] ^ x[23];
  assign t[48] = t[60] ^ x[24];
  assign t[49] = t[61] ^ x[25];
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[62] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[63] & ~t[64] & ~t[67] & ~t[68]) | (~t[62] & t[63] & t[64] & t[65] & ~t[68]) | (~t[62] & t[63] & t[66] & t[67] & ~t[68]) | (t[62] & ~t[64] & ~t[66] & t[68]) | (~t[62] & t[64] & t[66] & t[68]);
  assign t[51] = (t[62] & t[63] & ~t[64] & ~t[66] & t[67] & ~t[68]) | (t[62] & t[64] & ~t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & t[66] & ~t[67] & ~t[68]) | (~t[62] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[62] & ~t[63] & ~t[65] & t[66] & ~t[68]) | (~t[62] & ~t[64] & t[65] & t[66] & t[67]) | (t[65] & t[66] & ~t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[70] & ~t[71] & ~t[74] & ~t[75]) | (~t[69] & t[70] & t[71] & t[72] & ~t[75]) | (~t[69] & t[70] & t[73] & t[74] & ~t[75]) | (t[69] & ~t[71] & ~t[73] & t[75]) | (~t[69] & t[71] & t[73] & t[75]);
  assign t[53] = (t[69] & t[70] & ~t[71] & t[72] & ~t[73] & ~t[75]) | (t[69] & ~t[71] & ~t[72] & t[73] & ~t[74] & t[75]) | (~t[70] & t[71] & ~t[72] & ~t[73] & ~t[75]) | (~t[69] & t[71] & ~t[72] & ~t[73] & ~t[74]) | (~t[69] & ~t[70] & t[71] & ~t[74] & ~t[75]) | (~t[69] & t[71] & t[72] & ~t[73] & t[74]) | (t[71] & ~t[72] & t[74] & ~t[75]);
  assign t[54] = (t[70] & ~t[71] & ~t[72] & ~t[73] & ~t[74]) | (~t[69] & t[70] & ~t[72] & ~t[73] & ~t[75]) | (~t[69] & t[70] & ~t[71] & ~t[74] & ~t[75]) | (t[69] & ~t[70] & t[71] & t[72] & ~t[75]) | (t[69] & ~t[70] & t[73] & t[74] & ~t[75]) | (t[70] & ~t[72] & ~t[74] & t[75]) | (~t[70] & t[72] & t[74] & t[75]);
  assign t[55] = (t[69] & t[70] & t[71] & ~t[72] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & ~t[72] & ~t[73] & t[74] & t[75]) | (~t[70] & ~t[71] & t[72] & ~t[73] & ~t[74]) | (~t[69] & ~t[71] & t[72] & ~t[74] & ~t[75]) | (~t[69] & ~t[70] & t[72] & ~t[73] & ~t[75]) | (~t[70] & t[71] & t[72] & t[73] & ~t[74]) | (~t[71] & t[72] & t[73] & ~t[75]);
  assign t[56] = (t[69] & t[70] & ~t[71] & ~t[73] & t[74] & ~t[75]) | (t[69] & t[71] & ~t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & t[73] & ~t[74] & ~t[75]) | (~t[69] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[69] & ~t[70] & ~t[72] & t[73] & ~t[75]) | (~t[69] & ~t[71] & t[72] & t[73] & t[74]) | (t[72] & t[73] & ~t[74] & ~t[75]);
  assign t[57] = (t[69] & t[70] & ~t[72] & t[73] & ~t[74] & ~t[75]) | (t[70] & ~t[71] & t[72] & ~t[73] & ~t[74] & t[75]) | (~t[70] & ~t[71] & ~t[72] & ~t[73] & t[74]) | (~t[69] & ~t[72] & ~t[73] & t[74] & ~t[75]) | (~t[69] & ~t[70] & ~t[71] & t[74] & ~t[75]) | (~t[70] & t[71] & ~t[72] & t[73] & t[74]) | (t[71] & ~t[73] & t[74] & ~t[75]);
  assign t[58] = (t[62] & t[63] & ~t[64] & t[65] & ~t[66] & ~t[68]) | (t[62] & ~t[64] & ~t[65] & t[66] & ~t[67] & t[68]) | (~t[63] & t[64] & ~t[65] & ~t[66] & ~t[68]) | (~t[62] & t[64] & ~t[65] & ~t[66] & ~t[67]) | (~t[62] & ~t[63] & t[64] & ~t[67] & ~t[68]) | (~t[62] & t[64] & t[65] & ~t[66] & t[67]) | (t[64] & ~t[65] & t[67] & ~t[68]);
  assign t[59] = (t[63] & ~t[64] & ~t[65] & ~t[66] & ~t[67]) | (~t[62] & t[63] & ~t[65] & ~t[66] & ~t[68]) | (~t[62] & t[63] & ~t[64] & ~t[67] & ~t[68]) | (t[62] & ~t[63] & t[64] & t[65] & ~t[68]) | (t[62] & ~t[63] & t[66] & t[67] & ~t[68]) | (t[63] & ~t[65] & ~t[67] & t[68]) | (~t[63] & t[65] & t[67] & t[68]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[62] & t[63] & t[64] & ~t[65] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & ~t[65] & ~t[66] & t[67] & t[68]) | (~t[63] & ~t[64] & t[65] & ~t[66] & ~t[67]) | (~t[62] & ~t[64] & t[65] & ~t[67] & ~t[68]) | (~t[62] & ~t[63] & t[65] & ~t[66] & ~t[68]) | (~t[63] & t[64] & t[65] & t[66] & ~t[67]) | (~t[64] & t[65] & t[66] & ~t[68]);
  assign t[61] = (t[62] & t[63] & ~t[65] & t[66] & ~t[67] & ~t[68]) | (t[63] & ~t[64] & t[65] & ~t[66] & ~t[67] & t[68]) | (~t[63] & ~t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[65] & ~t[66] & t[67] & ~t[68]) | (~t[62] & ~t[63] & ~t[64] & t[67] & ~t[68]) | (~t[63] & t[64] & ~t[65] & t[66] & t[67]) | (t[64] & ~t[66] & t[67] & ~t[68]);
  assign t[62] = t[76] ^ x[7];
  assign t[63] = t[77] ^ x[23];
  assign t[64] = t[78] ^ x[21];
  assign t[65] = t[79] ^ x[24];
  assign t[66] = t[80] ^ x[8];
  assign t[67] = t[81] ^ x[25];
  assign t[68] = t[82] ^ x[6];
  assign t[69] = t[83] ^ x[14];
  assign t[6] = t[32] & t[10];
  assign t[70] = t[84] ^ x[16];
  assign t[71] = t[85] ^ x[15];
  assign t[72] = t[86] ^ x[17];
  assign t[73] = t[87] ^ x[18];
  assign t[74] = t[88] ^ x[19];
  assign t[75] = t[89] ^ x[13];
  assign t[76] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[77] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[78] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[79] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[81] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[82] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[83] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[84] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[85] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[86] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[87] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[88] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[89] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19] & ~t[27]) | (~t[0] & t[19] & ~t[27]) | (~t[0] & ~t[19] & t[27]) | (t[0] & t[19] & t[27]);
endmodule

module R2ind128(x, y);
 input [24:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[26]);
  assign t[12] = ~(t[25] ^ t[11]);
  assign t[13] = t[27] ^ t[26];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[25] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[25] ^ t[18];
  assign t[18] = t[26] ^ t[28];
  assign t[19] = x[0] ? x[21] : t[20];
  assign t[1] = ~(t[2] ^ t[24]);
  assign t[20] = ~(t[21] ^ t[29]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[18] ^ t[7];
  assign t[24] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[25] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[26] = (t[32] & ~t[35] & ~t[37]) | (~t[34] & t[35] & ~t[36]) | (~t[32] & ~t[35] & t[37]) | (t[34] & t[35] & t[36]);
  assign t[27] = (t[32] & ~t[36]) | (~t[32] & t[36]);
  assign t[28] = (t[32] & ~t[35] & ~t[36]) | (~t[34] & t[35] & ~t[37]) | (~t[32] & ~t[35] & t[36]) | (t[34] & t[35] & t[37]);
  assign t[29] = (t[30] & ~t[39] & ~t[40]) | (~t[38] & t[39] & ~t[31]) | (~t[30] & ~t[39] & t[40]) | (t[38] & t[39] & t[31]);
  assign t[2] = ~t[3];
  assign t[30] = t[41] ^ x[8];
  assign t[31] = t[42] ^ x[9];
  assign t[32] = t[43] ^ x[15];
  assign t[33] = t[44] ^ x[16];
  assign t[34] = t[45] ^ x[17];
  assign t[35] = t[46] ^ x[18];
  assign t[36] = t[47] ^ x[19];
  assign t[37] = t[48] ^ x[20];
  assign t[38] = t[49] ^ x[22];
  assign t[39] = t[50] ^ x[23];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[51] ^ x[24];
  assign t[41] = (t[52] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (t[52] & ~t[53] & ~t[55] & ~t[56] & ~t[58]) | (t[52] & ~t[53] & ~t[54] & ~t[57] & ~t[58]) | (~t[52] & t[53] & t[54] & t[55] & ~t[58]) | (~t[52] & t[53] & t[56] & t[57] & ~t[58]) | (t[52] & ~t[54] & ~t[56] & t[58]) | (~t[52] & t[54] & t[56] & t[58]);
  assign t[42] = (t[52] & t[53] & ~t[54] & ~t[56] & t[57] & ~t[58]) | (t[52] & t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[58]) | (~t[52] & ~t[54] & ~t[55] & t[56] & ~t[57]) | (~t[52] & ~t[53] & ~t[55] & t[56] & ~t[58]) | (~t[52] & ~t[54] & t[55] & t[56] & t[57]) | (t[55] & t[56] & ~t[57] & ~t[58]);
  assign t[43] = (t[59] & ~t[61] & ~t[62] & ~t[63] & ~t[64]) | (t[59] & ~t[60] & ~t[62] & ~t[63] & ~t[65]) | (t[59] & ~t[60] & ~t[61] & ~t[64] & ~t[65]) | (~t[59] & t[60] & t[61] & t[62] & ~t[65]) | (~t[59] & t[60] & t[63] & t[64] & ~t[65]) | (t[59] & ~t[61] & ~t[63] & t[65]) | (~t[59] & t[61] & t[63] & t[65]);
  assign t[44] = (t[59] & t[60] & ~t[61] & t[62] & ~t[63] & ~t[65]) | (t[59] & ~t[61] & ~t[62] & t[63] & ~t[64] & t[65]) | (~t[60] & t[61] & ~t[62] & ~t[63] & ~t[65]) | (~t[59] & t[61] & ~t[62] & ~t[63] & ~t[64]) | (~t[59] & ~t[60] & t[61] & ~t[64] & ~t[65]) | (~t[59] & t[61] & t[62] & ~t[63] & t[64]) | (t[61] & ~t[62] & t[64] & ~t[65]);
  assign t[45] = (t[60] & ~t[61] & ~t[62] & ~t[63] & ~t[64]) | (~t[59] & t[60] & ~t[62] & ~t[63] & ~t[65]) | (~t[59] & t[60] & ~t[61] & ~t[64] & ~t[65]) | (t[59] & ~t[60] & t[61] & t[62] & ~t[65]) | (t[59] & ~t[60] & t[63] & t[64] & ~t[65]) | (t[60] & ~t[62] & ~t[64] & t[65]) | (~t[60] & t[62] & t[64] & t[65]);
  assign t[46] = (t[59] & t[60] & t[61] & ~t[62] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[62] & ~t[63] & t[64] & t[65]) | (~t[60] & ~t[61] & t[62] & ~t[63] & ~t[64]) | (~t[59] & ~t[61] & t[62] & ~t[64] & ~t[65]) | (~t[59] & ~t[60] & t[62] & ~t[63] & ~t[65]) | (~t[60] & t[61] & t[62] & t[63] & ~t[64]) | (~t[61] & t[62] & t[63] & ~t[65]);
  assign t[47] = (t[59] & t[60] & ~t[61] & ~t[63] & t[64] & ~t[65]) | (t[59] & t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[65]) | (~t[59] & ~t[61] & ~t[62] & t[63] & ~t[64]) | (~t[59] & ~t[60] & ~t[62] & t[63] & ~t[65]) | (~t[59] & ~t[61] & t[62] & t[63] & t[64]) | (t[62] & t[63] & ~t[64] & ~t[65]);
  assign t[48] = (t[59] & t[60] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[61] & ~t[62] & ~t[63] & t[64]) | (~t[59] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[59] & ~t[60] & ~t[61] & t[64] & ~t[65]) | (~t[60] & t[61] & ~t[62] & t[63] & t[64]) | (t[61] & ~t[63] & t[64] & ~t[65]);
  assign t[49] = (t[53] & ~t[54] & ~t[55] & ~t[56] & ~t[57]) | (~t[52] & t[53] & ~t[55] & ~t[56] & ~t[58]) | (~t[52] & t[53] & ~t[54] & ~t[57] & ~t[58]) | (t[52] & ~t[53] & t[54] & t[55] & ~t[58]) | (t[52] & ~t[53] & t[56] & t[57] & ~t[58]) | (t[53] & ~t[55] & ~t[57] & t[58]) | (~t[53] & t[55] & t[57] & t[58]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[52] & t[53] & t[54] & ~t[55] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[55] & ~t[56] & t[57] & t[58]) | (~t[53] & ~t[54] & t[55] & ~t[56] & ~t[57]) | (~t[52] & ~t[54] & t[55] & ~t[57] & ~t[58]) | (~t[52] & ~t[53] & t[55] & ~t[56] & ~t[58]) | (~t[53] & t[54] & t[55] & t[56] & ~t[57]) | (~t[54] & t[55] & t[56] & ~t[58]);
  assign t[51] = (t[52] & t[53] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[54] & ~t[55] & ~t[56] & t[57]) | (~t[52] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[52] & ~t[53] & ~t[54] & t[57] & ~t[58]) | (~t[53] & t[54] & ~t[55] & t[56] & t[57]) | (t[54] & ~t[56] & t[57] & ~t[58]);
  assign t[52] = t[66] ^ x[8];
  assign t[53] = t[67] ^ x[22];
  assign t[54] = t[68] ^ x[6];
  assign t[55] = t[69] ^ x[23];
  assign t[56] = t[70] ^ x[9];
  assign t[57] = t[71] ^ x[24];
  assign t[58] = t[72] ^ x[7];
  assign t[59] = t[73] ^ x[15];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[74] ^ x[17];
  assign t[61] = t[75] ^ x[16];
  assign t[62] = t[76] ^ x[18];
  assign t[63] = t[77] ^ x[19];
  assign t[64] = t[78] ^ x[20];
  assign t[65] = t[79] ^ x[14];
  assign t[66] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[67] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[68] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[69] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[6] = t[25] & t[10];
  assign t[70] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[71] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[72] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[73] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[74] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[75] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[76] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[77] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[78] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[79] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[7] = t[11] & t[12];
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind129(x, y);
 input [24:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[15] ^ t[16];
  assign t[11] = ~(t[27]);
  assign t[12] = ~(t[26] ^ t[11]);
  assign t[13] = t[28] ^ t[27];
  assign t[14] = ~(t[17] ^ t[8]);
  assign t[15] = t[26] ^ t[13];
  assign t[16] = t[11] & t[17];
  assign t[17] = t[26] ^ t[18];
  assign t[18] = t[27] ^ t[29];
  assign t[19] = x[0] ? x[21] : t[20];
  assign t[1] = ~(t[2] ^ t[25]);
  assign t[20] = ~(t[21] ^ t[30]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[24] ^ t[7];
  assign t[24] = t[13] ^ t[16];
  assign t[25] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[26] = (t[33] & ~t[34]) | (~t[33] & t[34]);
  assign t[27] = (t[33] & ~t[36] & ~t[38]) | (~t[35] & t[36] & ~t[37]) | (~t[33] & ~t[36] & t[38]) | (t[35] & t[36] & t[37]);
  assign t[28] = (t[33] & ~t[37]) | (~t[33] & t[37]);
  assign t[29] = (t[33] & ~t[36] & ~t[37]) | (~t[35] & t[36] & ~t[38]) | (~t[33] & ~t[36] & t[37]) | (t[35] & t[36] & t[38]);
  assign t[2] = ~t[3];
  assign t[30] = (t[31] & ~t[40] & ~t[32]) | (~t[39] & t[40] & ~t[41]) | (~t[31] & ~t[40] & t[32]) | (t[39] & t[40] & t[41]);
  assign t[31] = t[42] ^ x[8];
  assign t[32] = t[43] ^ x[9];
  assign t[33] = t[44] ^ x[15];
  assign t[34] = t[45] ^ x[16];
  assign t[35] = t[46] ^ x[17];
  assign t[36] = t[47] ^ x[18];
  assign t[37] = t[48] ^ x[19];
  assign t[38] = t[49] ^ x[20];
  assign t[39] = t[50] ^ x[22];
  assign t[3] = t[4] ^ t[5];
  assign t[40] = t[51] ^ x[23];
  assign t[41] = t[52] ^ x[24];
  assign t[42] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[43] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[45] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[51] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[8];
  assign t[54] = t[68] ^ x[22];
  assign t[55] = t[69] ^ x[6];
  assign t[56] = t[70] ^ x[23];
  assign t[57] = t[71] ^ x[9];
  assign t[58] = t[72] ^ x[24];
  assign t[59] = t[73] ^ x[7];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[74] ^ x[15];
  assign t[61] = t[75] ^ x[17];
  assign t[62] = t[76] ^ x[16];
  assign t[63] = t[77] ^ x[18];
  assign t[64] = t[78] ^ x[19];
  assign t[65] = t[79] ^ x[20];
  assign t[66] = t[80] ^ x[14];
  assign t[67] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[68] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[69] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[6] = t[26] & t[10];
  assign t[70] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[71] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[72] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[73] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[74] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[75] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[76] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[77] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[78] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[79] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[7] = t[11] & t[12];
  assign t[80] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[8] = t[13] ^ t[11];
  assign t[9] = t[14] ^ t[7];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind130(x, y);
 input [24:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[26] ^ t[27];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[27]);
  assign t[13] = ~(t[25] ^ t[12]);
  assign t[14] = t[25] & t[16];
  assign t[15] = t[25] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[27] ^ t[28];
  assign t[18] = t[25] ^ t[10];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[24]);
  assign t[20] = ~(t[21] ^ t[29]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[23]);
  assign t[23] = t[17] ^ t[7];
  assign t[24] = (t[30] & ~t[31]) | (~t[30] & t[31]);
  assign t[25] = (t[32] & ~t[33]) | (~t[32] & t[33]);
  assign t[26] = (t[32] & ~t[34]) | (~t[32] & t[34]);
  assign t[27] = (t[32] & ~t[36] & ~t[37]) | (~t[35] & t[36] & ~t[34]) | (~t[32] & ~t[36] & t[37]) | (t[35] & t[36] & t[34]);
  assign t[28] = (t[32] & ~t[36] & ~t[34]) | (~t[35] & t[36] & ~t[37]) | (~t[32] & ~t[36] & t[34]) | (t[35] & t[36] & t[37]);
  assign t[29] = (t[30] & ~t[39] & ~t[41]) | (~t[38] & t[39] & ~t[40]) | (~t[30] & ~t[39] & t[41]) | (t[38] & t[39] & t[40]);
  assign t[2] = ~t[3];
  assign t[30] = t[42] ^ x[7];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[16];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[18];
  assign t[37] = t[49] ^ x[19];
  assign t[38] = t[50] ^ x[21];
  assign t[39] = t[51] ^ x[22];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[52] ^ x[23];
  assign t[41] = t[53] ^ x[24];
  assign t[42] = (t[54] & ~t[56] & ~t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[57] & ~t[58] & ~t[60]) | (t[54] & ~t[55] & ~t[56] & ~t[59] & ~t[60]) | (~t[54] & t[55] & t[56] & t[57] & ~t[60]) | (~t[54] & t[55] & t[58] & t[59] & ~t[60]) | (t[54] & ~t[56] & ~t[58] & t[60]) | (~t[54] & t[56] & t[58] & t[60]);
  assign t[43] = (t[54] & t[55] & ~t[56] & t[57] & ~t[58] & ~t[60]) | (t[54] & ~t[56] & ~t[57] & t[58] & ~t[59] & t[60]) | (~t[55] & t[56] & ~t[57] & ~t[58] & ~t[60]) | (~t[54] & t[56] & ~t[57] & ~t[58] & ~t[59]) | (~t[54] & ~t[55] & t[56] & ~t[59] & ~t[60]) | (~t[54] & t[56] & t[57] & ~t[58] & t[59]) | (t[56] & ~t[57] & t[59] & ~t[60]);
  assign t[44] = (t[61] & ~t[63] & ~t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[64] & ~t[65] & ~t[67]) | (t[61] & ~t[62] & ~t[63] & ~t[66] & ~t[67]) | (~t[61] & t[62] & t[63] & t[64] & ~t[67]) | (~t[61] & t[62] & t[65] & t[66] & ~t[67]) | (t[61] & ~t[63] & ~t[65] & t[67]) | (~t[61] & t[63] & t[65] & t[67]);
  assign t[45] = (t[61] & t[62] & ~t[63] & t[64] & ~t[65] & ~t[67]) | (t[61] & ~t[63] & ~t[64] & t[65] & ~t[66] & t[67]) | (~t[62] & t[63] & ~t[64] & ~t[65] & ~t[67]) | (~t[61] & t[63] & ~t[64] & ~t[65] & ~t[66]) | (~t[61] & ~t[62] & t[63] & ~t[66] & ~t[67]) | (~t[61] & t[63] & t[64] & ~t[65] & t[66]) | (t[63] & ~t[64] & t[66] & ~t[67]);
  assign t[46] = (t[61] & t[62] & ~t[63] & ~t[65] & t[66] & ~t[67]) | (t[61] & t[63] & ~t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[63] & t[65] & ~t[66] & ~t[67]) | (~t[61] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[61] & ~t[62] & ~t[64] & t[65] & ~t[67]) | (~t[61] & ~t[63] & t[64] & t[65] & t[66]) | (t[64] & t[65] & ~t[66] & ~t[67]);
  assign t[47] = (t[62] & ~t[63] & ~t[64] & ~t[65] & ~t[66]) | (~t[61] & t[62] & ~t[64] & ~t[65] & ~t[67]) | (~t[61] & t[62] & ~t[63] & ~t[66] & ~t[67]) | (t[61] & ~t[62] & t[63] & t[64] & ~t[67]) | (t[61] & ~t[62] & t[65] & t[66] & ~t[67]) | (t[62] & ~t[64] & ~t[66] & t[67]) | (~t[62] & t[64] & t[66] & t[67]);
  assign t[48] = (t[61] & t[62] & t[63] & ~t[64] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & ~t[64] & ~t[65] & t[66] & t[67]) | (~t[62] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (~t[61] & ~t[63] & t[64] & ~t[66] & ~t[67]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[67]) | (~t[62] & t[63] & t[64] & t[65] & ~t[66]) | (~t[63] & t[64] & t[65] & ~t[67]);
  assign t[49] = (t[61] & t[62] & ~t[64] & t[65] & ~t[66] & ~t[67]) | (t[62] & ~t[63] & t[64] & ~t[65] & ~t[66] & t[67]) | (~t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[64] & ~t[65] & t[66] & ~t[67]) | (~t[61] & ~t[62] & ~t[63] & t[66] & ~t[67]) | (~t[62] & t[63] & ~t[64] & t[65] & t[66]) | (t[63] & ~t[65] & t[66] & ~t[67]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[55] & ~t[56] & ~t[57] & ~t[58] & ~t[59]) | (~t[54] & t[55] & ~t[57] & ~t[58] & ~t[60]) | (~t[54] & t[55] & ~t[56] & ~t[59] & ~t[60]) | (t[54] & ~t[55] & t[56] & t[57] & ~t[60]) | (t[54] & ~t[55] & t[58] & t[59] & ~t[60]) | (t[55] & ~t[57] & ~t[59] & t[60]) | (~t[55] & t[57] & t[59] & t[60]);
  assign t[51] = (t[54] & t[55] & t[56] & ~t[57] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & ~t[57] & ~t[58] & t[59] & t[60]) | (~t[55] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (~t[54] & ~t[56] & t[57] & ~t[59] & ~t[60]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[60]) | (~t[55] & t[56] & t[57] & t[58] & ~t[59]) | (~t[56] & t[57] & t[58] & ~t[60]);
  assign t[52] = (t[54] & t[55] & ~t[56] & ~t[58] & t[59] & ~t[60]) | (t[54] & t[56] & ~t[57] & ~t[58] & ~t[59] & t[60]) | (~t[55] & ~t[56] & t[58] & ~t[59] & ~t[60]) | (~t[54] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[54] & ~t[55] & ~t[57] & t[58] & ~t[60]) | (~t[54] & ~t[56] & t[57] & t[58] & t[59]) | (t[57] & t[58] & ~t[59] & ~t[60]);
  assign t[53] = (t[54] & t[55] & ~t[57] & t[58] & ~t[59] & ~t[60]) | (t[55] & ~t[56] & t[57] & ~t[58] & ~t[59] & t[60]) | (~t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[57] & ~t[58] & t[59] & ~t[60]) | (~t[54] & ~t[55] & ~t[56] & t[59] & ~t[60]) | (~t[55] & t[56] & ~t[57] & t[58] & t[59]) | (t[56] & ~t[58] & t[59] & ~t[60]);
  assign t[54] = t[68] ^ x[7];
  assign t[55] = t[69] ^ x[21];
  assign t[56] = t[70] ^ x[8];
  assign t[57] = t[71] ^ x[22];
  assign t[58] = t[72] ^ x[23];
  assign t[59] = t[73] ^ x[24];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[74] ^ x[6];
  assign t[61] = t[75] ^ x[14];
  assign t[62] = t[76] ^ x[17];
  assign t[63] = t[77] ^ x[15];
  assign t[64] = t[78] ^ x[18];
  assign t[65] = t[79] ^ x[16];
  assign t[66] = t[80] ^ x[19];
  assign t[67] = t[81] ^ x[13];
  assign t[68] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[69] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[71] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[72] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[73] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[74] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[75] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[76] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[77] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[78] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[79] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[7] = t[12] & t[13];
  assign t[80] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[81] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[25] ^ t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind131(x, y);
 input [24:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = t[25] ^ t[26];
  assign t[11] = t[12] & t[15];
  assign t[12] = ~(t[26]);
  assign t[13] = ~(t[24] ^ t[12]);
  assign t[14] = t[24] & t[16];
  assign t[15] = t[24] ^ t[17];
  assign t[16] = t[18] ^ t[11];
  assign t[17] = t[26] ^ t[27];
  assign t[18] = t[24] ^ t[10];
  assign t[19] = x[0] ? x[20] : t[20];
  assign t[1] = ~(t[2] ^ t[23]);
  assign t[20] = ~(t[21] ^ t[28]);
  assign t[21] = ~t[22];
  assign t[22] = ~(t[4]);
  assign t[23] = (t[29] & ~t[30]) | (~t[29] & t[30]);
  assign t[24] = (t[31] & ~t[32]) | (~t[31] & t[32]);
  assign t[25] = (t[31] & ~t[33]) | (~t[31] & t[33]);
  assign t[26] = (t[31] & ~t[35] & ~t[36]) | (~t[34] & t[35] & ~t[33]) | (~t[31] & ~t[35] & t[36]) | (t[34] & t[35] & t[33]);
  assign t[27] = (t[31] & ~t[35] & ~t[33]) | (~t[34] & t[35] & ~t[36]) | (~t[31] & ~t[35] & t[33]) | (t[34] & t[35] & t[36]);
  assign t[28] = (t[29] & ~t[38] & ~t[39]) | (~t[37] & t[38] & ~t[40]) | (~t[29] & ~t[38] & t[39]) | (t[37] & t[38] & t[40]);
  assign t[29] = t[41] ^ x[7];
  assign t[2] = ~t[3];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[14];
  assign t[32] = t[44] ^ x[15];
  assign t[33] = t[45] ^ x[16];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[18];
  assign t[36] = t[48] ^ x[19];
  assign t[37] = t[49] ^ x[21];
  assign t[38] = t[50] ^ x[22];
  assign t[39] = t[51] ^ x[23];
  assign t[3] = ~(t[4] ^ t[5]);
  assign t[40] = t[52] ^ x[24];
  assign t[41] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[42] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[44] = (t[60] & t[61] & ~t[62] & t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[62] & ~t[63] & t[64] & ~t[65] & t[66]) | (~t[61] & t[62] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[61] & t[62] & ~t[65] & ~t[66]) | (~t[60] & t[62] & t[63] & ~t[64] & t[65]) | (t[62] & ~t[63] & t[65] & ~t[66]);
  assign t[45] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[49] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[4] = t[6] ^ t[7];
  assign t[50] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[51] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[52] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[53] = t[67] ^ x[7];
  assign t[54] = t[68] ^ x[21];
  assign t[55] = t[69] ^ x[8];
  assign t[56] = t[70] ^ x[22];
  assign t[57] = t[71] ^ x[23];
  assign t[58] = t[72] ^ x[24];
  assign t[59] = t[73] ^ x[6];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = t[74] ^ x[14];
  assign t[61] = t[75] ^ x[17];
  assign t[62] = t[76] ^ x[15];
  assign t[63] = t[77] ^ x[18];
  assign t[64] = t[78] ^ x[16];
  assign t[65] = t[79] ^ x[19];
  assign t[66] = t[80] ^ x[13];
  assign t[67] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[68] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[69] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[71] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[72] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[73] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[74] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[75] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[76] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[77] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[78] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[79] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[7] = t[12] & t[13];
  assign t[80] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[8] = t[14] ^ t[7];
  assign t[9] = t[24] ^ t[12];
  assign y = (t[0] & ~t[19]) | (~t[0] & t[19]);
endmodule

module R2ind132(x, y);
 input [24:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[10] = ~(t[11] ^ t[22]);
  assign t[11] = ~t[12];
  assign t[12] = ~(t[13]);
  assign t[13] = t[14] ^ t[6];
  assign t[14] = t[15] ^ t[16];
  assign t[15] = t[23] ^ t[19];
  assign t[16] = t[7] & t[17];
  assign t[17] = t[21] ^ t[5];
  assign t[18] = (t[24] & ~t[26] & ~t[28]) | (~t[25] & t[26] & ~t[27]) | (~t[24] & ~t[26] & t[28]) | (t[25] & t[26] & t[27]);
  assign t[19] = (t[29] & ~t[31] & ~t[33]) | (~t[30] & t[31] & ~t[32]) | (~t[29] & ~t[31] & t[33]) | (t[30] & t[31] & t[32]);
  assign t[1] = ~(t[2] ^ t[18]);
  assign t[20] = (t[29] & ~t[31] & ~t[32]) | (~t[30] & t[31] & ~t[33]) | (~t[29] & ~t[31] & t[32]) | (t[30] & t[31] & t[33]);
  assign t[21] = (t[29] & ~t[34]) | (~t[29] & t[34]);
  assign t[22] = (t[24] & ~t[26] & ~t[27]) | (~t[25] & t[26] & ~t[28]) | (~t[24] & ~t[26] & t[27]) | (t[25] & t[26] & t[28]);
  assign t[23] = (t[29] & ~t[32]) | (~t[29] & t[32]);
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[9];
  assign t[26] = t[37] ^ x[10];
  assign t[27] = t[38] ^ x[11];
  assign t[28] = t[39] ^ x[12];
  assign t[29] = t[40] ^ x[18];
  assign t[2] = ~t[3];
  assign t[30] = t[41] ^ x[19];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[23];
  assign t[35] = (t[46] & ~t[48] & ~t[49] & ~t[50] & ~t[51]) | (t[46] & ~t[47] & ~t[49] & ~t[50] & ~t[52]) | (t[46] & ~t[47] & ~t[48] & ~t[51] & ~t[52]) | (~t[46] & t[47] & t[48] & t[49] & ~t[52]) | (~t[46] & t[47] & t[50] & t[51] & ~t[52]) | (t[46] & ~t[48] & ~t[50] & t[52]) | (~t[46] & t[48] & t[50] & t[52]);
  assign t[36] = (t[47] & ~t[48] & ~t[49] & ~t[50] & ~t[51]) | (~t[46] & t[47] & ~t[49] & ~t[50] & ~t[52]) | (~t[46] & t[47] & ~t[48] & ~t[51] & ~t[52]) | (t[46] & ~t[47] & t[48] & t[49] & ~t[52]) | (t[46] & ~t[47] & t[50] & t[51] & ~t[52]) | (t[47] & ~t[49] & ~t[51] & t[52]) | (~t[47] & t[49] & t[51] & t[52]);
  assign t[37] = (t[46] & t[47] & t[48] & ~t[49] & ~t[51] & ~t[52]) | (t[47] & ~t[48] & ~t[49] & ~t[50] & t[51] & t[52]) | (~t[47] & ~t[48] & t[49] & ~t[50] & ~t[51]) | (~t[46] & ~t[48] & t[49] & ~t[51] & ~t[52]) | (~t[46] & ~t[47] & t[49] & ~t[50] & ~t[52]) | (~t[47] & t[48] & t[49] & t[50] & ~t[51]) | (~t[48] & t[49] & t[50] & ~t[52]);
  assign t[38] = (t[46] & t[47] & ~t[48] & ~t[50] & t[51] & ~t[52]) | (t[46] & t[48] & ~t[49] & ~t[50] & ~t[51] & t[52]) | (~t[47] & ~t[48] & t[50] & ~t[51] & ~t[52]) | (~t[46] & ~t[48] & ~t[49] & t[50] & ~t[51]) | (~t[46] & ~t[47] & ~t[49] & t[50] & ~t[52]) | (~t[46] & ~t[48] & t[49] & t[50] & t[51]) | (t[49] & t[50] & ~t[51] & ~t[52]);
  assign t[39] = (t[46] & t[47] & ~t[49] & t[50] & ~t[51] & ~t[52]) | (t[47] & ~t[48] & t[49] & ~t[50] & ~t[51] & t[52]) | (~t[47] & ~t[48] & ~t[49] & ~t[50] & t[51]) | (~t[46] & ~t[49] & ~t[50] & t[51] & ~t[52]) | (~t[46] & ~t[47] & ~t[48] & t[51] & ~t[52]) | (~t[47] & t[48] & ~t[49] & t[50] & t[51]) | (t[48] & ~t[50] & t[51] & ~t[52]);
  assign t[3] = ~(t[4]);
  assign t[40] = (t[53] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (t[53] & ~t[54] & ~t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[54] & ~t[55] & ~t[58] & ~t[59]) | (~t[53] & t[54] & t[55] & t[56] & ~t[59]) | (~t[53] & t[54] & t[57] & t[58] & ~t[59]) | (t[53] & ~t[55] & ~t[57] & t[59]) | (~t[53] & t[55] & t[57] & t[59]);
  assign t[41] = (t[54] & ~t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & t[54] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[54] & ~t[55] & ~t[58] & ~t[59]) | (t[53] & ~t[54] & t[55] & t[56] & ~t[59]) | (t[53] & ~t[54] & t[57] & t[58] & ~t[59]) | (t[54] & ~t[56] & ~t[58] & t[59]) | (~t[54] & t[56] & t[58] & t[59]);
  assign t[42] = (t[53] & t[54] & t[55] & ~t[56] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & ~t[56] & ~t[57] & t[58] & t[59]) | (~t[54] & ~t[55] & t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[55] & t[56] & ~t[58] & ~t[59]) | (~t[53] & ~t[54] & t[56] & ~t[57] & ~t[59]) | (~t[54] & t[55] & t[56] & t[57] & ~t[58]) | (~t[55] & t[56] & t[57] & ~t[59]);
  assign t[43] = (t[53] & t[54] & ~t[55] & ~t[57] & t[58] & ~t[59]) | (t[53] & t[55] & ~t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & t[57] & ~t[58] & ~t[59]) | (~t[53] & ~t[55] & ~t[56] & t[57] & ~t[58]) | (~t[53] & ~t[54] & ~t[56] & t[57] & ~t[59]) | (~t[53] & ~t[55] & t[56] & t[57] & t[58]) | (t[56] & t[57] & ~t[58] & ~t[59]);
  assign t[44] = (t[53] & t[54] & ~t[56] & t[57] & ~t[58] & ~t[59]) | (t[54] & ~t[55] & t[56] & ~t[57] & ~t[58] & t[59]) | (~t[54] & ~t[55] & ~t[56] & ~t[57] & t[58]) | (~t[53] & ~t[56] & ~t[57] & t[58] & ~t[59]) | (~t[53] & ~t[54] & ~t[55] & t[58] & ~t[59]) | (~t[54] & t[55] & ~t[56] & t[57] & t[58]) | (t[55] & ~t[57] & t[58] & ~t[59]);
  assign t[45] = (t[53] & t[54] & ~t[55] & t[56] & ~t[57] & ~t[59]) | (t[53] & ~t[55] & ~t[56] & t[57] & ~t[58] & t[59]) | (~t[54] & t[55] & ~t[56] & ~t[57] & ~t[59]) | (~t[53] & t[55] & ~t[56] & ~t[57] & ~t[58]) | (~t[53] & ~t[54] & t[55] & ~t[58] & ~t[59]) | (~t[53] & t[55] & t[56] & ~t[57] & t[58]) | (t[55] & ~t[56] & t[58] & ~t[59]);
  assign t[46] = t[60] ^ x[8];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[6];
  assign t[49] = t[63] ^ x[10];
  assign t[4] = t[5] ^ t[6];
  assign t[50] = t[64] ^ x[11];
  assign t[51] = t[65] ^ x[12];
  assign t[52] = t[66] ^ x[7];
  assign t[53] = t[67] ^ x[18];
  assign t[54] = t[68] ^ x[19];
  assign t[55] = t[69] ^ x[23];
  assign t[56] = t[70] ^ x[20];
  assign t[57] = t[71] ^ x[21];
  assign t[58] = t[72] ^ x[22];
  assign t[59] = t[73] ^ x[17];
  assign t[5] = t[19] ^ t[20];
  assign t[60] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[61] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[62] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[63] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[64] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[65] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[66] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[67] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[68] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[69] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[6] = t[7] & t[8];
  assign t[70] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[71] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[72] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[73] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[7] = ~(t[19]);
  assign t[8] = ~(t[21] ^ t[7]);
  assign t[9] = x[0] ? x[24] : t[10];
  assign y = (t[0] & ~t[9]) | (~t[0] & t[9]);
endmodule

module R2ind133(x, y);
 input [49:0] x;
 output y;

 wire [153:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[135] ^ x[23];
  assign t[101] = t[136] ^ x[25];
  assign t[102] = t[137] ^ x[26];
  assign t[103] = t[138] ^ x[27];
  assign t[104] = t[139] ^ x[21];
  assign t[105] = t[140] ^ x[36];
  assign t[106] = t[141] ^ x[31];
  assign t[107] = t[142] ^ x[32];
  assign t[108] = t[143] ^ x[33];
  assign t[109] = t[144] ^ x[37];
  assign t[10] = t[15] ^ t[13];
  assign t[110] = t[145] ^ x[34];
  assign t[111] = t[146] ^ x[35];
  assign t[112] = t[147] ^ x[48];
  assign t[113] = t[148] ^ x[43];
  assign t[114] = t[149] ^ x[44];
  assign t[115] = t[150] ^ x[45];
  assign t[116] = t[151] ^ x[49];
  assign t[117] = t[152] ^ x[46];
  assign t[118] = t[153] ^ x[47];
  assign t[119] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[11] = t[16] ^ t[9];
  assign t[120] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[121] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[122] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[123] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[124] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[125] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[126] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[127] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[128] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[129] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[12] = t[17] ^ t[18];
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[133] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[134] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[135] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[136] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[137] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[138] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[139] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[13] = ~(t[41]);
  assign t[140] = (x[30] & ~1'b0 & ~1'b0) | (~x[30] & 1'b0 & ~1'b0) | (~x[30] & ~1'b0 & 1'b0) | (x[30] & 1'b0 & 1'b0);
  assign t[141] = (x[30] & ~1'b0 & ~1'b0) | (~x[30] & 1'b0 & ~1'b0) | (~x[30] & ~1'b0 & 1'b0) | (x[30] & 1'b0 & 1'b0);
  assign t[142] = (x[30] & ~1'b0) | (~x[30] & 1'b0);
  assign t[143] = (x[30] & ~1'b0) | (~x[30] & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[147] = (x[42] & ~1'b0 & ~1'b0) | (~x[42] & 1'b0 & ~1'b0) | (~x[42] & ~1'b0 & 1'b0) | (x[42] & 1'b0 & 1'b0);
  assign t[148] = (x[42] & ~1'b0 & ~1'b0) | (~x[42] & 1'b0 & ~1'b0) | (~x[42] & ~1'b0 & 1'b0) | (x[42] & 1'b0 & 1'b0);
  assign t[149] = (x[42] & ~1'b0) | (~x[42] & 1'b0);
  assign t[14] = ~(t[40] ^ t[13]);
  assign t[150] = (x[42] & ~1'b0) | (~x[42] & 1'b0);
  assign t[151] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[152] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[153] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = t[42] ^ t[41];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[40] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[40] ^ t[20];
  assign t[1] = ~(t[2] ^ t[38]);
  assign t[20] = t[41] ^ t[43];
  assign t[21] = x[0] ? x[28] : t[22];
  assign t[22] = ~(t[23] ^ t[44]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[45]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = t[29] ^ t[9];
  assign t[28] = t[6] ^ t[30];
  assign t[29] = t[15] ^ t[18];
  assign t[2] = ~t[3];
  assign t[30] = t[40] ^ t[13];
  assign t[31] = x[0] ? x[38] : t[32];
  assign t[32] = ~(t[33] ^ t[46]);
  assign t[33] = ~t[34];
  assign t[34] = ~(t[35] ^ t[47]);
  assign t[35] = ~t[36];
  assign t[36] = ~(t[37]);
  assign t[37] = t[20] ^ t[9];
  assign t[38] = (t[48] & ~t[49]) | (~t[48] & t[49]);
  assign t[39] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[3] = ~(t[4] ^ t[39]);
  assign t[40] = (t[52] & ~t[53]) | (~t[52] & t[53]);
  assign t[41] = (t[52] & ~t[55] & ~t[57]) | (~t[54] & t[55] & ~t[56]) | (~t[52] & ~t[55] & t[57]) | (t[54] & t[55] & t[56]);
  assign t[42] = (t[52] & ~t[56]) | (~t[52] & t[56]);
  assign t[43] = (t[52] & ~t[55] & ~t[56]) | (~t[54] & t[55] & ~t[57]) | (~t[52] & ~t[55] & t[56]) | (t[54] & t[55] & t[57]);
  assign t[44] = (t[48] & ~t[58]) | (~t[48] & t[58]);
  assign t[45] = (t[59] & ~t[60]) | (~t[59] & t[60]);
  assign t[46] = (t[48] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[49]) | (~t[48] & ~t[62] & t[63]) | (t[61] & t[62] & t[49]);
  assign t[47] = (t[64] & ~t[65]) | (~t[64] & t[65]);
  assign t[48] = t[66] ^ x[7];
  assign t[49] = t[67] ^ x[8];
  assign t[4] = ~t[5];
  assign t[50] = t[68] ^ x[15];
  assign t[51] = t[69] ^ x[16];
  assign t[52] = t[70] ^ x[22];
  assign t[53] = t[71] ^ x[23];
  assign t[54] = t[72] ^ x[24];
  assign t[55] = t[73] ^ x[25];
  assign t[56] = t[74] ^ x[26];
  assign t[57] = t[75] ^ x[27];
  assign t[58] = t[76] ^ x[29];
  assign t[59] = t[77] ^ x[36];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[78] ^ x[37];
  assign t[61] = t[79] ^ x[39];
  assign t[62] = t[80] ^ x[40];
  assign t[63] = t[81] ^ x[41];
  assign t[64] = t[82] ^ x[48];
  assign t[65] = t[83] ^ x[49];
  assign t[66] = (t[84] & ~t[86] & ~t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[87] & ~t[88] & ~t[90]) | (t[84] & ~t[85] & ~t[86] & ~t[89] & ~t[90]) | (~t[84] & t[85] & t[86] & t[87] & ~t[90]) | (~t[84] & t[85] & t[88] & t[89] & ~t[90]) | (t[84] & ~t[86] & ~t[88] & t[90]) | (~t[84] & t[86] & t[88] & t[90]);
  assign t[67] = (t[84] & t[85] & ~t[86] & ~t[88] & t[89] & ~t[90]) | (t[84] & t[86] & ~t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[86] & t[88] & ~t[89] & ~t[90]) | (~t[84] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[84] & ~t[85] & ~t[87] & t[88] & ~t[90]) | (~t[84] & ~t[86] & t[87] & t[88] & t[89]) | (t[87] & t[88] & ~t[89] & ~t[90]);
  assign t[68] = (t[91] & ~t[93] & ~t[94] & ~t[95] & ~t[96]) | (t[91] & ~t[92] & ~t[94] & ~t[95] & ~t[97]) | (t[91] & ~t[92] & ~t[93] & ~t[96] & ~t[97]) | (~t[91] & t[92] & t[93] & t[94] & ~t[97]) | (~t[91] & t[92] & t[95] & t[96] & ~t[97]) | (t[91] & ~t[93] & ~t[95] & t[97]) | (~t[91] & t[93] & t[95] & t[97]);
  assign t[69] = (t[91] & t[92] & ~t[93] & ~t[95] & t[96] & ~t[97]) | (t[91] & t[93] & ~t[94] & ~t[95] & ~t[96] & t[97]) | (~t[92] & ~t[93] & t[95] & ~t[96] & ~t[97]) | (~t[91] & ~t[93] & ~t[94] & t[95] & ~t[96]) | (~t[91] & ~t[92] & ~t[94] & t[95] & ~t[97]) | (~t[91] & ~t[93] & t[94] & t[95] & t[96]) | (t[94] & t[95] & ~t[96] & ~t[97]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (t[98] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[99] & ~t[100] & ~t[103] & ~t[104]) | (~t[98] & t[99] & t[100] & t[101] & ~t[104]) | (~t[98] & t[99] & t[102] & t[103] & ~t[104]) | (t[98] & ~t[100] & ~t[102] & t[104]) | (~t[98] & t[100] & t[102] & t[104]);
  assign t[71] = (t[98] & t[99] & ~t[100] & t[101] & ~t[102] & ~t[104]) | (t[98] & ~t[100] & ~t[101] & t[102] & ~t[103] & t[104]) | (~t[99] & t[100] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[99] & t[100] & ~t[103] & ~t[104]) | (~t[98] & t[100] & t[101] & ~t[102] & t[103]) | (t[100] & ~t[101] & t[103] & ~t[104]);
  assign t[72] = (t[99] & ~t[100] & ~t[101] & ~t[102] & ~t[103]) | (~t[98] & t[99] & ~t[101] & ~t[102] & ~t[104]) | (~t[98] & t[99] & ~t[100] & ~t[103] & ~t[104]) | (t[98] & ~t[99] & t[100] & t[101] & ~t[104]) | (t[98] & ~t[99] & t[102] & t[103] & ~t[104]) | (t[99] & ~t[101] & ~t[103] & t[104]) | (~t[99] & t[101] & t[103] & t[104]);
  assign t[73] = (t[98] & t[99] & t[100] & ~t[101] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & ~t[101] & ~t[102] & t[103] & t[104]) | (~t[99] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (~t[98] & ~t[100] & t[101] & ~t[103] & ~t[104]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[104]) | (~t[99] & t[100] & t[101] & t[102] & ~t[103]) | (~t[100] & t[101] & t[102] & ~t[104]);
  assign t[74] = (t[98] & t[99] & ~t[100] & ~t[102] & t[103] & ~t[104]) | (t[98] & t[100] & ~t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & t[102] & ~t[103] & ~t[104]) | (~t[98] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[98] & ~t[99] & ~t[101] & t[102] & ~t[104]) | (~t[98] & ~t[100] & t[101] & t[102] & t[103]) | (t[101] & t[102] & ~t[103] & ~t[104]);
  assign t[75] = (t[98] & t[99] & ~t[101] & t[102] & ~t[103] & ~t[104]) | (t[99] & ~t[100] & t[101] & ~t[102] & ~t[103] & t[104]) | (~t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[101] & ~t[102] & t[103] & ~t[104]) | (~t[98] & ~t[99] & ~t[100] & t[103] & ~t[104]) | (~t[99] & t[100] & ~t[101] & t[102] & t[103]) | (t[100] & ~t[102] & t[103] & ~t[104]);
  assign t[76] = (t[84] & t[85] & ~t[86] & t[87] & ~t[88] & ~t[90]) | (t[84] & ~t[86] & ~t[87] & t[88] & ~t[89] & t[90]) | (~t[85] & t[86] & ~t[87] & ~t[88] & ~t[90]) | (~t[84] & t[86] & ~t[87] & ~t[88] & ~t[89]) | (~t[84] & ~t[85] & t[86] & ~t[89] & ~t[90]) | (~t[84] & t[86] & t[87] & ~t[88] & t[89]) | (t[86] & ~t[87] & t[89] & ~t[90]);
  assign t[77] = (t[105] & ~t[107] & ~t[108] & ~t[109] & ~t[110]) | (t[105] & ~t[106] & ~t[108] & ~t[109] & ~t[111]) | (t[105] & ~t[106] & ~t[107] & ~t[110] & ~t[111]) | (~t[105] & t[106] & t[107] & t[108] & ~t[111]) | (~t[105] & t[106] & t[109] & t[110] & ~t[111]) | (t[105] & ~t[107] & ~t[109] & t[111]) | (~t[105] & t[107] & t[109] & t[111]);
  assign t[78] = (t[105] & t[106] & ~t[107] & ~t[109] & t[110] & ~t[111]) | (t[105] & t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[111]) | (~t[105] & ~t[107] & ~t[108] & t[109] & ~t[110]) | (~t[105] & ~t[106] & ~t[108] & t[109] & ~t[111]) | (~t[105] & ~t[107] & t[108] & t[109] & t[110]) | (t[108] & t[109] & ~t[110] & ~t[111]);
  assign t[79] = (t[85] & ~t[86] & ~t[87] & ~t[88] & ~t[89]) | (~t[84] & t[85] & ~t[87] & ~t[88] & ~t[90]) | (~t[84] & t[85] & ~t[86] & ~t[89] & ~t[90]) | (t[84] & ~t[85] & t[86] & t[87] & ~t[90]) | (t[84] & ~t[85] & t[88] & t[89] & ~t[90]) | (t[85] & ~t[87] & ~t[89] & t[90]) | (~t[85] & t[87] & t[89] & t[90]);
  assign t[7] = t[10] & t[11];
  assign t[80] = (t[84] & t[85] & t[86] & ~t[87] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & ~t[87] & ~t[88] & t[89] & t[90]) | (~t[85] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (~t[84] & ~t[86] & t[87] & ~t[89] & ~t[90]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[90]) | (~t[85] & t[86] & t[87] & t[88] & ~t[89]) | (~t[86] & t[87] & t[88] & ~t[90]);
  assign t[81] = (t[84] & t[85] & ~t[87] & t[88] & ~t[89] & ~t[90]) | (t[85] & ~t[86] & t[87] & ~t[88] & ~t[89] & t[90]) | (~t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[87] & ~t[88] & t[89] & ~t[90]) | (~t[84] & ~t[85] & ~t[86] & t[89] & ~t[90]) | (~t[85] & t[86] & ~t[87] & t[88] & t[89]) | (t[86] & ~t[88] & t[89] & ~t[90]);
  assign t[82] = (t[112] & ~t[114] & ~t[115] & ~t[116] & ~t[117]) | (t[112] & ~t[113] & ~t[115] & ~t[116] & ~t[118]) | (t[112] & ~t[113] & ~t[114] & ~t[117] & ~t[118]) | (~t[112] & t[113] & t[114] & t[115] & ~t[118]) | (~t[112] & t[113] & t[116] & t[117] & ~t[118]) | (t[112] & ~t[114] & ~t[116] & t[118]) | (~t[112] & t[114] & t[116] & t[118]);
  assign t[83] = (t[112] & t[113] & ~t[114] & ~t[116] & t[117] & ~t[118]) | (t[112] & t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[118]) | (~t[112] & ~t[114] & ~t[115] & t[116] & ~t[117]) | (~t[112] & ~t[113] & ~t[115] & t[116] & ~t[118]) | (~t[112] & ~t[114] & t[115] & t[116] & t[117]) | (t[115] & t[116] & ~t[117] & ~t[118]);
  assign t[84] = t[119] ^ x[7];
  assign t[85] = t[120] ^ x[39];
  assign t[86] = t[121] ^ x[29];
  assign t[87] = t[122] ^ x[40];
  assign t[88] = t[123] ^ x[8];
  assign t[89] = t[124] ^ x[41];
  assign t[8] = t[40] & t[12];
  assign t[90] = t[125] ^ x[6];
  assign t[91] = t[126] ^ x[15];
  assign t[92] = t[127] ^ x[10];
  assign t[93] = t[128] ^ x[11];
  assign t[94] = t[129] ^ x[12];
  assign t[95] = t[130] ^ x[16];
  assign t[96] = t[131] ^ x[13];
  assign t[97] = t[132] ^ x[14];
  assign t[98] = t[133] ^ x[22];
  assign t[99] = t[134] ^ x[24];
  assign t[9] = t[13] & t[14];
  assign y = (t[0] & ~t[21] & ~t[31]) | (~t[0] & t[21] & ~t[31]) | (~t[0] & ~t[21] & t[31]) | (t[0] & t[21] & t[31]);
endmodule

module R2ind134(x, y);
 input [49:0] x;
 output y;

 wire [152:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[135] ^ x[25];
  assign t[101] = t[136] ^ x[26];
  assign t[102] = t[137] ^ x[27];
  assign t[103] = t[138] ^ x[21];
  assign t[104] = t[139] ^ x[36];
  assign t[105] = t[140] ^ x[31];
  assign t[106] = t[141] ^ x[32];
  assign t[107] = t[142] ^ x[33];
  assign t[108] = t[143] ^ x[37];
  assign t[109] = t[144] ^ x[34];
  assign t[10] = t[15] ^ t[13];
  assign t[110] = t[145] ^ x[35];
  assign t[111] = t[146] ^ x[48];
  assign t[112] = t[147] ^ x[43];
  assign t[113] = t[148] ^ x[44];
  assign t[114] = t[149] ^ x[45];
  assign t[115] = t[150] ^ x[49];
  assign t[116] = t[151] ^ x[46];
  assign t[117] = t[152] ^ x[47];
  assign t[118] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[119] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[11] = t[16] ^ t[9];
  assign t[120] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[121] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[122] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[123] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[124] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[125] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[126] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[127] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[128] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[129] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = t[17] ^ t[18];
  assign t[130] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[131] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[132] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[133] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[134] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[135] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[136] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[137] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[138] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[139] = (x[30] & ~1'b0 & ~1'b0) | (~x[30] & 1'b0 & ~1'b0) | (~x[30] & ~1'b0 & 1'b0) | (x[30] & 1'b0 & 1'b0);
  assign t[13] = ~(t[40]);
  assign t[140] = (x[30] & ~1'b0 & ~1'b0) | (~x[30] & 1'b0 & ~1'b0) | (~x[30] & ~1'b0 & 1'b0) | (x[30] & 1'b0 & 1'b0);
  assign t[141] = (x[30] & ~1'b0) | (~x[30] & 1'b0);
  assign t[142] = (x[30] & ~1'b0) | (~x[30] & 1'b0);
  assign t[143] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[144] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[145] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[146] = (x[42] & ~1'b0 & ~1'b0) | (~x[42] & 1'b0 & ~1'b0) | (~x[42] & ~1'b0 & 1'b0) | (x[42] & 1'b0 & 1'b0);
  assign t[147] = (x[42] & ~1'b0 & ~1'b0) | (~x[42] & 1'b0 & ~1'b0) | (~x[42] & ~1'b0 & 1'b0) | (x[42] & 1'b0 & 1'b0);
  assign t[148] = (x[42] & ~1'b0) | (~x[42] & 1'b0);
  assign t[149] = (x[42] & ~1'b0) | (~x[42] & 1'b0);
  assign t[14] = ~(t[39] ^ t[13]);
  assign t[150] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[151] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[152] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[15] = t[41] ^ t[40];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[39] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[39] ^ t[20];
  assign t[1] = ~(t[2] ^ t[37]);
  assign t[20] = t[40] ^ t[42];
  assign t[21] = x[0] ? x[28] : t[22];
  assign t[22] = ~(t[23] ^ t[43]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[44]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = t[29] ^ t[9];
  assign t[28] = t[6] ^ t[30];
  assign t[29] = t[15] ^ t[18];
  assign t[2] = ~t[3];
  assign t[30] = t[39] ^ t[13];
  assign t[31] = x[0] ? x[38] : t[32];
  assign t[32] = ~(t[33] ^ t[45]);
  assign t[33] = ~t[34];
  assign t[34] = ~(t[35] ^ t[46]);
  assign t[35] = ~t[36];
  assign t[36] = ~(t[27]);
  assign t[37] = (t[47] & ~t[48]) | (~t[47] & t[48]);
  assign t[38] = (t[49] & ~t[50]) | (~t[49] & t[50]);
  assign t[39] = (t[51] & ~t[52]) | (~t[51] & t[52]);
  assign t[3] = ~(t[4] ^ t[38]);
  assign t[40] = (t[51] & ~t[54] & ~t[56]) | (~t[53] & t[54] & ~t[55]) | (~t[51] & ~t[54] & t[56]) | (t[53] & t[54] & t[55]);
  assign t[41] = (t[51] & ~t[55]) | (~t[51] & t[55]);
  assign t[42] = (t[51] & ~t[54] & ~t[55]) | (~t[53] & t[54] & ~t[56]) | (~t[51] & ~t[54] & t[55]) | (t[53] & t[54] & t[56]);
  assign t[43] = (t[47] & ~t[57]) | (~t[47] & t[57]);
  assign t[44] = (t[58] & ~t[59]) | (~t[58] & t[59]);
  assign t[45] = (t[47] & ~t[61] & ~t[48]) | (~t[60] & t[61] & ~t[62]) | (~t[47] & ~t[61] & t[48]) | (t[60] & t[61] & t[62]);
  assign t[46] = (t[63] & ~t[64]) | (~t[63] & t[64]);
  assign t[47] = t[65] ^ x[7];
  assign t[48] = t[66] ^ x[8];
  assign t[49] = t[67] ^ x[15];
  assign t[4] = ~t[5];
  assign t[50] = t[68] ^ x[16];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[23];
  assign t[53] = t[71] ^ x[24];
  assign t[54] = t[72] ^ x[25];
  assign t[55] = t[73] ^ x[26];
  assign t[56] = t[74] ^ x[27];
  assign t[57] = t[75] ^ x[29];
  assign t[58] = t[76] ^ x[36];
  assign t[59] = t[77] ^ x[37];
  assign t[5] = t[6] ^ t[7];
  assign t[60] = t[78] ^ x[39];
  assign t[61] = t[79] ^ x[40];
  assign t[62] = t[80] ^ x[41];
  assign t[63] = t[81] ^ x[48];
  assign t[64] = t[82] ^ x[49];
  assign t[65] = (t[83] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[84] & ~t[85] & ~t[88] & ~t[89]) | (~t[83] & t[84] & t[85] & t[86] & ~t[89]) | (~t[83] & t[84] & t[87] & t[88] & ~t[89]) | (t[83] & ~t[85] & ~t[87] & t[89]) | (~t[83] & t[85] & t[87] & t[89]);
  assign t[66] = (t[83] & t[84] & ~t[85] & ~t[87] & t[88] & ~t[89]) | (t[83] & t[85] & ~t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & t[87] & ~t[88] & ~t[89]) | (~t[83] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[83] & ~t[84] & ~t[86] & t[87] & ~t[89]) | (~t[83] & ~t[85] & t[86] & t[87] & t[88]) | (t[86] & t[87] & ~t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[92] & ~t[93] & ~t[94] & ~t[95]) | (t[90] & ~t[91] & ~t[93] & ~t[94] & ~t[96]) | (t[90] & ~t[91] & ~t[92] & ~t[95] & ~t[96]) | (~t[90] & t[91] & t[92] & t[93] & ~t[96]) | (~t[90] & t[91] & t[94] & t[95] & ~t[96]) | (t[90] & ~t[92] & ~t[94] & t[96]) | (~t[90] & t[92] & t[94] & t[96]);
  assign t[68] = (t[90] & t[91] & ~t[92] & ~t[94] & t[95] & ~t[96]) | (t[90] & t[92] & ~t[93] & ~t[94] & ~t[95] & t[96]) | (~t[91] & ~t[92] & t[94] & ~t[95] & ~t[96]) | (~t[90] & ~t[92] & ~t[93] & t[94] & ~t[95]) | (~t[90] & ~t[91] & ~t[93] & t[94] & ~t[96]) | (~t[90] & ~t[92] & t[93] & t[94] & t[95]) | (t[93] & t[94] & ~t[95] & ~t[96]);
  assign t[69] = (t[97] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (t[97] & ~t[98] & ~t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[98] & ~t[99] & ~t[102] & ~t[103]) | (~t[97] & t[98] & t[99] & t[100] & ~t[103]) | (~t[97] & t[98] & t[101] & t[102] & ~t[103]) | (t[97] & ~t[99] & ~t[101] & t[103]) | (~t[97] & t[99] & t[101] & t[103]);
  assign t[6] = t[8] ^ t[9];
  assign t[70] = (t[97] & t[98] & ~t[99] & t[100] & ~t[101] & ~t[103]) | (t[97] & ~t[99] & ~t[100] & t[101] & ~t[102] & t[103]) | (~t[98] & t[99] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[98] & t[99] & ~t[102] & ~t[103]) | (~t[97] & t[99] & t[100] & ~t[101] & t[102]) | (t[99] & ~t[100] & t[102] & ~t[103]);
  assign t[71] = (t[98] & ~t[99] & ~t[100] & ~t[101] & ~t[102]) | (~t[97] & t[98] & ~t[100] & ~t[101] & ~t[103]) | (~t[97] & t[98] & ~t[99] & ~t[102] & ~t[103]) | (t[97] & ~t[98] & t[99] & t[100] & ~t[103]) | (t[97] & ~t[98] & t[101] & t[102] & ~t[103]) | (t[98] & ~t[100] & ~t[102] & t[103]) | (~t[98] & t[100] & t[102] & t[103]);
  assign t[72] = (t[97] & t[98] & t[99] & ~t[100] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & ~t[100] & ~t[101] & t[102] & t[103]) | (~t[98] & ~t[99] & t[100] & ~t[101] & ~t[102]) | (~t[97] & ~t[99] & t[100] & ~t[102] & ~t[103]) | (~t[97] & ~t[98] & t[100] & ~t[101] & ~t[103]) | (~t[98] & t[99] & t[100] & t[101] & ~t[102]) | (~t[99] & t[100] & t[101] & ~t[103]);
  assign t[73] = (t[97] & t[98] & ~t[99] & ~t[101] & t[102] & ~t[103]) | (t[97] & t[99] & ~t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & t[101] & ~t[102] & ~t[103]) | (~t[97] & ~t[99] & ~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[98] & ~t[100] & t[101] & ~t[103]) | (~t[97] & ~t[99] & t[100] & t[101] & t[102]) | (t[100] & t[101] & ~t[102] & ~t[103]);
  assign t[74] = (t[97] & t[98] & ~t[100] & t[101] & ~t[102] & ~t[103]) | (t[98] & ~t[99] & t[100] & ~t[101] & ~t[102] & t[103]) | (~t[98] & ~t[99] & ~t[100] & ~t[101] & t[102]) | (~t[97] & ~t[100] & ~t[101] & t[102] & ~t[103]) | (~t[97] & ~t[98] & ~t[99] & t[102] & ~t[103]) | (~t[98] & t[99] & ~t[100] & t[101] & t[102]) | (t[99] & ~t[101] & t[102] & ~t[103]);
  assign t[75] = (t[83] & t[84] & ~t[85] & t[86] & ~t[87] & ~t[89]) | (t[83] & ~t[85] & ~t[86] & t[87] & ~t[88] & t[89]) | (~t[84] & t[85] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[84] & t[85] & ~t[88] & ~t[89]) | (~t[83] & t[85] & t[86] & ~t[87] & t[88]) | (t[85] & ~t[86] & t[88] & ~t[89]);
  assign t[76] = (t[104] & ~t[106] & ~t[107] & ~t[108] & ~t[109]) | (t[104] & ~t[105] & ~t[107] & ~t[108] & ~t[110]) | (t[104] & ~t[105] & ~t[106] & ~t[109] & ~t[110]) | (~t[104] & t[105] & t[106] & t[107] & ~t[110]) | (~t[104] & t[105] & t[108] & t[109] & ~t[110]) | (t[104] & ~t[106] & ~t[108] & t[110]) | (~t[104] & t[106] & t[108] & t[110]);
  assign t[77] = (t[104] & t[105] & ~t[106] & ~t[108] & t[109] & ~t[110]) | (t[104] & t[106] & ~t[107] & ~t[108] & ~t[109] & t[110]) | (~t[105] & ~t[106] & t[108] & ~t[109] & ~t[110]) | (~t[104] & ~t[106] & ~t[107] & t[108] & ~t[109]) | (~t[104] & ~t[105] & ~t[107] & t[108] & ~t[110]) | (~t[104] & ~t[106] & t[107] & t[108] & t[109]) | (t[107] & t[108] & ~t[109] & ~t[110]);
  assign t[78] = (t[84] & ~t[85] & ~t[86] & ~t[87] & ~t[88]) | (~t[83] & t[84] & ~t[86] & ~t[87] & ~t[89]) | (~t[83] & t[84] & ~t[85] & ~t[88] & ~t[89]) | (t[83] & ~t[84] & t[85] & t[86] & ~t[89]) | (t[83] & ~t[84] & t[87] & t[88] & ~t[89]) | (t[84] & ~t[86] & ~t[88] & t[89]) | (~t[84] & t[86] & t[88] & t[89]);
  assign t[79] = (t[83] & t[84] & t[85] & ~t[86] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & ~t[86] & ~t[87] & t[88] & t[89]) | (~t[84] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (~t[83] & ~t[85] & t[86] & ~t[88] & ~t[89]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[89]) | (~t[84] & t[85] & t[86] & t[87] & ~t[88]) | (~t[85] & t[86] & t[87] & ~t[89]);
  assign t[7] = t[10] & t[11];
  assign t[80] = (t[83] & t[84] & ~t[86] & t[87] & ~t[88] & ~t[89]) | (t[84] & ~t[85] & t[86] & ~t[87] & ~t[88] & t[89]) | (~t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[86] & ~t[87] & t[88] & ~t[89]) | (~t[83] & ~t[84] & ~t[85] & t[88] & ~t[89]) | (~t[84] & t[85] & ~t[86] & t[87] & t[88]) | (t[85] & ~t[87] & t[88] & ~t[89]);
  assign t[81] = (t[111] & ~t[113] & ~t[114] & ~t[115] & ~t[116]) | (t[111] & ~t[112] & ~t[114] & ~t[115] & ~t[117]) | (t[111] & ~t[112] & ~t[113] & ~t[116] & ~t[117]) | (~t[111] & t[112] & t[113] & t[114] & ~t[117]) | (~t[111] & t[112] & t[115] & t[116] & ~t[117]) | (t[111] & ~t[113] & ~t[115] & t[117]) | (~t[111] & t[113] & t[115] & t[117]);
  assign t[82] = (t[111] & t[112] & ~t[113] & ~t[115] & t[116] & ~t[117]) | (t[111] & t[113] & ~t[114] & ~t[115] & ~t[116] & t[117]) | (~t[112] & ~t[113] & t[115] & ~t[116] & ~t[117]) | (~t[111] & ~t[113] & ~t[114] & t[115] & ~t[116]) | (~t[111] & ~t[112] & ~t[114] & t[115] & ~t[117]) | (~t[111] & ~t[113] & t[114] & t[115] & t[116]) | (t[114] & t[115] & ~t[116] & ~t[117]);
  assign t[83] = t[118] ^ x[7];
  assign t[84] = t[119] ^ x[39];
  assign t[85] = t[120] ^ x[29];
  assign t[86] = t[121] ^ x[40];
  assign t[87] = t[122] ^ x[8];
  assign t[88] = t[123] ^ x[41];
  assign t[89] = t[124] ^ x[6];
  assign t[8] = t[39] & t[12];
  assign t[90] = t[125] ^ x[15];
  assign t[91] = t[126] ^ x[10];
  assign t[92] = t[127] ^ x[11];
  assign t[93] = t[128] ^ x[12];
  assign t[94] = t[129] ^ x[16];
  assign t[95] = t[130] ^ x[13];
  assign t[96] = t[131] ^ x[14];
  assign t[97] = t[132] ^ x[22];
  assign t[98] = t[133] ^ x[24];
  assign t[99] = t[134] ^ x[23];
  assign t[9] = t[13] & t[14];
  assign y = (t[0] & ~t[21] & ~t[31]) | (~t[0] & t[21] & ~t[31]) | (~t[0] & ~t[21] & t[31]) | (t[0] & t[21] & t[31]);
endmodule

module R2ind135(x, y);
 input [40:0] x;
 output y;

 wire [121:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[101] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[102] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[103] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[104] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[105] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[106] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[107] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[108] = (x[18] & ~x[19] & ~x[20]) | (~x[18] & x[19] & ~x[20]) | (~x[18] & ~x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[109] = (x[18] & ~x[19] & ~x[21]) | (~x[18] & x[19] & ~x[21]) | (~x[18] & ~x[19] & x[21]) | (x[18] & x[19] & x[21]);
  assign t[10] = t[15] ^ t[13];
  assign t[110] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[111] = (x[18] & ~x[21]) | (~x[18] & x[21]);
  assign t[112] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[113] = (x[19] & ~x[21]) | (~x[19] & x[21]);
  assign t[114] = (x[20] & ~x[21]) | (~x[20] & x[21]);
  assign t[115] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[116] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[117] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[118] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[119] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = t[16] ^ t[9];
  assign t[120] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[121] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[31]);
  assign t[14] = ~(t[30] ^ t[13]);
  assign t[15] = t[32] ^ t[31];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[30] ^ t[20];
  assign t[1] = ~(t[2] ^ t[28]);
  assign t[20] = t[31] ^ t[33];
  assign t[21] = x[0] ? x[29] : t[22];
  assign t[22] = ~(t[23] ^ t[34]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[35]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[27]);
  assign t[27] = t[20] ^ t[9];
  assign t[28] = (t[36] & ~t[37]) | (~t[36] & t[37]);
  assign t[29] = (t[38] & ~t[39]) | (~t[38] & t[39]);
  assign t[2] = ~t[3];
  assign t[30] = (t[40] & ~t[41]) | (~t[40] & t[41]);
  assign t[31] = (t[40] & ~t[43] & ~t[45]) | (~t[42] & t[43] & ~t[44]) | (~t[40] & ~t[43] & t[45]) | (t[42] & t[43] & t[44]);
  assign t[32] = (t[40] & ~t[44]) | (~t[40] & t[44]);
  assign t[33] = (t[40] & ~t[43] & ~t[44]) | (~t[42] & t[43] & ~t[45]) | (~t[40] & ~t[43] & t[44]) | (t[42] & t[43] & t[45]);
  assign t[34] = (t[36] & ~t[47] & ~t[48]) | (~t[46] & t[47] & ~t[37]) | (~t[36] & ~t[47] & t[48]) | (t[46] & t[47] & t[37]);
  assign t[35] = (t[49] & ~t[50]) | (~t[49] & t[50]);
  assign t[36] = t[51] ^ x[8];
  assign t[37] = t[52] ^ x[9];
  assign t[38] = t[53] ^ x[16];
  assign t[39] = t[54] ^ x[17];
  assign t[3] = ~(t[4] ^ t[29]);
  assign t[40] = t[55] ^ x[23];
  assign t[41] = t[56] ^ x[24];
  assign t[42] = t[57] ^ x[25];
  assign t[43] = t[58] ^ x[26];
  assign t[44] = t[59] ^ x[27];
  assign t[45] = t[60] ^ x[28];
  assign t[46] = t[61] ^ x[30];
  assign t[47] = t[62] ^ x[31];
  assign t[48] = t[63] ^ x[32];
  assign t[49] = t[64] ^ x[39];
  assign t[4] = ~t[5];
  assign t[50] = t[65] ^ x[40];
  assign t[51] = (t[66] & ~t[68] & ~t[69] & ~t[70] & ~t[71]) | (t[66] & ~t[67] & ~t[69] & ~t[70] & ~t[72]) | (t[66] & ~t[67] & ~t[68] & ~t[71] & ~t[72]) | (~t[66] & t[67] & t[68] & t[69] & ~t[72]) | (~t[66] & t[67] & t[70] & t[71] & ~t[72]) | (t[66] & ~t[68] & ~t[70] & t[72]) | (~t[66] & t[68] & t[70] & t[72]);
  assign t[52] = (t[66] & t[67] & ~t[68] & ~t[70] & t[71] & ~t[72]) | (t[66] & t[68] & ~t[69] & ~t[70] & ~t[71] & t[72]) | (~t[67] & ~t[68] & t[70] & ~t[71] & ~t[72]) | (~t[66] & ~t[68] & ~t[69] & t[70] & ~t[71]) | (~t[66] & ~t[67] & ~t[69] & t[70] & ~t[72]) | (~t[66] & ~t[68] & t[69] & t[70] & t[71]) | (t[69] & t[70] & ~t[71] & ~t[72]);
  assign t[53] = (t[73] & ~t[75] & ~t[76] & ~t[77] & ~t[78]) | (t[73] & ~t[74] & ~t[76] & ~t[77] & ~t[79]) | (t[73] & ~t[74] & ~t[75] & ~t[78] & ~t[79]) | (~t[73] & t[74] & t[75] & t[76] & ~t[79]) | (~t[73] & t[74] & t[77] & t[78] & ~t[79]) | (t[73] & ~t[75] & ~t[77] & t[79]) | (~t[73] & t[75] & t[77] & t[79]);
  assign t[54] = (t[73] & t[74] & ~t[75] & ~t[77] & t[78] & ~t[79]) | (t[73] & t[75] & ~t[76] & ~t[77] & ~t[78] & t[79]) | (~t[74] & ~t[75] & t[77] & ~t[78] & ~t[79]) | (~t[73] & ~t[75] & ~t[76] & t[77] & ~t[78]) | (~t[73] & ~t[74] & ~t[76] & t[77] & ~t[79]) | (~t[73] & ~t[75] & t[76] & t[77] & t[78]) | (t[76] & t[77] & ~t[78] & ~t[79]);
  assign t[55] = (t[80] & ~t[82] & ~t[83] & ~t[84] & ~t[85]) | (t[80] & ~t[81] & ~t[83] & ~t[84] & ~t[86]) | (t[80] & ~t[81] & ~t[82] & ~t[85] & ~t[86]) | (~t[80] & t[81] & t[82] & t[83] & ~t[86]) | (~t[80] & t[81] & t[84] & t[85] & ~t[86]) | (t[80] & ~t[82] & ~t[84] & t[86]) | (~t[80] & t[82] & t[84] & t[86]);
  assign t[56] = (t[80] & t[81] & ~t[82] & t[83] & ~t[84] & ~t[86]) | (t[80] & ~t[82] & ~t[83] & t[84] & ~t[85] & t[86]) | (~t[81] & t[82] & ~t[83] & ~t[84] & ~t[86]) | (~t[80] & t[82] & ~t[83] & ~t[84] & ~t[85]) | (~t[80] & ~t[81] & t[82] & ~t[85] & ~t[86]) | (~t[80] & t[82] & t[83] & ~t[84] & t[85]) | (t[82] & ~t[83] & t[85] & ~t[86]);
  assign t[57] = (t[81] & ~t[82] & ~t[83] & ~t[84] & ~t[85]) | (~t[80] & t[81] & ~t[83] & ~t[84] & ~t[86]) | (~t[80] & t[81] & ~t[82] & ~t[85] & ~t[86]) | (t[80] & ~t[81] & t[82] & t[83] & ~t[86]) | (t[80] & ~t[81] & t[84] & t[85] & ~t[86]) | (t[81] & ~t[83] & ~t[85] & t[86]) | (~t[81] & t[83] & t[85] & t[86]);
  assign t[58] = (t[80] & t[81] & t[82] & ~t[83] & ~t[85] & ~t[86]) | (t[81] & ~t[82] & ~t[83] & ~t[84] & t[85] & t[86]) | (~t[81] & ~t[82] & t[83] & ~t[84] & ~t[85]) | (~t[80] & ~t[82] & t[83] & ~t[85] & ~t[86]) | (~t[80] & ~t[81] & t[83] & ~t[84] & ~t[86]) | (~t[81] & t[82] & t[83] & t[84] & ~t[85]) | (~t[82] & t[83] & t[84] & ~t[86]);
  assign t[59] = (t[80] & t[81] & ~t[82] & ~t[84] & t[85] & ~t[86]) | (t[80] & t[82] & ~t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[82] & t[84] & ~t[85] & ~t[86]) | (~t[80] & ~t[82] & ~t[83] & t[84] & ~t[85]) | (~t[80] & ~t[81] & ~t[83] & t[84] & ~t[86]) | (~t[80] & ~t[82] & t[83] & t[84] & t[85]) | (t[83] & t[84] & ~t[85] & ~t[86]);
  assign t[5] = t[6] ^ t[7];
  assign t[60] = (t[80] & t[81] & ~t[83] & t[84] & ~t[85] & ~t[86]) | (t[81] & ~t[82] & t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[82] & ~t[83] & ~t[84] & t[85]) | (~t[80] & ~t[83] & ~t[84] & t[85] & ~t[86]) | (~t[80] & ~t[81] & ~t[82] & t[85] & ~t[86]) | (~t[81] & t[82] & ~t[83] & t[84] & t[85]) | (t[82] & ~t[84] & t[85] & ~t[86]);
  assign t[61] = (t[67] & ~t[68] & ~t[69] & ~t[70] & ~t[71]) | (~t[66] & t[67] & ~t[69] & ~t[70] & ~t[72]) | (~t[66] & t[67] & ~t[68] & ~t[71] & ~t[72]) | (t[66] & ~t[67] & t[68] & t[69] & ~t[72]) | (t[66] & ~t[67] & t[70] & t[71] & ~t[72]) | (t[67] & ~t[69] & ~t[71] & t[72]) | (~t[67] & t[69] & t[71] & t[72]);
  assign t[62] = (t[66] & t[67] & t[68] & ~t[69] & ~t[71] & ~t[72]) | (t[67] & ~t[68] & ~t[69] & ~t[70] & t[71] & t[72]) | (~t[67] & ~t[68] & t[69] & ~t[70] & ~t[71]) | (~t[66] & ~t[68] & t[69] & ~t[71] & ~t[72]) | (~t[66] & ~t[67] & t[69] & ~t[70] & ~t[72]) | (~t[67] & t[68] & t[69] & t[70] & ~t[71]) | (~t[68] & t[69] & t[70] & ~t[72]);
  assign t[63] = (t[66] & t[67] & ~t[69] & t[70] & ~t[71] & ~t[72]) | (t[67] & ~t[68] & t[69] & ~t[70] & ~t[71] & t[72]) | (~t[67] & ~t[68] & ~t[69] & ~t[70] & t[71]) | (~t[66] & ~t[69] & ~t[70] & t[71] & ~t[72]) | (~t[66] & ~t[67] & ~t[68] & t[71] & ~t[72]) | (~t[67] & t[68] & ~t[69] & t[70] & t[71]) | (t[68] & ~t[70] & t[71] & ~t[72]);
  assign t[64] = (t[87] & ~t[89] & ~t[90] & ~t[91] & ~t[92]) | (t[87] & ~t[88] & ~t[90] & ~t[91] & ~t[93]) | (t[87] & ~t[88] & ~t[89] & ~t[92] & ~t[93]) | (~t[87] & t[88] & t[89] & t[90] & ~t[93]) | (~t[87] & t[88] & t[91] & t[92] & ~t[93]) | (t[87] & ~t[89] & ~t[91] & t[93]) | (~t[87] & t[89] & t[91] & t[93]);
  assign t[65] = (t[87] & t[88] & ~t[89] & ~t[91] & t[92] & ~t[93]) | (t[87] & t[89] & ~t[90] & ~t[91] & ~t[92] & t[93]) | (~t[88] & ~t[89] & t[91] & ~t[92] & ~t[93]) | (~t[87] & ~t[89] & ~t[90] & t[91] & ~t[92]) | (~t[87] & ~t[88] & ~t[90] & t[91] & ~t[93]) | (~t[87] & ~t[89] & t[90] & t[91] & t[92]) | (t[90] & t[91] & ~t[92] & ~t[93]);
  assign t[66] = t[94] ^ x[8];
  assign t[67] = t[95] ^ x[30];
  assign t[68] = t[96] ^ x[6];
  assign t[69] = t[97] ^ x[31];
  assign t[6] = t[8] ^ t[9];
  assign t[70] = t[98] ^ x[9];
  assign t[71] = t[99] ^ x[32];
  assign t[72] = t[100] ^ x[7];
  assign t[73] = t[101] ^ x[16];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[12];
  assign t[76] = t[104] ^ x[13];
  assign t[77] = t[105] ^ x[17];
  assign t[78] = t[106] ^ x[14];
  assign t[79] = t[107] ^ x[15];
  assign t[7] = t[10] & t[11];
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[24];
  assign t[83] = t[111] ^ x[26];
  assign t[84] = t[112] ^ x[27];
  assign t[85] = t[113] ^ x[28];
  assign t[86] = t[114] ^ x[22];
  assign t[87] = t[115] ^ x[39];
  assign t[88] = t[116] ^ x[34];
  assign t[89] = t[117] ^ x[35];
  assign t[8] = t[30] & t[12];
  assign t[90] = t[118] ^ x[36];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = t[120] ^ x[37];
  assign t[93] = t[121] ^ x[38];
  assign t[94] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[95] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[96] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[97] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[98] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[99] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[9] = t[13] & t[14];
  assign y = (t[0] & ~t[21]) | (~t[0] & t[21]);
endmodule

module R2ind136(x, y);
 input [40:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[101] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[102] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[103] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[104] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[105] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[106] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[107] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (x[18] & ~x[19] & ~x[20]) | (~x[18] & x[19] & ~x[20]) | (~x[18] & ~x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[10] = t[15] ^ t[13];
  assign t[110] = (x[18] & ~x[19] & ~x[21]) | (~x[18] & x[19] & ~x[21]) | (~x[18] & ~x[19] & x[21]) | (x[18] & x[19] & x[21]);
  assign t[111] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[112] = (x[18] & ~x[21]) | (~x[18] & x[21]);
  assign t[113] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[114] = (x[19] & ~x[21]) | (~x[19] & x[21]);
  assign t[115] = (x[20] & ~x[21]) | (~x[20] & x[21]);
  assign t[116] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[117] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[118] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[119] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[11] = t[16] ^ t[9];
  assign t[120] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[121] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = t[17] ^ t[18];
  assign t[13] = ~(t[32]);
  assign t[14] = ~(t[31] ^ t[13]);
  assign t[15] = t[33] ^ t[32];
  assign t[16] = ~(t[19] ^ t[10]);
  assign t[17] = t[31] ^ t[15];
  assign t[18] = t[13] & t[19];
  assign t[19] = t[31] ^ t[20];
  assign t[1] = ~(t[2] ^ t[29]);
  assign t[20] = t[32] ^ t[34];
  assign t[21] = x[0] ? x[29] : t[22];
  assign t[22] = ~(t[23] ^ t[35]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[36]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[27]);
  assign t[27] = t[28] ^ t[9];
  assign t[28] = t[15] ^ t[18];
  assign t[29] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[2] = ~t[3];
  assign t[30] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[31] = (t[41] & ~t[42]) | (~t[41] & t[42]);
  assign t[32] = (t[41] & ~t[44] & ~t[46]) | (~t[43] & t[44] & ~t[45]) | (~t[41] & ~t[44] & t[46]) | (t[43] & t[44] & t[45]);
  assign t[33] = (t[41] & ~t[45]) | (~t[41] & t[45]);
  assign t[34] = (t[41] & ~t[44] & ~t[45]) | (~t[43] & t[44] & ~t[46]) | (~t[41] & ~t[44] & t[45]) | (t[43] & t[44] & t[46]);
  assign t[35] = (t[37] & ~t[48] & ~t[38]) | (~t[47] & t[48] & ~t[49]) | (~t[37] & ~t[48] & t[38]) | (t[47] & t[48] & t[49]);
  assign t[36] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[37] = t[52] ^ x[8];
  assign t[38] = t[53] ^ x[9];
  assign t[39] = t[54] ^ x[16];
  assign t[3] = ~(t[4] ^ t[30]);
  assign t[40] = t[55] ^ x[17];
  assign t[41] = t[56] ^ x[23];
  assign t[42] = t[57] ^ x[24];
  assign t[43] = t[58] ^ x[25];
  assign t[44] = t[59] ^ x[26];
  assign t[45] = t[60] ^ x[27];
  assign t[46] = t[61] ^ x[28];
  assign t[47] = t[62] ^ x[30];
  assign t[48] = t[63] ^ x[31];
  assign t[49] = t[64] ^ x[32];
  assign t[4] = ~t[5];
  assign t[50] = t[65] ^ x[39];
  assign t[51] = t[66] ^ x[40];
  assign t[52] = (t[67] & ~t[69] & ~t[70] & ~t[71] & ~t[72]) | (t[67] & ~t[68] & ~t[70] & ~t[71] & ~t[73]) | (t[67] & ~t[68] & ~t[69] & ~t[72] & ~t[73]) | (~t[67] & t[68] & t[69] & t[70] & ~t[73]) | (~t[67] & t[68] & t[71] & t[72] & ~t[73]) | (t[67] & ~t[69] & ~t[71] & t[73]) | (~t[67] & t[69] & t[71] & t[73]);
  assign t[53] = (t[67] & t[68] & ~t[69] & ~t[71] & t[72] & ~t[73]) | (t[67] & t[69] & ~t[70] & ~t[71] & ~t[72] & t[73]) | (~t[68] & ~t[69] & t[71] & ~t[72] & ~t[73]) | (~t[67] & ~t[69] & ~t[70] & t[71] & ~t[72]) | (~t[67] & ~t[68] & ~t[70] & t[71] & ~t[73]) | (~t[67] & ~t[69] & t[70] & t[71] & t[72]) | (t[70] & t[71] & ~t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[76] & ~t[77] & ~t[78] & ~t[79]) | (t[74] & ~t[75] & ~t[77] & ~t[78] & ~t[80]) | (t[74] & ~t[75] & ~t[76] & ~t[79] & ~t[80]) | (~t[74] & t[75] & t[76] & t[77] & ~t[80]) | (~t[74] & t[75] & t[78] & t[79] & ~t[80]) | (t[74] & ~t[76] & ~t[78] & t[80]) | (~t[74] & t[76] & t[78] & t[80]);
  assign t[55] = (t[74] & t[75] & ~t[76] & ~t[78] & t[79] & ~t[80]) | (t[74] & t[76] & ~t[77] & ~t[78] & ~t[79] & t[80]) | (~t[75] & ~t[76] & t[78] & ~t[79] & ~t[80]) | (~t[74] & ~t[76] & ~t[77] & t[78] & ~t[79]) | (~t[74] & ~t[75] & ~t[77] & t[78] & ~t[80]) | (~t[74] & ~t[76] & t[77] & t[78] & t[79]) | (t[77] & t[78] & ~t[79] & ~t[80]);
  assign t[56] = (t[81] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (t[81] & ~t[82] & ~t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[82] & ~t[83] & ~t[86] & ~t[87]) | (~t[81] & t[82] & t[83] & t[84] & ~t[87]) | (~t[81] & t[82] & t[85] & t[86] & ~t[87]) | (t[81] & ~t[83] & ~t[85] & t[87]) | (~t[81] & t[83] & t[85] & t[87]);
  assign t[57] = (t[81] & t[82] & ~t[83] & t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[83] & ~t[84] & t[85] & ~t[86] & t[87]) | (~t[82] & t[83] & ~t[84] & ~t[85] & ~t[87]) | (~t[81] & t[83] & ~t[84] & ~t[85] & ~t[86]) | (~t[81] & ~t[82] & t[83] & ~t[86] & ~t[87]) | (~t[81] & t[83] & t[84] & ~t[85] & t[86]) | (t[83] & ~t[84] & t[86] & ~t[87]);
  assign t[58] = (t[82] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (~t[81] & t[82] & ~t[84] & ~t[85] & ~t[87]) | (~t[81] & t[82] & ~t[83] & ~t[86] & ~t[87]) | (t[81] & ~t[82] & t[83] & t[84] & ~t[87]) | (t[81] & ~t[82] & t[85] & t[86] & ~t[87]) | (t[82] & ~t[84] & ~t[86] & t[87]) | (~t[82] & t[84] & t[86] & t[87]);
  assign t[59] = (t[81] & t[82] & t[83] & ~t[84] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & ~t[84] & ~t[85] & t[86] & t[87]) | (~t[82] & ~t[83] & t[84] & ~t[85] & ~t[86]) | (~t[81] & ~t[83] & t[84] & ~t[86] & ~t[87]) | (~t[81] & ~t[82] & t[84] & ~t[85] & ~t[87]) | (~t[82] & t[83] & t[84] & t[85] & ~t[86]) | (~t[83] & t[84] & t[85] & ~t[87]);
  assign t[5] = t[6] ^ t[7];
  assign t[60] = (t[81] & t[82] & ~t[83] & ~t[85] & t[86] & ~t[87]) | (t[81] & t[83] & ~t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & t[85] & ~t[86] & ~t[87]) | (~t[81] & ~t[83] & ~t[84] & t[85] & ~t[86]) | (~t[81] & ~t[82] & ~t[84] & t[85] & ~t[87]) | (~t[81] & ~t[83] & t[84] & t[85] & t[86]) | (t[84] & t[85] & ~t[86] & ~t[87]);
  assign t[61] = (t[81] & t[82] & ~t[84] & t[85] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[84] & ~t[85] & t[86] & ~t[87]) | (~t[81] & ~t[82] & ~t[83] & t[86] & ~t[87]) | (~t[82] & t[83] & ~t[84] & t[85] & t[86]) | (t[83] & ~t[85] & t[86] & ~t[87]);
  assign t[62] = (t[68] & ~t[69] & ~t[70] & ~t[71] & ~t[72]) | (~t[67] & t[68] & ~t[70] & ~t[71] & ~t[73]) | (~t[67] & t[68] & ~t[69] & ~t[72] & ~t[73]) | (t[67] & ~t[68] & t[69] & t[70] & ~t[73]) | (t[67] & ~t[68] & t[71] & t[72] & ~t[73]) | (t[68] & ~t[70] & ~t[72] & t[73]) | (~t[68] & t[70] & t[72] & t[73]);
  assign t[63] = (t[67] & t[68] & t[69] & ~t[70] & ~t[72] & ~t[73]) | (t[68] & ~t[69] & ~t[70] & ~t[71] & t[72] & t[73]) | (~t[68] & ~t[69] & t[70] & ~t[71] & ~t[72]) | (~t[67] & ~t[69] & t[70] & ~t[72] & ~t[73]) | (~t[67] & ~t[68] & t[70] & ~t[71] & ~t[73]) | (~t[68] & t[69] & t[70] & t[71] & ~t[72]) | (~t[69] & t[70] & t[71] & ~t[73]);
  assign t[64] = (t[67] & t[68] & ~t[70] & t[71] & ~t[72] & ~t[73]) | (t[68] & ~t[69] & t[70] & ~t[71] & ~t[72] & t[73]) | (~t[68] & ~t[69] & ~t[70] & ~t[71] & t[72]) | (~t[67] & ~t[70] & ~t[71] & t[72] & ~t[73]) | (~t[67] & ~t[68] & ~t[69] & t[72] & ~t[73]) | (~t[68] & t[69] & ~t[70] & t[71] & t[72]) | (t[69] & ~t[71] & t[72] & ~t[73]);
  assign t[65] = (t[88] & ~t[90] & ~t[91] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & ~t[91] & ~t[92] & ~t[94]) | (t[88] & ~t[89] & ~t[90] & ~t[93] & ~t[94]) | (~t[88] & t[89] & t[90] & t[91] & ~t[94]) | (~t[88] & t[89] & t[92] & t[93] & ~t[94]) | (t[88] & ~t[90] & ~t[92] & t[94]) | (~t[88] & t[90] & t[92] & t[94]);
  assign t[66] = (t[88] & t[89] & ~t[90] & ~t[92] & t[93] & ~t[94]) | (t[88] & t[90] & ~t[91] & ~t[92] & ~t[93] & t[94]) | (~t[89] & ~t[90] & t[92] & ~t[93] & ~t[94]) | (~t[88] & ~t[90] & ~t[91] & t[92] & ~t[93]) | (~t[88] & ~t[89] & ~t[91] & t[92] & ~t[94]) | (~t[88] & ~t[90] & t[91] & t[92] & t[93]) | (t[91] & t[92] & ~t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[8];
  assign t[68] = t[96] ^ x[30];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = t[8] ^ t[9];
  assign t[70] = t[98] ^ x[31];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[32];
  assign t[73] = t[101] ^ x[7];
  assign t[74] = t[102] ^ x[16];
  assign t[75] = t[103] ^ x[11];
  assign t[76] = t[104] ^ x[12];
  assign t[77] = t[105] ^ x[13];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[14];
  assign t[7] = t[10] & t[11];
  assign t[80] = t[108] ^ x[15];
  assign t[81] = t[109] ^ x[23];
  assign t[82] = t[110] ^ x[25];
  assign t[83] = t[111] ^ x[24];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[27];
  assign t[86] = t[114] ^ x[28];
  assign t[87] = t[115] ^ x[22];
  assign t[88] = t[116] ^ x[39];
  assign t[89] = t[117] ^ x[34];
  assign t[8] = t[31] & t[12];
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[36];
  assign t[92] = t[120] ^ x[40];
  assign t[93] = t[121] ^ x[37];
  assign t[94] = t[122] ^ x[38];
  assign t[95] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[96] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[97] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[98] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[99] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[9] = t[13] & t[14];
  assign y = (t[0] & ~t[21]) | (~t[0] & t[21]);
endmodule

module R2ind137(x, y);
 input [40:0] x;
 output y;

 wire [123:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[101] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[102] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[103] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[104] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[105] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[106] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[107] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[10] = t[16] ^ t[9];
  assign t[110] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[111] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[112] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[113] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[114] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[115] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[116] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[117] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[118] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[119] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[11] = t[30] ^ t[14];
  assign t[120] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[121] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[123] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = t[31] ^ t[32];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[32]);
  assign t[15] = ~(t[30] ^ t[14]);
  assign t[16] = t[30] & t[18];
  assign t[17] = t[30] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[28]);
  assign t[20] = t[30] ^ t[12];
  assign t[21] = x[0] ? x[28] : t[22];
  assign t[22] = ~(t[23] ^ t[34]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[35]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[27]);
  assign t[27] = t[19] ^ t[9];
  assign t[28] = (t[36] & ~t[37]) | (~t[36] & t[37]);
  assign t[29] = (t[38] & ~t[39]) | (~t[38] & t[39]);
  assign t[2] = ~t[3];
  assign t[30] = (t[40] & ~t[41]) | (~t[40] & t[41]);
  assign t[31] = (t[40] & ~t[42]) | (~t[40] & t[42]);
  assign t[32] = (t[40] & ~t[44] & ~t[45]) | (~t[43] & t[44] & ~t[42]) | (~t[40] & ~t[44] & t[45]) | (t[43] & t[44] & t[42]);
  assign t[33] = (t[40] & ~t[44] & ~t[42]) | (~t[43] & t[44] & ~t[45]) | (~t[40] & ~t[44] & t[42]) | (t[43] & t[44] & t[45]);
  assign t[34] = (t[36] & ~t[47] & ~t[49]) | (~t[46] & t[47] & ~t[48]) | (~t[36] & ~t[47] & t[49]) | (t[46] & t[47] & t[48]);
  assign t[35] = (t[50] & ~t[51]) | (~t[50] & t[51]);
  assign t[36] = t[52] ^ x[7];
  assign t[37] = t[53] ^ x[8];
  assign t[38] = t[54] ^ x[15];
  assign t[39] = t[55] ^ x[16];
  assign t[3] = ~(t[4] ^ t[29]);
  assign t[40] = t[56] ^ x[22];
  assign t[41] = t[57] ^ x[23];
  assign t[42] = t[58] ^ x[24];
  assign t[43] = t[59] ^ x[25];
  assign t[44] = t[60] ^ x[26];
  assign t[45] = t[61] ^ x[27];
  assign t[46] = t[62] ^ x[29];
  assign t[47] = t[63] ^ x[30];
  assign t[48] = t[64] ^ x[31];
  assign t[49] = t[65] ^ x[32];
  assign t[4] = ~t[5];
  assign t[50] = t[66] ^ x[39];
  assign t[51] = t[67] ^ x[40];
  assign t[52] = (t[68] & ~t[70] & ~t[71] & ~t[72] & ~t[73]) | (t[68] & ~t[69] & ~t[71] & ~t[72] & ~t[74]) | (t[68] & ~t[69] & ~t[70] & ~t[73] & ~t[74]) | (~t[68] & t[69] & t[70] & t[71] & ~t[74]) | (~t[68] & t[69] & t[72] & t[73] & ~t[74]) | (t[68] & ~t[70] & ~t[72] & t[74]) | (~t[68] & t[70] & t[72] & t[74]);
  assign t[53] = (t[68] & t[69] & ~t[70] & t[71] & ~t[72] & ~t[74]) | (t[68] & ~t[70] & ~t[71] & t[72] & ~t[73] & t[74]) | (~t[69] & t[70] & ~t[71] & ~t[72] & ~t[74]) | (~t[68] & t[70] & ~t[71] & ~t[72] & ~t[73]) | (~t[68] & ~t[69] & t[70] & ~t[73] & ~t[74]) | (~t[68] & t[70] & t[71] & ~t[72] & t[73]) | (t[70] & ~t[71] & t[73] & ~t[74]);
  assign t[54] = (t[75] & ~t[77] & ~t[78] & ~t[79] & ~t[80]) | (t[75] & ~t[76] & ~t[78] & ~t[79] & ~t[81]) | (t[75] & ~t[76] & ~t[77] & ~t[80] & ~t[81]) | (~t[75] & t[76] & t[77] & t[78] & ~t[81]) | (~t[75] & t[76] & t[79] & t[80] & ~t[81]) | (t[75] & ~t[77] & ~t[79] & t[81]) | (~t[75] & t[77] & t[79] & t[81]);
  assign t[55] = (t[75] & t[76] & ~t[77] & ~t[79] & t[80] & ~t[81]) | (t[75] & t[77] & ~t[78] & ~t[79] & ~t[80] & t[81]) | (~t[76] & ~t[77] & t[79] & ~t[80] & ~t[81]) | (~t[75] & ~t[77] & ~t[78] & t[79] & ~t[80]) | (~t[75] & ~t[76] & ~t[78] & t[79] & ~t[81]) | (~t[75] & ~t[77] & t[78] & t[79] & t[80]) | (t[78] & t[79] & ~t[80] & ~t[81]);
  assign t[56] = (t[82] & ~t[84] & ~t[85] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & ~t[85] & ~t[86] & ~t[88]) | (t[82] & ~t[83] & ~t[84] & ~t[87] & ~t[88]) | (~t[82] & t[83] & t[84] & t[85] & ~t[88]) | (~t[82] & t[83] & t[86] & t[87] & ~t[88]) | (t[82] & ~t[84] & ~t[86] & t[88]) | (~t[82] & t[84] & t[86] & t[88]);
  assign t[57] = (t[82] & t[83] & ~t[84] & t[85] & ~t[86] & ~t[88]) | (t[82] & ~t[84] & ~t[85] & t[86] & ~t[87] & t[88]) | (~t[83] & t[84] & ~t[85] & ~t[86] & ~t[88]) | (~t[82] & t[84] & ~t[85] & ~t[86] & ~t[87]) | (~t[82] & ~t[83] & t[84] & ~t[87] & ~t[88]) | (~t[82] & t[84] & t[85] & ~t[86] & t[87]) | (t[84] & ~t[85] & t[87] & ~t[88]);
  assign t[58] = (t[82] & t[83] & ~t[84] & ~t[86] & t[87] & ~t[88]) | (t[82] & t[84] & ~t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[84] & t[86] & ~t[87] & ~t[88]) | (~t[82] & ~t[84] & ~t[85] & t[86] & ~t[87]) | (~t[82] & ~t[83] & ~t[85] & t[86] & ~t[88]) | (~t[82] & ~t[84] & t[85] & t[86] & t[87]) | (t[85] & t[86] & ~t[87] & ~t[88]);
  assign t[59] = (t[83] & ~t[84] & ~t[85] & ~t[86] & ~t[87]) | (~t[82] & t[83] & ~t[85] & ~t[86] & ~t[88]) | (~t[82] & t[83] & ~t[84] & ~t[87] & ~t[88]) | (t[82] & ~t[83] & t[84] & t[85] & ~t[88]) | (t[82] & ~t[83] & t[86] & t[87] & ~t[88]) | (t[83] & ~t[85] & ~t[87] & t[88]) | (~t[83] & t[85] & t[87] & t[88]);
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[60] = (t[82] & t[83] & t[84] & ~t[85] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & ~t[85] & ~t[86] & t[87] & t[88]) | (~t[83] & ~t[84] & t[85] & ~t[86] & ~t[87]) | (~t[82] & ~t[84] & t[85] & ~t[87] & ~t[88]) | (~t[82] & ~t[83] & t[85] & ~t[86] & ~t[88]) | (~t[83] & t[84] & t[85] & t[86] & ~t[87]) | (~t[84] & t[85] & t[86] & ~t[88]);
  assign t[61] = (t[82] & t[83] & ~t[85] & t[86] & ~t[87] & ~t[88]) | (t[83] & ~t[84] & t[85] & ~t[86] & ~t[87] & t[88]) | (~t[83] & ~t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[85] & ~t[86] & t[87] & ~t[88]) | (~t[82] & ~t[83] & ~t[84] & t[87] & ~t[88]) | (~t[83] & t[84] & ~t[85] & t[86] & t[87]) | (t[84] & ~t[86] & t[87] & ~t[88]);
  assign t[62] = (t[69] & ~t[70] & ~t[71] & ~t[72] & ~t[73]) | (~t[68] & t[69] & ~t[71] & ~t[72] & ~t[74]) | (~t[68] & t[69] & ~t[70] & ~t[73] & ~t[74]) | (t[68] & ~t[69] & t[70] & t[71] & ~t[74]) | (t[68] & ~t[69] & t[72] & t[73] & ~t[74]) | (t[69] & ~t[71] & ~t[73] & t[74]) | (~t[69] & t[71] & t[73] & t[74]);
  assign t[63] = (t[68] & t[69] & t[70] & ~t[71] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & ~t[71] & ~t[72] & t[73] & t[74]) | (~t[69] & ~t[70] & t[71] & ~t[72] & ~t[73]) | (~t[68] & ~t[70] & t[71] & ~t[73] & ~t[74]) | (~t[68] & ~t[69] & t[71] & ~t[72] & ~t[74]) | (~t[69] & t[70] & t[71] & t[72] & ~t[73]) | (~t[70] & t[71] & t[72] & ~t[74]);
  assign t[64] = (t[68] & t[69] & ~t[70] & ~t[72] & t[73] & ~t[74]) | (t[68] & t[70] & ~t[71] & ~t[72] & ~t[73] & t[74]) | (~t[69] & ~t[70] & t[72] & ~t[73] & ~t[74]) | (~t[68] & ~t[70] & ~t[71] & t[72] & ~t[73]) | (~t[68] & ~t[69] & ~t[71] & t[72] & ~t[74]) | (~t[68] & ~t[70] & t[71] & t[72] & t[73]) | (t[71] & t[72] & ~t[73] & ~t[74]);
  assign t[65] = (t[68] & t[69] & ~t[71] & t[72] & ~t[73] & ~t[74]) | (t[69] & ~t[70] & t[71] & ~t[72] & ~t[73] & t[74]) | (~t[69] & ~t[70] & ~t[71] & ~t[72] & t[73]) | (~t[68] & ~t[71] & ~t[72] & t[73] & ~t[74]) | (~t[68] & ~t[69] & ~t[70] & t[73] & ~t[74]) | (~t[69] & t[70] & ~t[71] & t[72] & t[73]) | (t[70] & ~t[72] & t[73] & ~t[74]);
  assign t[66] = (t[89] & ~t[91] & ~t[92] & ~t[93] & ~t[94]) | (t[89] & ~t[90] & ~t[92] & ~t[93] & ~t[95]) | (t[89] & ~t[90] & ~t[91] & ~t[94] & ~t[95]) | (~t[89] & t[90] & t[91] & t[92] & ~t[95]) | (~t[89] & t[90] & t[93] & t[94] & ~t[95]) | (t[89] & ~t[91] & ~t[93] & t[95]) | (~t[89] & t[91] & t[93] & t[95]);
  assign t[67] = (t[89] & t[90] & ~t[91] & ~t[93] & t[94] & ~t[95]) | (t[89] & t[91] & ~t[92] & ~t[93] & ~t[94] & t[95]) | (~t[90] & ~t[91] & t[93] & ~t[94] & ~t[95]) | (~t[89] & ~t[91] & ~t[92] & t[93] & ~t[94]) | (~t[89] & ~t[90] & ~t[92] & t[93] & ~t[95]) | (~t[89] & ~t[91] & t[92] & t[93] & t[94]) | (t[92] & t[93] & ~t[94] & ~t[95]);
  assign t[68] = t[96] ^ x[7];
  assign t[69] = t[97] ^ x[29];
  assign t[6] = t[8] ^ t[9];
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[30];
  assign t[72] = t[100] ^ x[31];
  assign t[73] = t[101] ^ x[32];
  assign t[74] = t[102] ^ x[6];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[10];
  assign t[77] = t[105] ^ x[11];
  assign t[78] = t[106] ^ x[12];
  assign t[79] = t[107] ^ x[16];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[108] ^ x[13];
  assign t[81] = t[109] ^ x[14];
  assign t[82] = t[110] ^ x[22];
  assign t[83] = t[111] ^ x[25];
  assign t[84] = t[112] ^ x[23];
  assign t[85] = t[113] ^ x[26];
  assign t[86] = t[114] ^ x[24];
  assign t[87] = t[115] ^ x[27];
  assign t[88] = t[116] ^ x[21];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[118] ^ x[34];
  assign t[91] = t[119] ^ x[35];
  assign t[92] = t[120] ^ x[36];
  assign t[93] = t[121] ^ x[40];
  assign t[94] = t[122] ^ x[37];
  assign t[95] = t[123] ^ x[38];
  assign t[96] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[97] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[98] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[99] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[21]) | (~t[0] & t[21]);
endmodule

module R2ind138(x, y);
 input [40:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[101] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[102] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[103] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[104] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[105] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[106] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[107] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[108] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[109] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[10] = t[16] ^ t[9];
  assign t[110] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[111] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[112] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[113] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[114] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[115] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[116] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[117] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[118] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[119] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[11] = t[29] ^ t[14];
  assign t[120] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[121] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[122] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[12] = t[30] ^ t[31];
  assign t[13] = t[14] & t[17];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[29] ^ t[14]);
  assign t[16] = t[29] & t[18];
  assign t[17] = t[29] ^ t[19];
  assign t[18] = t[20] ^ t[13];
  assign t[19] = t[31] ^ t[32];
  assign t[1] = ~(t[2] ^ t[27]);
  assign t[20] = t[29] ^ t[12];
  assign t[21] = x[0] ? x[28] : t[22];
  assign t[22] = ~(t[23] ^ t[33]);
  assign t[23] = ~t[24];
  assign t[24] = ~(t[25] ^ t[34]);
  assign t[25] = ~t[26];
  assign t[26] = ~(t[6]);
  assign t[27] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[28] = (t[37] & ~t[38]) | (~t[37] & t[38]);
  assign t[29] = (t[39] & ~t[40]) | (~t[39] & t[40]);
  assign t[2] = ~t[3];
  assign t[30] = (t[39] & ~t[41]) | (~t[39] & t[41]);
  assign t[31] = (t[39] & ~t[43] & ~t[44]) | (~t[42] & t[43] & ~t[41]) | (~t[39] & ~t[43] & t[44]) | (t[42] & t[43] & t[41]);
  assign t[32] = (t[39] & ~t[43] & ~t[41]) | (~t[42] & t[43] & ~t[44]) | (~t[39] & ~t[43] & t[41]) | (t[42] & t[43] & t[44]);
  assign t[33] = (t[35] & ~t[46] & ~t[47]) | (~t[45] & t[46] & ~t[48]) | (~t[35] & ~t[46] & t[47]) | (t[45] & t[46] & t[48]);
  assign t[34] = (t[49] & ~t[50]) | (~t[49] & t[50]);
  assign t[35] = t[51] ^ x[7];
  assign t[36] = t[52] ^ x[8];
  assign t[37] = t[53] ^ x[15];
  assign t[38] = t[54] ^ x[16];
  assign t[39] = t[55] ^ x[22];
  assign t[3] = ~(t[4] ^ t[28]);
  assign t[40] = t[56] ^ x[23];
  assign t[41] = t[57] ^ x[24];
  assign t[42] = t[58] ^ x[25];
  assign t[43] = t[59] ^ x[26];
  assign t[44] = t[60] ^ x[27];
  assign t[45] = t[61] ^ x[29];
  assign t[46] = t[62] ^ x[30];
  assign t[47] = t[63] ^ x[31];
  assign t[48] = t[64] ^ x[32];
  assign t[49] = t[65] ^ x[39];
  assign t[4] = ~t[5];
  assign t[50] = t[66] ^ x[40];
  assign t[51] = (t[67] & ~t[69] & ~t[70] & ~t[71] & ~t[72]) | (t[67] & ~t[68] & ~t[70] & ~t[71] & ~t[73]) | (t[67] & ~t[68] & ~t[69] & ~t[72] & ~t[73]) | (~t[67] & t[68] & t[69] & t[70] & ~t[73]) | (~t[67] & t[68] & t[71] & t[72] & ~t[73]) | (t[67] & ~t[69] & ~t[71] & t[73]) | (~t[67] & t[69] & t[71] & t[73]);
  assign t[52] = (t[67] & t[68] & ~t[69] & t[70] & ~t[71] & ~t[73]) | (t[67] & ~t[69] & ~t[70] & t[71] & ~t[72] & t[73]) | (~t[68] & t[69] & ~t[70] & ~t[71] & ~t[73]) | (~t[67] & t[69] & ~t[70] & ~t[71] & ~t[72]) | (~t[67] & ~t[68] & t[69] & ~t[72] & ~t[73]) | (~t[67] & t[69] & t[70] & ~t[71] & t[72]) | (t[69] & ~t[70] & t[72] & ~t[73]);
  assign t[53] = (t[74] & ~t[76] & ~t[77] & ~t[78] & ~t[79]) | (t[74] & ~t[75] & ~t[77] & ~t[78] & ~t[80]) | (t[74] & ~t[75] & ~t[76] & ~t[79] & ~t[80]) | (~t[74] & t[75] & t[76] & t[77] & ~t[80]) | (~t[74] & t[75] & t[78] & t[79] & ~t[80]) | (t[74] & ~t[76] & ~t[78] & t[80]) | (~t[74] & t[76] & t[78] & t[80]);
  assign t[54] = (t[74] & t[75] & ~t[76] & ~t[78] & t[79] & ~t[80]) | (t[74] & t[76] & ~t[77] & ~t[78] & ~t[79] & t[80]) | (~t[75] & ~t[76] & t[78] & ~t[79] & ~t[80]) | (~t[74] & ~t[76] & ~t[77] & t[78] & ~t[79]) | (~t[74] & ~t[75] & ~t[77] & t[78] & ~t[80]) | (~t[74] & ~t[76] & t[77] & t[78] & t[79]) | (t[77] & t[78] & ~t[79] & ~t[80]);
  assign t[55] = (t[81] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (t[81] & ~t[82] & ~t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[82] & ~t[83] & ~t[86] & ~t[87]) | (~t[81] & t[82] & t[83] & t[84] & ~t[87]) | (~t[81] & t[82] & t[85] & t[86] & ~t[87]) | (t[81] & ~t[83] & ~t[85] & t[87]) | (~t[81] & t[83] & t[85] & t[87]);
  assign t[56] = (t[81] & t[82] & ~t[83] & t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[83] & ~t[84] & t[85] & ~t[86] & t[87]) | (~t[82] & t[83] & ~t[84] & ~t[85] & ~t[87]) | (~t[81] & t[83] & ~t[84] & ~t[85] & ~t[86]) | (~t[81] & ~t[82] & t[83] & ~t[86] & ~t[87]) | (~t[81] & t[83] & t[84] & ~t[85] & t[86]) | (t[83] & ~t[84] & t[86] & ~t[87]);
  assign t[57] = (t[81] & t[82] & ~t[83] & ~t[85] & t[86] & ~t[87]) | (t[81] & t[83] & ~t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & t[85] & ~t[86] & ~t[87]) | (~t[81] & ~t[83] & ~t[84] & t[85] & ~t[86]) | (~t[81] & ~t[82] & ~t[84] & t[85] & ~t[87]) | (~t[81] & ~t[83] & t[84] & t[85] & t[86]) | (t[84] & t[85] & ~t[86] & ~t[87]);
  assign t[58] = (t[82] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (~t[81] & t[82] & ~t[84] & ~t[85] & ~t[87]) | (~t[81] & t[82] & ~t[83] & ~t[86] & ~t[87]) | (t[81] & ~t[82] & t[83] & t[84] & ~t[87]) | (t[81] & ~t[82] & t[85] & t[86] & ~t[87]) | (t[82] & ~t[84] & ~t[86] & t[87]) | (~t[82] & t[84] & t[86] & t[87]);
  assign t[59] = (t[81] & t[82] & t[83] & ~t[84] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & ~t[84] & ~t[85] & t[86] & t[87]) | (~t[82] & ~t[83] & t[84] & ~t[85] & ~t[86]) | (~t[81] & ~t[83] & t[84] & ~t[86] & ~t[87]) | (~t[81] & ~t[82] & t[84] & ~t[85] & ~t[87]) | (~t[82] & t[83] & t[84] & t[85] & ~t[86]) | (~t[83] & t[84] & t[85] & ~t[87]);
  assign t[5] = ~(t[6] ^ t[7]);
  assign t[60] = (t[81] & t[82] & ~t[84] & t[85] & ~t[86] & ~t[87]) | (t[82] & ~t[83] & t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & ~t[84] & ~t[85] & t[86]) | (~t[81] & ~t[84] & ~t[85] & t[86] & ~t[87]) | (~t[81] & ~t[82] & ~t[83] & t[86] & ~t[87]) | (~t[82] & t[83] & ~t[84] & t[85] & t[86]) | (t[83] & ~t[85] & t[86] & ~t[87]);
  assign t[61] = (t[68] & ~t[69] & ~t[70] & ~t[71] & ~t[72]) | (~t[67] & t[68] & ~t[70] & ~t[71] & ~t[73]) | (~t[67] & t[68] & ~t[69] & ~t[72] & ~t[73]) | (t[67] & ~t[68] & t[69] & t[70] & ~t[73]) | (t[67] & ~t[68] & t[71] & t[72] & ~t[73]) | (t[68] & ~t[70] & ~t[72] & t[73]) | (~t[68] & t[70] & t[72] & t[73]);
  assign t[62] = (t[67] & t[68] & t[69] & ~t[70] & ~t[72] & ~t[73]) | (t[68] & ~t[69] & ~t[70] & ~t[71] & t[72] & t[73]) | (~t[68] & ~t[69] & t[70] & ~t[71] & ~t[72]) | (~t[67] & ~t[69] & t[70] & ~t[72] & ~t[73]) | (~t[67] & ~t[68] & t[70] & ~t[71] & ~t[73]) | (~t[68] & t[69] & t[70] & t[71] & ~t[72]) | (~t[69] & t[70] & t[71] & ~t[73]);
  assign t[63] = (t[67] & t[68] & ~t[69] & ~t[71] & t[72] & ~t[73]) | (t[67] & t[69] & ~t[70] & ~t[71] & ~t[72] & t[73]) | (~t[68] & ~t[69] & t[71] & ~t[72] & ~t[73]) | (~t[67] & ~t[69] & ~t[70] & t[71] & ~t[72]) | (~t[67] & ~t[68] & ~t[70] & t[71] & ~t[73]) | (~t[67] & ~t[69] & t[70] & t[71] & t[72]) | (t[70] & t[71] & ~t[72] & ~t[73]);
  assign t[64] = (t[67] & t[68] & ~t[70] & t[71] & ~t[72] & ~t[73]) | (t[68] & ~t[69] & t[70] & ~t[71] & ~t[72] & t[73]) | (~t[68] & ~t[69] & ~t[70] & ~t[71] & t[72]) | (~t[67] & ~t[70] & ~t[71] & t[72] & ~t[73]) | (~t[67] & ~t[68] & ~t[69] & t[72] & ~t[73]) | (~t[68] & t[69] & ~t[70] & t[71] & t[72]) | (t[69] & ~t[71] & t[72] & ~t[73]);
  assign t[65] = (t[88] & ~t[90] & ~t[91] & ~t[92] & ~t[93]) | (t[88] & ~t[89] & ~t[91] & ~t[92] & ~t[94]) | (t[88] & ~t[89] & ~t[90] & ~t[93] & ~t[94]) | (~t[88] & t[89] & t[90] & t[91] & ~t[94]) | (~t[88] & t[89] & t[92] & t[93] & ~t[94]) | (t[88] & ~t[90] & ~t[92] & t[94]) | (~t[88] & t[90] & t[92] & t[94]);
  assign t[66] = (t[88] & t[89] & ~t[90] & ~t[92] & t[93] & ~t[94]) | (t[88] & t[90] & ~t[91] & ~t[92] & ~t[93] & t[94]) | (~t[89] & ~t[90] & t[92] & ~t[93] & ~t[94]) | (~t[88] & ~t[90] & ~t[91] & t[92] & ~t[93]) | (~t[88] & ~t[89] & ~t[91] & t[92] & ~t[94]) | (~t[88] & ~t[90] & t[91] & t[92] & t[93]) | (t[91] & t[92] & ~t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[7];
  assign t[68] = t[96] ^ x[29];
  assign t[69] = t[97] ^ x[8];
  assign t[6] = t[8] ^ t[9];
  assign t[70] = t[98] ^ x[30];
  assign t[71] = t[99] ^ x[31];
  assign t[72] = t[100] ^ x[32];
  assign t[73] = t[101] ^ x[6];
  assign t[74] = t[102] ^ x[15];
  assign t[75] = t[103] ^ x[10];
  assign t[76] = t[104] ^ x[11];
  assign t[77] = t[105] ^ x[12];
  assign t[78] = t[106] ^ x[16];
  assign t[79] = t[107] ^ x[13];
  assign t[7] = t[10] ^ t[11];
  assign t[80] = t[108] ^ x[14];
  assign t[81] = t[109] ^ x[22];
  assign t[82] = t[110] ^ x[25];
  assign t[83] = t[111] ^ x[23];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[24];
  assign t[86] = t[114] ^ x[27];
  assign t[87] = t[115] ^ x[21];
  assign t[88] = t[116] ^ x[39];
  assign t[89] = t[117] ^ x[34];
  assign t[8] = t[12] ^ t[13];
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[36];
  assign t[92] = t[120] ^ x[40];
  assign t[93] = t[121] ^ x[37];
  assign t[94] = t[122] ^ x[38];
  assign t[95] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[96] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[97] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[98] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[99] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[9] = t[14] & t[15];
  assign y = (t[0] & ~t[21]) | (~t[0] & t[21]);
endmodule

module R2ind139(x, y);
 input [40:0] x;
 output y;

 wire [115:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[101] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[102] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[103] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[104] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[105] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[106] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[107] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[108] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[109] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[10] = ~(t[26] ^ t[9]);
  assign t[110] = (x[33] & ~1'b0 & ~1'b0) | (~x[33] & 1'b0 & ~1'b0) | (~x[33] & ~1'b0 & 1'b0) | (x[33] & 1'b0 & 1'b0);
  assign t[111] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[112] = (x[33] & ~1'b0) | (~x[33] & 1'b0);
  assign t[113] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[114] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[115] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[11] = x[0] ? x[32] : t[12];
  assign t[12] = ~(t[13] ^ t[27]);
  assign t[13] = ~t[14];
  assign t[14] = ~(t[15] ^ t[28]);
  assign t[15] = ~t[16];
  assign t[16] = ~(t[17]);
  assign t[17] = t[18] ^ t[8];
  assign t[18] = t[19] ^ t[20];
  assign t[19] = t[29] ^ t[24];
  assign t[1] = ~(t[2] ^ t[22]);
  assign t[20] = t[9] & t[21];
  assign t[21] = t[26] ^ t[7];
  assign t[22] = (t[30] & ~t[32] & ~t[34]) | (~t[31] & t[32] & ~t[33]) | (~t[30] & ~t[32] & t[34]) | (t[31] & t[32] & t[33]);
  assign t[23] = (t[35] & ~t[36]) | (~t[35] & t[36]);
  assign t[24] = (t[37] & ~t[39] & ~t[41]) | (~t[38] & t[39] & ~t[40]) | (~t[37] & ~t[39] & t[41]) | (t[38] & t[39] & t[40]);
  assign t[25] = (t[37] & ~t[39] & ~t[40]) | (~t[38] & t[39] & ~t[41]) | (~t[37] & ~t[39] & t[40]) | (t[38] & t[39] & t[41]);
  assign t[26] = (t[37] & ~t[42]) | (~t[37] & t[42]);
  assign t[27] = (t[30] & ~t[32] & ~t[33]) | (~t[31] & t[32] & ~t[34]) | (~t[30] & ~t[32] & t[33]) | (t[31] & t[32] & t[34]);
  assign t[28] = (t[43] & ~t[44]) | (~t[43] & t[44]);
  assign t[29] = (t[37] & ~t[40]) | (~t[37] & t[40]);
  assign t[2] = ~t[3];
  assign t[30] = t[45] ^ x[8];
  assign t[31] = t[46] ^ x[9];
  assign t[32] = t[47] ^ x[10];
  assign t[33] = t[48] ^ x[11];
  assign t[34] = t[49] ^ x[12];
  assign t[35] = t[50] ^ x[19];
  assign t[36] = t[51] ^ x[20];
  assign t[37] = t[52] ^ x[26];
  assign t[38] = t[53] ^ x[27];
  assign t[39] = t[54] ^ x[28];
  assign t[3] = ~(t[4] ^ t[23]);
  assign t[40] = t[55] ^ x[29];
  assign t[41] = t[56] ^ x[30];
  assign t[42] = t[57] ^ x[31];
  assign t[43] = t[58] ^ x[39];
  assign t[44] = t[59] ^ x[40];
  assign t[45] = (t[60] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (t[60] & ~t[61] & ~t[63] & ~t[64] & ~t[66]) | (t[60] & ~t[61] & ~t[62] & ~t[65] & ~t[66]) | (~t[60] & t[61] & t[62] & t[63] & ~t[66]) | (~t[60] & t[61] & t[64] & t[65] & ~t[66]) | (t[60] & ~t[62] & ~t[64] & t[66]) | (~t[60] & t[62] & t[64] & t[66]);
  assign t[46] = (t[61] & ~t[62] & ~t[63] & ~t[64] & ~t[65]) | (~t[60] & t[61] & ~t[63] & ~t[64] & ~t[66]) | (~t[60] & t[61] & ~t[62] & ~t[65] & ~t[66]) | (t[60] & ~t[61] & t[62] & t[63] & ~t[66]) | (t[60] & ~t[61] & t[64] & t[65] & ~t[66]) | (t[61] & ~t[63] & ~t[65] & t[66]) | (~t[61] & t[63] & t[65] & t[66]);
  assign t[47] = (t[60] & t[61] & t[62] & ~t[63] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & ~t[63] & ~t[64] & t[65] & t[66]) | (~t[61] & ~t[62] & t[63] & ~t[64] & ~t[65]) | (~t[60] & ~t[62] & t[63] & ~t[65] & ~t[66]) | (~t[60] & ~t[61] & t[63] & ~t[64] & ~t[66]) | (~t[61] & t[62] & t[63] & t[64] & ~t[65]) | (~t[62] & t[63] & t[64] & ~t[66]);
  assign t[48] = (t[60] & t[61] & ~t[62] & ~t[64] & t[65] & ~t[66]) | (t[60] & t[62] & ~t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & t[64] & ~t[65] & ~t[66]) | (~t[60] & ~t[62] & ~t[63] & t[64] & ~t[65]) | (~t[60] & ~t[61] & ~t[63] & t[64] & ~t[66]) | (~t[60] & ~t[62] & t[63] & t[64] & t[65]) | (t[63] & t[64] & ~t[65] & ~t[66]);
  assign t[49] = (t[60] & t[61] & ~t[63] & t[64] & ~t[65] & ~t[66]) | (t[61] & ~t[62] & t[63] & ~t[64] & ~t[65] & t[66]) | (~t[61] & ~t[62] & ~t[63] & ~t[64] & t[65]) | (~t[60] & ~t[63] & ~t[64] & t[65] & ~t[66]) | (~t[60] & ~t[61] & ~t[62] & t[65] & ~t[66]) | (~t[61] & t[62] & ~t[63] & t[64] & t[65]) | (t[62] & ~t[64] & t[65] & ~t[66]);
  assign t[4] = ~t[5];
  assign t[50] = (t[67] & ~t[69] & ~t[70] & ~t[71] & ~t[72]) | (t[67] & ~t[68] & ~t[70] & ~t[71] & ~t[73]) | (t[67] & ~t[68] & ~t[69] & ~t[72] & ~t[73]) | (~t[67] & t[68] & t[69] & t[70] & ~t[73]) | (~t[67] & t[68] & t[71] & t[72] & ~t[73]) | (t[67] & ~t[69] & ~t[71] & t[73]) | (~t[67] & t[69] & t[71] & t[73]);
  assign t[51] = (t[67] & t[68] & ~t[69] & ~t[71] & t[72] & ~t[73]) | (t[67] & t[69] & ~t[70] & ~t[71] & ~t[72] & t[73]) | (~t[68] & ~t[69] & t[71] & ~t[72] & ~t[73]) | (~t[67] & ~t[69] & ~t[70] & t[71] & ~t[72]) | (~t[67] & ~t[68] & ~t[70] & t[71] & ~t[73]) | (~t[67] & ~t[69] & t[70] & t[71] & t[72]) | (t[70] & t[71] & ~t[72] & ~t[73]);
  assign t[52] = (t[74] & ~t[76] & ~t[77] & ~t[78] & ~t[79]) | (t[74] & ~t[75] & ~t[77] & ~t[78] & ~t[80]) | (t[74] & ~t[75] & ~t[76] & ~t[79] & ~t[80]) | (~t[74] & t[75] & t[76] & t[77] & ~t[80]) | (~t[74] & t[75] & t[78] & t[79] & ~t[80]) | (t[74] & ~t[76] & ~t[78] & t[80]) | (~t[74] & t[76] & t[78] & t[80]);
  assign t[53] = (t[75] & ~t[76] & ~t[77] & ~t[78] & ~t[79]) | (~t[74] & t[75] & ~t[77] & ~t[78] & ~t[80]) | (~t[74] & t[75] & ~t[76] & ~t[79] & ~t[80]) | (t[74] & ~t[75] & t[76] & t[77] & ~t[80]) | (t[74] & ~t[75] & t[78] & t[79] & ~t[80]) | (t[75] & ~t[77] & ~t[79] & t[80]) | (~t[75] & t[77] & t[79] & t[80]);
  assign t[54] = (t[74] & t[75] & t[76] & ~t[77] & ~t[79] & ~t[80]) | (t[75] & ~t[76] & ~t[77] & ~t[78] & t[79] & t[80]) | (~t[75] & ~t[76] & t[77] & ~t[78] & ~t[79]) | (~t[74] & ~t[76] & t[77] & ~t[79] & ~t[80]) | (~t[74] & ~t[75] & t[77] & ~t[78] & ~t[80]) | (~t[75] & t[76] & t[77] & t[78] & ~t[79]) | (~t[76] & t[77] & t[78] & ~t[80]);
  assign t[55] = (t[74] & t[75] & ~t[76] & ~t[78] & t[79] & ~t[80]) | (t[74] & t[76] & ~t[77] & ~t[78] & ~t[79] & t[80]) | (~t[75] & ~t[76] & t[78] & ~t[79] & ~t[80]) | (~t[74] & ~t[76] & ~t[77] & t[78] & ~t[79]) | (~t[74] & ~t[75] & ~t[77] & t[78] & ~t[80]) | (~t[74] & ~t[76] & t[77] & t[78] & t[79]) | (t[77] & t[78] & ~t[79] & ~t[80]);
  assign t[56] = (t[74] & t[75] & ~t[77] & t[78] & ~t[79] & ~t[80]) | (t[75] & ~t[76] & t[77] & ~t[78] & ~t[79] & t[80]) | (~t[75] & ~t[76] & ~t[77] & ~t[78] & t[79]) | (~t[74] & ~t[77] & ~t[78] & t[79] & ~t[80]) | (~t[74] & ~t[75] & ~t[76] & t[79] & ~t[80]) | (~t[75] & t[76] & ~t[77] & t[78] & t[79]) | (t[76] & ~t[78] & t[79] & ~t[80]);
  assign t[57] = (t[74] & t[75] & ~t[76] & t[77] & ~t[78] & ~t[80]) | (t[74] & ~t[76] & ~t[77] & t[78] & ~t[79] & t[80]) | (~t[75] & t[76] & ~t[77] & ~t[78] & ~t[80]) | (~t[74] & t[76] & ~t[77] & ~t[78] & ~t[79]) | (~t[74] & ~t[75] & t[76] & ~t[79] & ~t[80]) | (~t[74] & t[76] & t[77] & ~t[78] & t[79]) | (t[76] & ~t[77] & t[79] & ~t[80]);
  assign t[58] = (t[81] & ~t[83] & ~t[84] & ~t[85] & ~t[86]) | (t[81] & ~t[82] & ~t[84] & ~t[85] & ~t[87]) | (t[81] & ~t[82] & ~t[83] & ~t[86] & ~t[87]) | (~t[81] & t[82] & t[83] & t[84] & ~t[87]) | (~t[81] & t[82] & t[85] & t[86] & ~t[87]) | (t[81] & ~t[83] & ~t[85] & t[87]) | (~t[81] & t[83] & t[85] & t[87]);
  assign t[59] = (t[81] & t[82] & ~t[83] & ~t[85] & t[86] & ~t[87]) | (t[81] & t[83] & ~t[84] & ~t[85] & ~t[86] & t[87]) | (~t[82] & ~t[83] & t[85] & ~t[86] & ~t[87]) | (~t[81] & ~t[83] & ~t[84] & t[85] & ~t[86]) | (~t[81] & ~t[82] & ~t[84] & t[85] & ~t[87]) | (~t[81] & ~t[83] & t[84] & t[85] & t[86]) | (t[84] & t[85] & ~t[86] & ~t[87]);
  assign t[5] = ~(t[6]);
  assign t[60] = t[88] ^ x[8];
  assign t[61] = t[89] ^ x[9];
  assign t[62] = t[90] ^ x[6];
  assign t[63] = t[91] ^ x[10];
  assign t[64] = t[92] ^ x[11];
  assign t[65] = t[93] ^ x[12];
  assign t[66] = t[94] ^ x[7];
  assign t[67] = t[95] ^ x[19];
  assign t[68] = t[96] ^ x[14];
  assign t[69] = t[97] ^ x[15];
  assign t[6] = t[7] ^ t[8];
  assign t[70] = t[98] ^ x[16];
  assign t[71] = t[99] ^ x[20];
  assign t[72] = t[100] ^ x[17];
  assign t[73] = t[101] ^ x[18];
  assign t[74] = t[102] ^ x[26];
  assign t[75] = t[103] ^ x[27];
  assign t[76] = t[104] ^ x[31];
  assign t[77] = t[105] ^ x[28];
  assign t[78] = t[106] ^ x[29];
  assign t[79] = t[107] ^ x[30];
  assign t[7] = t[24] ^ t[25];
  assign t[80] = t[108] ^ x[25];
  assign t[81] = t[109] ^ x[39];
  assign t[82] = t[110] ^ x[34];
  assign t[83] = t[111] ^ x[35];
  assign t[84] = t[112] ^ x[36];
  assign t[85] = t[113] ^ x[40];
  assign t[86] = t[114] ^ x[37];
  assign t[87] = t[115] ^ x[38];
  assign t[88] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[89] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[8] = t[9] & t[10];
  assign t[90] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[91] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[92] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[93] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[94] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[95] = (x[13] & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0);
  assign t[96] = (x[13] & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0);
  assign t[97] = (x[13] & ~1'b0) | (~x[13] & 1'b0);
  assign t[98] = (x[13] & ~1'b0) | (~x[13] & 1'b0);
  assign t[99] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[9] = ~(t[24]);
  assign y = (t[0] & ~t[11]) | (~t[0] & t[11]);
endmodule

module R2ind140(x, y);
 input [47:0] x;
 output y;

 wire [202:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[8];
  assign t[101] = t[125] ^ x[14];
  assign t[102] = t[126] ^ x[15];
  assign t[103] = t[127] ^ x[21];
  assign t[104] = t[128] ^ x[22];
  assign t[105] = t[129] ^ x[28];
  assign t[106] = t[130] ^ x[29];
  assign t[107] = t[131] ^ x[30];
  assign t[108] = t[132] ^ x[31];
  assign t[109] = t[133] ^ x[32];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[134] ^ x[33];
  assign t[111] = t[135] ^ x[34];
  assign t[112] = t[136] ^ x[35];
  assign t[113] = t[137] ^ x[36];
  assign t[114] = t[138] ^ x[37];
  assign t[115] = t[139] ^ x[38];
  assign t[116] = t[140] ^ x[39];
  assign t[117] = t[141] ^ x[40];
  assign t[118] = t[142] ^ x[41];
  assign t[119] = t[143] ^ x[43];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[144] ^ x[45];
  assign t[121] = t[145] ^ x[46];
  assign t[122] = t[146] ^ x[47];
  assign t[123] = (t[147] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (t[147] & ~t[148] & ~t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[148] & ~t[149] & ~t[152] & ~t[153]) | (~t[147] & t[148] & t[149] & t[150] & ~t[153]) | (~t[147] & t[148] & t[151] & t[152] & ~t[153]) | (t[147] & ~t[149] & ~t[151] & t[153]) | (~t[147] & t[149] & t[151] & t[153]);
  assign t[124] = (t[147] & t[148] & ~t[149] & ~t[151] & t[152] & ~t[153]) | (t[147] & t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[153]) | (~t[147] & ~t[149] & ~t[150] & t[151] & ~t[152]) | (~t[147] & ~t[148] & ~t[150] & t[151] & ~t[153]) | (~t[147] & ~t[149] & t[150] & t[151] & t[152]) | (t[150] & t[151] & ~t[152] & ~t[153]);
  assign t[125] = (t[154] & ~t[156] & ~t[157] & ~t[158] & ~t[159]) | (t[154] & ~t[155] & ~t[157] & ~t[158] & ~t[160]) | (t[154] & ~t[155] & ~t[156] & ~t[159] & ~t[160]) | (~t[154] & t[155] & t[156] & t[157] & ~t[160]) | (~t[154] & t[155] & t[158] & t[159] & ~t[160]) | (t[154] & ~t[156] & ~t[158] & t[160]) | (~t[154] & t[156] & t[158] & t[160]);
  assign t[126] = (t[154] & t[155] & ~t[156] & t[157] & ~t[158] & ~t[160]) | (t[154] & ~t[156] & ~t[157] & t[158] & ~t[159] & t[160]) | (~t[155] & t[156] & ~t[157] & ~t[158] & ~t[160]) | (~t[154] & t[156] & ~t[157] & ~t[158] & ~t[159]) | (~t[154] & ~t[155] & t[156] & ~t[159] & ~t[160]) | (~t[154] & t[156] & t[157] & ~t[158] & t[159]) | (t[156] & ~t[157] & t[159] & ~t[160]);
  assign t[127] = (t[161] & ~t[163] & ~t[164] & ~t[165] & ~t[166]) | (t[161] & ~t[162] & ~t[164] & ~t[165] & ~t[167]) | (t[161] & ~t[162] & ~t[163] & ~t[166] & ~t[167]) | (~t[161] & t[162] & t[163] & t[164] & ~t[167]) | (~t[161] & t[162] & t[165] & t[166] & ~t[167]) | (t[161] & ~t[163] & ~t[165] & t[167]) | (~t[161] & t[163] & t[165] & t[167]);
  assign t[128] = (t[161] & t[162] & ~t[163] & t[164] & ~t[165] & ~t[167]) | (t[161] & ~t[163] & ~t[164] & t[165] & ~t[166] & t[167]) | (~t[162] & t[163] & ~t[164] & ~t[165] & ~t[167]) | (~t[161] & t[163] & ~t[164] & ~t[165] & ~t[166]) | (~t[161] & ~t[162] & t[163] & ~t[166] & ~t[167]) | (~t[161] & t[163] & t[164] & ~t[165] & t[166]) | (t[163] & ~t[164] & t[166] & ~t[167]);
  assign t[129] = (t[168] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (t[168] & ~t[169] & ~t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[169] & ~t[170] & ~t[173] & ~t[174]) | (~t[168] & t[169] & t[170] & t[171] & ~t[174]) | (~t[168] & t[169] & t[172] & t[173] & ~t[174]) | (t[168] & ~t[170] & ~t[172] & t[174]) | (~t[168] & t[170] & t[172] & t[174]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (t[168] & t[169] & ~t[170] & t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[170] & ~t[171] & t[172] & ~t[173] & t[174]) | (~t[169] & t[170] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[169] & t[170] & ~t[173] & ~t[174]) | (~t[168] & t[170] & t[171] & ~t[172] & t[173]) | (t[170] & ~t[171] & t[173] & ~t[174]);
  assign t[131] = (t[155] & ~t[156] & ~t[157] & ~t[158] & ~t[159]) | (~t[154] & t[155] & ~t[157] & ~t[158] & ~t[160]) | (~t[154] & t[155] & ~t[156] & ~t[159] & ~t[160]) | (t[154] & ~t[155] & t[156] & t[157] & ~t[160]) | (t[154] & ~t[155] & t[158] & t[159] & ~t[160]) | (t[155] & ~t[157] & ~t[159] & t[160]) | (~t[155] & t[157] & t[159] & t[160]);
  assign t[132] = (t[154] & t[155] & t[156] & ~t[157] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[157] & ~t[158] & t[159] & t[160]) | (~t[155] & ~t[156] & t[157] & ~t[158] & ~t[159]) | (~t[154] & ~t[156] & t[157] & ~t[159] & ~t[160]) | (~t[154] & ~t[155] & t[157] & ~t[158] & ~t[160]) | (~t[155] & t[156] & t[157] & t[158] & ~t[159]) | (~t[156] & t[157] & t[158] & ~t[160]);
  assign t[133] = (t[154] & t[155] & ~t[156] & ~t[158] & t[159] & ~t[160]) | (t[154] & t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[160]) | (~t[154] & ~t[156] & ~t[157] & t[158] & ~t[159]) | (~t[154] & ~t[155] & ~t[157] & t[158] & ~t[160]) | (~t[154] & ~t[156] & t[157] & t[158] & t[159]) | (t[157] & t[158] & ~t[159] & ~t[160]);
  assign t[134] = (t[154] & t[155] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[156] & ~t[157] & ~t[158] & t[159]) | (~t[154] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[154] & ~t[155] & ~t[156] & t[159] & ~t[160]) | (~t[155] & t[156] & ~t[157] & t[158] & t[159]) | (t[156] & ~t[158] & t[159] & ~t[160]);
  assign t[135] = (t[162] & ~t[163] & ~t[164] & ~t[165] & ~t[166]) | (~t[161] & t[162] & ~t[164] & ~t[165] & ~t[167]) | (~t[161] & t[162] & ~t[163] & ~t[166] & ~t[167]) | (t[161] & ~t[162] & t[163] & t[164] & ~t[167]) | (t[161] & ~t[162] & t[165] & t[166] & ~t[167]) | (t[162] & ~t[164] & ~t[166] & t[167]) | (~t[162] & t[164] & t[166] & t[167]);
  assign t[136] = (t[161] & t[162] & t[163] & ~t[164] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & ~t[164] & ~t[165] & t[166] & t[167]) | (~t[162] & ~t[163] & t[164] & ~t[165] & ~t[166]) | (~t[161] & ~t[163] & t[164] & ~t[166] & ~t[167]) | (~t[161] & ~t[162] & t[164] & ~t[165] & ~t[167]) | (~t[162] & t[163] & t[164] & t[165] & ~t[166]) | (~t[163] & t[164] & t[165] & ~t[167]);
  assign t[137] = (t[161] & t[162] & ~t[163] & ~t[165] & t[166] & ~t[167]) | (t[161] & t[163] & ~t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[163] & t[165] & ~t[166] & ~t[167]) | (~t[161] & ~t[163] & ~t[164] & t[165] & ~t[166]) | (~t[161] & ~t[162] & ~t[164] & t[165] & ~t[167]) | (~t[161] & ~t[163] & t[164] & t[165] & t[166]) | (t[164] & t[165] & ~t[166] & ~t[167]);
  assign t[138] = (t[161] & t[162] & ~t[164] & t[165] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[163] & ~t[164] & ~t[165] & t[166]) | (~t[161] & ~t[164] & ~t[165] & t[166] & ~t[167]) | (~t[161] & ~t[162] & ~t[163] & t[166] & ~t[167]) | (~t[162] & t[163] & ~t[164] & t[165] & t[166]) | (t[163] & ~t[165] & t[166] & ~t[167]);
  assign t[139] = (t[169] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & t[169] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[169] & ~t[170] & ~t[173] & ~t[174]) | (t[168] & ~t[169] & t[170] & t[171] & ~t[174]) | (t[168] & ~t[169] & t[172] & t[173] & ~t[174]) | (t[169] & ~t[171] & ~t[173] & t[174]) | (~t[169] & t[171] & t[173] & t[174]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (t[168] & t[169] & t[170] & ~t[171] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & ~t[171] & ~t[172] & t[173] & t[174]) | (~t[169] & ~t[170] & t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[170] & t[171] & ~t[173] & ~t[174]) | (~t[168] & ~t[169] & t[171] & ~t[172] & ~t[174]) | (~t[169] & t[170] & t[171] & t[172] & ~t[173]) | (~t[170] & t[171] & t[172] & ~t[174]);
  assign t[141] = (t[168] & t[169] & ~t[170] & ~t[172] & t[173] & ~t[174]) | (t[168] & t[170] & ~t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & t[172] & ~t[173] & ~t[174]) | (~t[168] & ~t[170] & ~t[171] & t[172] & ~t[173]) | (~t[168] & ~t[169] & ~t[171] & t[172] & ~t[174]) | (~t[168] & ~t[170] & t[171] & t[172] & t[173]) | (t[171] & t[172] & ~t[173] & ~t[174]);
  assign t[142] = (t[168] & t[169] & ~t[171] & t[172] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & ~t[171] & ~t[172] & t[173]) | (~t[168] & ~t[171] & ~t[172] & t[173] & ~t[174]) | (~t[168] & ~t[169] & ~t[170] & t[173] & ~t[174]) | (~t[169] & t[170] & ~t[171] & t[172] & t[173]) | (t[170] & ~t[172] & t[173] & ~t[174]);
  assign t[143] = (t[147] & t[148] & ~t[149] & t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[149] & ~t[150] & t[151] & ~t[152] & t[153]) | (~t[148] & t[149] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[148] & t[149] & ~t[152] & ~t[153]) | (~t[147] & t[149] & t[150] & ~t[151] & t[152]) | (t[149] & ~t[150] & t[152] & ~t[153]);
  assign t[144] = (t[148] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & t[148] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[148] & ~t[149] & ~t[152] & ~t[153]) | (t[147] & ~t[148] & t[149] & t[150] & ~t[153]) | (t[147] & ~t[148] & t[151] & t[152] & ~t[153]) | (t[148] & ~t[150] & ~t[152] & t[153]) | (~t[148] & t[150] & t[152] & t[153]);
  assign t[145] = (t[147] & t[148] & t[149] & ~t[150] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[150] & ~t[151] & t[152] & t[153]) | (~t[148] & ~t[149] & t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[149] & t[150] & ~t[152] & ~t[153]) | (~t[147] & ~t[148] & t[150] & ~t[151] & ~t[153]) | (~t[148] & t[149] & t[150] & t[151] & ~t[152]) | (~t[149] & t[150] & t[151] & ~t[153]);
  assign t[146] = (t[147] & t[148] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & ~t[150] & ~t[151] & t[152]) | (~t[147] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[147] & ~t[148] & ~t[149] & t[152] & ~t[153]) | (~t[148] & t[149] & ~t[150] & t[151] & t[152]) | (t[149] & ~t[151] & t[152] & ~t[153]);
  assign t[147] = t[175] ^ x[7];
  assign t[148] = t[176] ^ x[45];
  assign t[149] = t[177] ^ x[43];
  assign t[14] = t[85] & t[26];
  assign t[150] = t[178] ^ x[46];
  assign t[151] = t[179] ^ x[8];
  assign t[152] = t[180] ^ x[47];
  assign t[153] = t[181] ^ x[6];
  assign t[154] = t[182] ^ x[14];
  assign t[155] = t[183] ^ x[30];
  assign t[156] = t[184] ^ x[15];
  assign t[157] = t[185] ^ x[31];
  assign t[158] = t[186] ^ x[32];
  assign t[159] = t[187] ^ x[33];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[188] ^ x[13];
  assign t[161] = t[189] ^ x[21];
  assign t[162] = t[190] ^ x[34];
  assign t[163] = t[191] ^ x[22];
  assign t[164] = t[192] ^ x[35];
  assign t[165] = t[193] ^ x[36];
  assign t[166] = t[194] ^ x[37];
  assign t[167] = t[195] ^ x[20];
  assign t[168] = t[196] ^ x[28];
  assign t[169] = t[197] ^ x[38];
  assign t[16] = t[29] ^ t[27];
  assign t[170] = t[198] ^ x[29];
  assign t[171] = t[199] ^ x[39];
  assign t[172] = t[200] ^ x[40];
  assign t[173] = t[201] ^ x[41];
  assign t[174] = t[202] ^ x[27];
  assign t[175] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[176] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[177] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[178] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[179] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[181] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[182] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[183] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[184] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[185] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[186] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[187] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[188] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[189] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[18] = t[86] & t[31];
  assign t[190] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[191] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[192] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[193] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[194] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[195] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[196] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[197] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[198] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[199] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[201] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[202] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[87] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[88]);
  assign t[28] = ~(t[85] ^ t[27]);
  assign t[29] = t[89] ^ t[88];
  assign t[2] = ~(t[4] ^ t[84]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[90]);
  assign t[33] = ~(t[86] ^ t[32]);
  assign t[34] = t[91] ^ t[90];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[92]);
  assign t[38] = ~(t[87] ^ t[37]);
  assign t[39] = t[93] ^ t[92];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[85] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[85] ^ t[50];
  assign t[44] = t[86] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[86] ^ t[51];
  assign t[47] = t[87] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[87] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[88] ^ t[94];
  assign t[51] = t[90] ^ t[95];
  assign t[52] = t[92] ^ t[96];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[97]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61] ^ t[62]);
  assign t[59] = ~(t[63] ^ t[64]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[65] ^ t[66]);
  assign t[61] = t[67] ^ t[15];
  assign t[62] = t[8] ^ t[68];
  assign t[63] = t[69] ^ t[19];
  assign t[64] = t[10] ^ t[70];
  assign t[65] = t[71] ^ t[23];
  assign t[66] = t[12] ^ t[72];
  assign t[67] = t[29] ^ t[42];
  assign t[68] = t[85] ^ t[27];
  assign t[69] = t[34] ^ t[45];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[86] ^ t[32];
  assign t[71] = t[39] ^ t[48];
  assign t[72] = t[87] ^ t[37];
  assign t[73] = x[0] ? x[44] : t[74];
  assign t[74] = ~(t[75] ^ t[76]);
  assign t[75] = ~(t[77] ^ t[98]);
  assign t[76] = ~(t[78] ^ t[79]);
  assign t[77] = ~t[80];
  assign t[78] = ~(t[81]);
  assign t[79] = ~(t[82]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[83]);
  assign t[81] = t[50] ^ t[15];
  assign t[82] = t[51] ^ t[19];
  assign t[83] = t[52] ^ t[23];
  assign t[84] = (t[99] & ~t[100]) | (~t[99] & t[100]);
  assign t[85] = (t[101] & ~t[102]) | (~t[101] & t[102]);
  assign t[86] = (t[103] & ~t[104]) | (~t[103] & t[104]);
  assign t[87] = (t[105] & ~t[106]) | (~t[105] & t[106]);
  assign t[88] = (t[101] & ~t[108] & ~t[110]) | (~t[107] & t[108] & ~t[109]) | (~t[101] & ~t[108] & t[110]) | (t[107] & t[108] & t[109]);
  assign t[89] = (t[101] & ~t[109]) | (~t[101] & t[109]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (t[103] & ~t[112] & ~t[114]) | (~t[111] & t[112] & ~t[113]) | (~t[103] & ~t[112] & t[114]) | (t[111] & t[112] & t[113]);
  assign t[91] = (t[103] & ~t[113]) | (~t[103] & t[113]);
  assign t[92] = (t[105] & ~t[116] & ~t[118]) | (~t[115] & t[116] & ~t[117]) | (~t[105] & ~t[116] & t[118]) | (t[115] & t[116] & t[117]);
  assign t[93] = (t[105] & ~t[117]) | (~t[105] & t[117]);
  assign t[94] = (t[101] & ~t[108] & ~t[109]) | (~t[107] & t[108] & ~t[110]) | (~t[101] & ~t[108] & t[109]) | (t[107] & t[108] & t[110]);
  assign t[95] = (t[103] & ~t[112] & ~t[113]) | (~t[111] & t[112] & ~t[114]) | (~t[103] & ~t[112] & t[113]) | (t[111] & t[112] & t[114]);
  assign t[96] = (t[105] & ~t[116] & ~t[117]) | (~t[115] & t[116] & ~t[118]) | (~t[105] & ~t[116] & t[117]) | (t[115] & t[116] & t[118]);
  assign t[97] = (t[99] & ~t[119]) | (~t[99] & t[119]);
  assign t[98] = (t[99] & ~t[121] & ~t[122]) | (~t[120] & t[121] & ~t[100]) | (~t[99] & ~t[121] & t[122]) | (t[120] & t[121] & t[100]);
  assign t[99] = t[123] ^ x[7];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[73]) | (~t[0] & t[53] & ~t[73]) | (~t[0] & ~t[53] & t[73]) | (t[0] & t[53] & t[73]);
endmodule

module R2ind141(x, y);
 input [47:0] x;
 output y;

 wire [199:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[21];
  assign t[101] = t[125] ^ x[22];
  assign t[102] = t[126] ^ x[28];
  assign t[103] = t[127] ^ x[29];
  assign t[104] = t[128] ^ x[30];
  assign t[105] = t[129] ^ x[31];
  assign t[106] = t[130] ^ x[32];
  assign t[107] = t[131] ^ x[33];
  assign t[108] = t[132] ^ x[34];
  assign t[109] = t[133] ^ x[35];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[134] ^ x[36];
  assign t[111] = t[135] ^ x[37];
  assign t[112] = t[136] ^ x[38];
  assign t[113] = t[137] ^ x[39];
  assign t[114] = t[138] ^ x[40];
  assign t[115] = t[139] ^ x[41];
  assign t[116] = t[140] ^ x[43];
  assign t[117] = t[141] ^ x[45];
  assign t[118] = t[142] ^ x[46];
  assign t[119] = t[143] ^ x[47];
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[121] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[122] = (t[151] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & ~t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[152] & ~t[153] & ~t[156] & ~t[157]) | (~t[151] & t[152] & t[153] & t[154] & ~t[157]) | (~t[151] & t[152] & t[155] & t[156] & ~t[157]) | (t[151] & ~t[153] & ~t[155] & t[157]) | (~t[151] & t[153] & t[155] & t[157]);
  assign t[123] = (t[151] & t[152] & ~t[153] & t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[153] & ~t[154] & t[155] & ~t[156] & t[157]) | (~t[152] & t[153] & ~t[154] & ~t[155] & ~t[157]) | (~t[151] & t[153] & ~t[154] & ~t[155] & ~t[156]) | (~t[151] & ~t[152] & t[153] & ~t[156] & ~t[157]) | (~t[151] & t[153] & t[154] & ~t[155] & t[156]) | (t[153] & ~t[154] & t[156] & ~t[157]);
  assign t[124] = (t[158] & ~t[160] & ~t[161] & ~t[162] & ~t[163]) | (t[158] & ~t[159] & ~t[161] & ~t[162] & ~t[164]) | (t[158] & ~t[159] & ~t[160] & ~t[163] & ~t[164]) | (~t[158] & t[159] & t[160] & t[161] & ~t[164]) | (~t[158] & t[159] & t[162] & t[163] & ~t[164]) | (t[158] & ~t[160] & ~t[162] & t[164]) | (~t[158] & t[160] & t[162] & t[164]);
  assign t[125] = (t[158] & t[159] & ~t[160] & t[161] & ~t[162] & ~t[164]) | (t[158] & ~t[160] & ~t[161] & t[162] & ~t[163] & t[164]) | (~t[159] & t[160] & ~t[161] & ~t[162] & ~t[164]) | (~t[158] & t[160] & ~t[161] & ~t[162] & ~t[163]) | (~t[158] & ~t[159] & t[160] & ~t[163] & ~t[164]) | (~t[158] & t[160] & t[161] & ~t[162] & t[163]) | (t[160] & ~t[161] & t[163] & ~t[164]);
  assign t[126] = (t[165] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (t[165] & ~t[166] & ~t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[166] & ~t[167] & ~t[170] & ~t[171]) | (~t[165] & t[166] & t[167] & t[168] & ~t[171]) | (~t[165] & t[166] & t[169] & t[170] & ~t[171]) | (t[165] & ~t[167] & ~t[169] & t[171]) | (~t[165] & t[167] & t[169] & t[171]);
  assign t[127] = (t[165] & t[166] & ~t[167] & t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[167] & ~t[168] & t[169] & ~t[170] & t[171]) | (~t[166] & t[167] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[166] & t[167] & ~t[170] & ~t[171]) | (~t[165] & t[167] & t[168] & ~t[169] & t[170]) | (t[167] & ~t[168] & t[170] & ~t[171]);
  assign t[128] = (t[152] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (~t[151] & t[152] & ~t[154] & ~t[155] & ~t[157]) | (~t[151] & t[152] & ~t[153] & ~t[156] & ~t[157]) | (t[151] & ~t[152] & t[153] & t[154] & ~t[157]) | (t[151] & ~t[152] & t[155] & t[156] & ~t[157]) | (t[152] & ~t[154] & ~t[156] & t[157]) | (~t[152] & t[154] & t[156] & t[157]);
  assign t[129] = (t[151] & t[152] & t[153] & ~t[154] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & ~t[154] & ~t[155] & t[156] & t[157]) | (~t[152] & ~t[153] & t[154] & ~t[155] & ~t[156]) | (~t[151] & ~t[153] & t[154] & ~t[156] & ~t[157]) | (~t[151] & ~t[152] & t[154] & ~t[155] & ~t[157]) | (~t[152] & t[153] & t[154] & t[155] & ~t[156]) | (~t[153] & t[154] & t[155] & ~t[157]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (t[151] & t[152] & ~t[153] & ~t[155] & t[156] & ~t[157]) | (t[151] & t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[157]) | (~t[151] & ~t[153] & ~t[154] & t[155] & ~t[156]) | (~t[151] & ~t[152] & ~t[154] & t[155] & ~t[157]) | (~t[151] & ~t[153] & t[154] & t[155] & t[156]) | (t[154] & t[155] & ~t[156] & ~t[157]);
  assign t[131] = (t[151] & t[152] & ~t[154] & t[155] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & ~t[154] & ~t[155] & t[156]) | (~t[151] & ~t[154] & ~t[155] & t[156] & ~t[157]) | (~t[151] & ~t[152] & ~t[153] & t[156] & ~t[157]) | (~t[152] & t[153] & ~t[154] & t[155] & t[156]) | (t[153] & ~t[155] & t[156] & ~t[157]);
  assign t[132] = (t[159] & ~t[160] & ~t[161] & ~t[162] & ~t[163]) | (~t[158] & t[159] & ~t[161] & ~t[162] & ~t[164]) | (~t[158] & t[159] & ~t[160] & ~t[163] & ~t[164]) | (t[158] & ~t[159] & t[160] & t[161] & ~t[164]) | (t[158] & ~t[159] & t[162] & t[163] & ~t[164]) | (t[159] & ~t[161] & ~t[163] & t[164]) | (~t[159] & t[161] & t[163] & t[164]);
  assign t[133] = (t[158] & t[159] & t[160] & ~t[161] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & ~t[161] & ~t[162] & t[163] & t[164]) | (~t[159] & ~t[160] & t[161] & ~t[162] & ~t[163]) | (~t[158] & ~t[160] & t[161] & ~t[163] & ~t[164]) | (~t[158] & ~t[159] & t[161] & ~t[162] & ~t[164]) | (~t[159] & t[160] & t[161] & t[162] & ~t[163]) | (~t[160] & t[161] & t[162] & ~t[164]);
  assign t[134] = (t[158] & t[159] & ~t[160] & ~t[162] & t[163] & ~t[164]) | (t[158] & t[160] & ~t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[160] & t[162] & ~t[163] & ~t[164]) | (~t[158] & ~t[160] & ~t[161] & t[162] & ~t[163]) | (~t[158] & ~t[159] & ~t[161] & t[162] & ~t[164]) | (~t[158] & ~t[160] & t[161] & t[162] & t[163]) | (t[161] & t[162] & ~t[163] & ~t[164]);
  assign t[135] = (t[158] & t[159] & ~t[161] & t[162] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[160] & ~t[161] & ~t[162] & t[163]) | (~t[158] & ~t[161] & ~t[162] & t[163] & ~t[164]) | (~t[158] & ~t[159] & ~t[160] & t[163] & ~t[164]) | (~t[159] & t[160] & ~t[161] & t[162] & t[163]) | (t[160] & ~t[162] & t[163] & ~t[164]);
  assign t[136] = (t[166] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & t[166] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[166] & ~t[167] & ~t[170] & ~t[171]) | (t[165] & ~t[166] & t[167] & t[168] & ~t[171]) | (t[165] & ~t[166] & t[169] & t[170] & ~t[171]) | (t[166] & ~t[168] & ~t[170] & t[171]) | (~t[166] & t[168] & t[170] & t[171]);
  assign t[137] = (t[165] & t[166] & t[167] & ~t[168] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & ~t[168] & ~t[169] & t[170] & t[171]) | (~t[166] & ~t[167] & t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[167] & t[168] & ~t[170] & ~t[171]) | (~t[165] & ~t[166] & t[168] & ~t[169] & ~t[171]) | (~t[166] & t[167] & t[168] & t[169] & ~t[170]) | (~t[167] & t[168] & t[169] & ~t[171]);
  assign t[138] = (t[165] & t[166] & ~t[167] & ~t[169] & t[170] & ~t[171]) | (t[165] & t[167] & ~t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & t[169] & ~t[170] & ~t[171]) | (~t[165] & ~t[167] & ~t[168] & t[169] & ~t[170]) | (~t[165] & ~t[166] & ~t[168] & t[169] & ~t[171]) | (~t[165] & ~t[167] & t[168] & t[169] & t[170]) | (t[168] & t[169] & ~t[170] & ~t[171]);
  assign t[139] = (t[165] & t[166] & ~t[168] & t[169] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & ~t[168] & ~t[169] & t[170]) | (~t[165] & ~t[168] & ~t[169] & t[170] & ~t[171]) | (~t[165] & ~t[166] & ~t[167] & t[170] & ~t[171]) | (~t[166] & t[167] & ~t[168] & t[169] & t[170]) | (t[167] & ~t[169] & t[170] & ~t[171]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (t[144] & t[145] & ~t[146] & t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[146] & ~t[147] & t[148] & ~t[149] & t[150]) | (~t[145] & t[146] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[145] & t[146] & ~t[149] & ~t[150]) | (~t[144] & t[146] & t[147] & ~t[148] & t[149]) | (t[146] & ~t[147] & t[149] & ~t[150]);
  assign t[141] = (t[145] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & t[145] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[145] & ~t[146] & ~t[149] & ~t[150]) | (t[144] & ~t[145] & t[146] & t[147] & ~t[150]) | (t[144] & ~t[145] & t[148] & t[149] & ~t[150]) | (t[145] & ~t[147] & ~t[149] & t[150]) | (~t[145] & t[147] & t[149] & t[150]);
  assign t[142] = (t[144] & t[145] & t[146] & ~t[147] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[147] & ~t[148] & t[149] & t[150]) | (~t[145] & ~t[146] & t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[146] & t[147] & ~t[149] & ~t[150]) | (~t[144] & ~t[145] & t[147] & ~t[148] & ~t[150]) | (~t[145] & t[146] & t[147] & t[148] & ~t[149]) | (~t[146] & t[147] & t[148] & ~t[150]);
  assign t[143] = (t[144] & t[145] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[144] & ~t[145] & ~t[146] & t[149] & ~t[150]) | (~t[145] & t[146] & ~t[147] & t[148] & t[149]) | (t[146] & ~t[148] & t[149] & ~t[150]);
  assign t[144] = t[172] ^ x[7];
  assign t[145] = t[173] ^ x[45];
  assign t[146] = t[174] ^ x[43];
  assign t[147] = t[175] ^ x[46];
  assign t[148] = t[176] ^ x[8];
  assign t[149] = t[177] ^ x[47];
  assign t[14] = t[82] & t[26];
  assign t[150] = t[178] ^ x[6];
  assign t[151] = t[179] ^ x[14];
  assign t[152] = t[180] ^ x[30];
  assign t[153] = t[181] ^ x[15];
  assign t[154] = t[182] ^ x[31];
  assign t[155] = t[183] ^ x[32];
  assign t[156] = t[184] ^ x[33];
  assign t[157] = t[185] ^ x[13];
  assign t[158] = t[186] ^ x[21];
  assign t[159] = t[187] ^ x[34];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[188] ^ x[22];
  assign t[161] = t[189] ^ x[35];
  assign t[162] = t[190] ^ x[36];
  assign t[163] = t[191] ^ x[37];
  assign t[164] = t[192] ^ x[20];
  assign t[165] = t[193] ^ x[28];
  assign t[166] = t[194] ^ x[38];
  assign t[167] = t[195] ^ x[29];
  assign t[168] = t[196] ^ x[39];
  assign t[169] = t[197] ^ x[40];
  assign t[16] = t[29] ^ t[27];
  assign t[170] = t[198] ^ x[41];
  assign t[171] = t[199] ^ x[27];
  assign t[172] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[173] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[174] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[175] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[176] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[177] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[178] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[179] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[181] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[182] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[183] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[184] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[185] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[186] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[187] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[188] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[189] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[18] = t[83] & t[31];
  assign t[190] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[191] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[192] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[193] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[194] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[195] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[196] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[197] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[198] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[199] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[84] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[85]);
  assign t[28] = ~(t[82] ^ t[27]);
  assign t[29] = t[86] ^ t[85];
  assign t[2] = ~(t[4] ^ t[81]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[87]);
  assign t[33] = ~(t[83] ^ t[32]);
  assign t[34] = t[88] ^ t[87];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[89]);
  assign t[38] = ~(t[84] ^ t[37]);
  assign t[39] = t[90] ^ t[89];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[82] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[82] ^ t[50];
  assign t[44] = t[83] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[83] ^ t[51];
  assign t[47] = t[84] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[84] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[85] ^ t[91];
  assign t[51] = t[87] ^ t[92];
  assign t[52] = t[89] ^ t[93];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[94]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61] ^ t[62]);
  assign t[59] = ~(t[63] ^ t[64]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[65] ^ t[66]);
  assign t[61] = t[67] ^ t[15];
  assign t[62] = t[8] ^ t[68];
  assign t[63] = t[69] ^ t[19];
  assign t[64] = t[10] ^ t[70];
  assign t[65] = t[71] ^ t[23];
  assign t[66] = t[12] ^ t[72];
  assign t[67] = t[29] ^ t[42];
  assign t[68] = t[82] ^ t[27];
  assign t[69] = t[34] ^ t[45];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ t[32];
  assign t[71] = t[39] ^ t[48];
  assign t[72] = t[84] ^ t[37];
  assign t[73] = x[0] ? x[44] : t[74];
  assign t[74] = ~(t[75] ^ t[76]);
  assign t[75] = ~(t[77] ^ t[95]);
  assign t[76] = ~(t[78] ^ t[79]);
  assign t[77] = ~t[80];
  assign t[78] = ~(t[61]);
  assign t[79] = ~(t[63]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[65]);
  assign t[81] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[82] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[83] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[84] = (t[102] & ~t[103]) | (~t[102] & t[103]);
  assign t[85] = (t[98] & ~t[105] & ~t[107]) | (~t[104] & t[105] & ~t[106]) | (~t[98] & ~t[105] & t[107]) | (t[104] & t[105] & t[106]);
  assign t[86] = (t[98] & ~t[106]) | (~t[98] & t[106]);
  assign t[87] = (t[100] & ~t[109] & ~t[111]) | (~t[108] & t[109] & ~t[110]) | (~t[100] & ~t[109] & t[111]) | (t[108] & t[109] & t[110]);
  assign t[88] = (t[100] & ~t[110]) | (~t[100] & t[110]);
  assign t[89] = (t[102] & ~t[113] & ~t[115]) | (~t[112] & t[113] & ~t[114]) | (~t[102] & ~t[113] & t[115]) | (t[112] & t[113] & t[114]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (t[102] & ~t[114]) | (~t[102] & t[114]);
  assign t[91] = (t[98] & ~t[105] & ~t[106]) | (~t[104] & t[105] & ~t[107]) | (~t[98] & ~t[105] & t[106]) | (t[104] & t[105] & t[107]);
  assign t[92] = (t[100] & ~t[109] & ~t[110]) | (~t[108] & t[109] & ~t[111]) | (~t[100] & ~t[109] & t[110]) | (t[108] & t[109] & t[111]);
  assign t[93] = (t[102] & ~t[113] & ~t[114]) | (~t[112] & t[113] & ~t[115]) | (~t[102] & ~t[113] & t[114]) | (t[112] & t[113] & t[115]);
  assign t[94] = (t[96] & ~t[116]) | (~t[96] & t[116]);
  assign t[95] = (t[96] & ~t[118] & ~t[97]) | (~t[117] & t[118] & ~t[119]) | (~t[96] & ~t[118] & t[97]) | (t[117] & t[118] & t[119]);
  assign t[96] = t[120] ^ x[7];
  assign t[97] = t[121] ^ x[8];
  assign t[98] = t[122] ^ x[14];
  assign t[99] = t[123] ^ x[15];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[73]) | (~t[0] & t[53] & ~t[73]) | (~t[0] & ~t[53] & t[73]) | (t[0] & t[53] & t[73]);
endmodule

module R2ind142(x, y);
 input [46:0] x;
 output y;

 wire [179:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[123] ^ x[46];
  assign t[101] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[102] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[103] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[104] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[105] = (t[138] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[139] & ~t[140] & ~t[143] & ~t[144]) | (~t[138] & t[139] & t[140] & t[141] & ~t[144]) | (~t[138] & t[139] & t[142] & t[143] & ~t[144]) | (t[138] & ~t[140] & ~t[142] & t[144]) | (~t[138] & t[140] & t[142] & t[144]);
  assign t[106] = (t[138] & t[139] & ~t[140] & t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[140] & ~t[141] & t[142] & ~t[143] & t[144]) | (~t[139] & t[140] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[139] & t[140] & ~t[143] & ~t[144]) | (~t[138] & t[140] & t[141] & ~t[142] & t[143]) | (t[140] & ~t[141] & t[143] & ~t[144]);
  assign t[107] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[108] = (t[145] & t[146] & ~t[147] & t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[147] & ~t[148] & t[149] & ~t[150] & t[151]) | (~t[146] & t[147] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[146] & t[147] & ~t[150] & ~t[151]) | (~t[145] & t[147] & t[148] & ~t[149] & t[150]) | (t[147] & ~t[148] & t[150] & ~t[151]);
  assign t[109] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[111] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[112] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[113] = (t[139] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & t[139] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[139] & ~t[140] & ~t[143] & ~t[144]) | (t[138] & ~t[139] & t[140] & t[141] & ~t[144]) | (t[138] & ~t[139] & t[142] & t[143] & ~t[144]) | (t[139] & ~t[141] & ~t[143] & t[144]) | (~t[139] & t[141] & t[143] & t[144]);
  assign t[114] = (t[138] & t[139] & t[140] & ~t[141] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & ~t[141] & ~t[142] & t[143] & t[144]) | (~t[139] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[140] & t[141] & ~t[143] & ~t[144]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[144]) | (~t[139] & t[140] & t[141] & t[142] & ~t[143]) | (~t[140] & t[141] & t[142] & ~t[144]);
  assign t[115] = (t[138] & t[139] & ~t[140] & ~t[142] & t[143] & ~t[144]) | (t[138] & t[140] & ~t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & t[142] & ~t[143] & ~t[144]) | (~t[138] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[138] & ~t[139] & ~t[141] & t[142] & ~t[144]) | (~t[138] & ~t[140] & t[141] & t[142] & t[143]) | (t[141] & t[142] & ~t[143] & ~t[144]);
  assign t[116] = (t[138] & t[139] & ~t[141] & t[142] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[141] & ~t[142] & t[143] & ~t[144]) | (~t[138] & ~t[139] & ~t[140] & t[143] & ~t[144]) | (~t[139] & t[140] & ~t[141] & t[142] & t[143]) | (t[140] & ~t[142] & t[143] & ~t[144]);
  assign t[117] = (t[146] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & t[146] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[146] & ~t[147] & ~t[150] & ~t[151]) | (t[145] & ~t[146] & t[147] & t[148] & ~t[151]) | (t[145] & ~t[146] & t[149] & t[150] & ~t[151]) | (t[146] & ~t[148] & ~t[150] & t[151]) | (~t[146] & t[148] & t[150] & t[151]);
  assign t[118] = (t[145] & t[146] & t[147] & ~t[148] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & ~t[148] & ~t[149] & t[150] & t[151]) | (~t[146] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[147] & t[148] & ~t[150] & ~t[151]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[151]) | (~t[146] & t[147] & t[148] & t[149] & ~t[150]) | (~t[147] & t[148] & t[149] & ~t[151]);
  assign t[119] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[145] & t[146] & ~t[148] & t[149] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[148] & ~t[149] & t[150] & ~t[151]) | (~t[145] & ~t[146] & ~t[147] & t[150] & ~t[151]) | (~t[146] & t[147] & ~t[148] & t[149] & t[150]) | (t[147] & ~t[149] & t[150] & ~t[151]);
  assign t[121] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[122] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[123] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[124] = t[152] ^ x[8];
  assign t[125] = t[153] ^ x[44];
  assign t[126] = t[154] ^ x[6];
  assign t[127] = t[155] ^ x[45];
  assign t[128] = t[156] ^ x[9];
  assign t[129] = t[157] ^ x[46];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[7];
  assign t[131] = t[159] ^ x[15];
  assign t[132] = t[160] ^ x[31];
  assign t[133] = t[161] ^ x[16];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = t[163] ^ x[33];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[14];
  assign t[138] = t[166] ^ x[22];
  assign t[139] = t[167] ^ x[35];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[168] ^ x[23];
  assign t[141] = t[169] ^ x[36];
  assign t[142] = t[170] ^ x[37];
  assign t[143] = t[171] ^ x[38];
  assign t[144] = t[172] ^ x[21];
  assign t[145] = t[173] ^ x[29];
  assign t[146] = t[174] ^ x[39];
  assign t[147] = t[175] ^ x[30];
  assign t[148] = t[176] ^ x[40];
  assign t[149] = t[177] ^ x[41];
  assign t[14] = t[65] & t[26];
  assign t[150] = t[178] ^ x[42];
  assign t[151] = t[179] ^ x[28];
  assign t[152] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[153] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[154] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[155] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[156] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[157] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[158] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[159] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[161] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[162] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[163] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[164] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[165] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[166] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[167] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[168] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[169] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[171] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[172] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[173] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[174] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[175] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[176] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[177] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[178] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[179] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[66] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[67] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[65] ^ t[27]);
  assign t[29] = t[69] ^ t[68];
  assign t[2] = ~(t[4] ^ t[64]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[70]);
  assign t[33] = ~(t[66] ^ t[32]);
  assign t[34] = t[71] ^ t[70];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[72]);
  assign t[38] = ~(t[67] ^ t[37]);
  assign t[39] = t[73] ^ t[72];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[65] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[65] ^ t[50];
  assign t[44] = t[66] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[66] ^ t[51];
  assign t[47] = t[67] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[67] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[68] ^ t[74];
  assign t[51] = t[70] ^ t[75];
  assign t[52] = t[72] ^ t[76];
  assign t[53] = x[0] ? x[43] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[77]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = t[50] ^ t[15];
  assign t[62] = t[51] ^ t[19];
  assign t[63] = t[52] ^ t[23];
  assign t[64] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[67] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[68] = (t[80] & ~t[87] & ~t[89]) | (~t[86] & t[87] & ~t[88]) | (~t[80] & ~t[87] & t[89]) | (t[86] & t[87] & t[88]);
  assign t[69] = (t[80] & ~t[88]) | (~t[80] & t[88]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[82] & ~t[91] & ~t[93]) | (~t[90] & t[91] & ~t[92]) | (~t[82] & ~t[91] & t[93]) | (t[90] & t[91] & t[92]);
  assign t[71] = (t[82] & ~t[92]) | (~t[82] & t[92]);
  assign t[72] = (t[84] & ~t[95] & ~t[97]) | (~t[94] & t[95] & ~t[96]) | (~t[84] & ~t[95] & t[97]) | (t[94] & t[95] & t[96]);
  assign t[73] = (t[84] & ~t[96]) | (~t[84] & t[96]);
  assign t[74] = (t[80] & ~t[87] & ~t[88]) | (~t[86] & t[87] & ~t[89]) | (~t[80] & ~t[87] & t[88]) | (t[86] & t[87] & t[89]);
  assign t[75] = (t[82] & ~t[91] & ~t[92]) | (~t[90] & t[91] & ~t[93]) | (~t[82] & ~t[91] & t[92]) | (t[90] & t[91] & t[93]);
  assign t[76] = (t[84] & ~t[95] & ~t[96]) | (~t[94] & t[95] & ~t[97]) | (~t[84] & ~t[95] & t[96]) | (t[94] & t[95] & t[97]);
  assign t[77] = (t[78] & ~t[99] & ~t[100]) | (~t[98] & t[99] & ~t[79]) | (~t[78] & ~t[99] & t[100]) | (t[98] & t[99] & t[79]);
  assign t[78] = t[101] ^ x[8];
  assign t[79] = t[102] ^ x[9];
  assign t[7] = t[12] ^ t[13];
  assign t[80] = t[103] ^ x[15];
  assign t[81] = t[104] ^ x[16];
  assign t[82] = t[105] ^ x[22];
  assign t[83] = t[106] ^ x[23];
  assign t[84] = t[107] ^ x[29];
  assign t[85] = t[108] ^ x[30];
  assign t[86] = t[109] ^ x[31];
  assign t[87] = t[110] ^ x[32];
  assign t[88] = t[111] ^ x[33];
  assign t[89] = t[112] ^ x[34];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[113] ^ x[35];
  assign t[91] = t[114] ^ x[36];
  assign t[92] = t[115] ^ x[37];
  assign t[93] = t[116] ^ x[38];
  assign t[94] = t[117] ^ x[39];
  assign t[95] = t[118] ^ x[40];
  assign t[96] = t[119] ^ x[41];
  assign t[97] = t[120] ^ x[42];
  assign t[98] = t[121] ^ x[44];
  assign t[99] = t[122] ^ x[45];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind143(x, y);
 input [46:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[123] ^ x[42];
  assign t[101] = t[124] ^ x[44];
  assign t[102] = t[125] ^ x[45];
  assign t[103] = t[126] ^ x[46];
  assign t[104] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[105] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[106] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[107] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[108] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[109] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[111] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[112] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[113] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[114] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[115] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[116] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[117] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[118] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[119] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[121] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[122] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[123] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[124] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[125] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[126] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[127] = t[155] ^ x[8];
  assign t[128] = t[156] ^ x[44];
  assign t[129] = t[157] ^ x[6];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[45];
  assign t[131] = t[159] ^ x[9];
  assign t[132] = t[160] ^ x[46];
  assign t[133] = t[161] ^ x[7];
  assign t[134] = t[162] ^ x[15];
  assign t[135] = t[163] ^ x[31];
  assign t[136] = t[164] ^ x[16];
  assign t[137] = t[165] ^ x[32];
  assign t[138] = t[166] ^ x[33];
  assign t[139] = t[167] ^ x[34];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[168] ^ x[14];
  assign t[141] = t[169] ^ x[22];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[23];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[21];
  assign t[148] = t[176] ^ x[29];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = t[68] & t[26];
  assign t[150] = t[178] ^ x[30];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[28];
  assign t[155] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[156] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[157] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[158] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[159] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[161] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[162] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[163] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[164] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[165] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[166] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[167] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[168] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[169] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[171] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[172] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[173] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[174] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[175] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[176] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[177] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[178] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[179] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[181] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[182] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[18] = t[69] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[70] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[71]);
  assign t[28] = ~(t[68] ^ t[27]);
  assign t[29] = t[72] ^ t[71];
  assign t[2] = ~(t[4] ^ t[67]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[73]);
  assign t[33] = ~(t[69] ^ t[32]);
  assign t[34] = t[74] ^ t[73];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[75]);
  assign t[38] = ~(t[70] ^ t[37]);
  assign t[39] = t[76] ^ t[75];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[68] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[68] ^ t[50];
  assign t[44] = t[69] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[69] ^ t[51];
  assign t[47] = t[70] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[70] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[71] ^ t[77];
  assign t[51] = t[73] ^ t[78];
  assign t[52] = t[75] ^ t[79];
  assign t[53] = x[0] ? x[43] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[80]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = t[64] ^ t[15];
  assign t[62] = t[65] ^ t[19];
  assign t[63] = t[66] ^ t[23];
  assign t[64] = t[29] ^ t[42];
  assign t[65] = t[34] ^ t[45];
  assign t[66] = t[39] ^ t[48];
  assign t[67] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[68] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[69] = (t[85] & ~t[86]) | (~t[85] & t[86]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[87] & ~t[88]) | (~t[87] & t[88]);
  assign t[71] = (t[83] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[83] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[72] = (t[83] & ~t[91]) | (~t[83] & t[91]);
  assign t[73] = (t[85] & ~t[94] & ~t[96]) | (~t[93] & t[94] & ~t[95]) | (~t[85] & ~t[94] & t[96]) | (t[93] & t[94] & t[95]);
  assign t[74] = (t[85] & ~t[95]) | (~t[85] & t[95]);
  assign t[75] = (t[87] & ~t[98] & ~t[100]) | (~t[97] & t[98] & ~t[99]) | (~t[87] & ~t[98] & t[100]) | (t[97] & t[98] & t[99]);
  assign t[76] = (t[87] & ~t[99]) | (~t[87] & t[99]);
  assign t[77] = (t[83] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[83] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[78] = (t[85] & ~t[94] & ~t[95]) | (~t[93] & t[94] & ~t[96]) | (~t[85] & ~t[94] & t[95]) | (t[93] & t[94] & t[96]);
  assign t[79] = (t[87] & ~t[98] & ~t[99]) | (~t[97] & t[98] & ~t[100]) | (~t[87] & ~t[98] & t[99]) | (t[97] & t[98] & t[100]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[81] & ~t[102] & ~t[82]) | (~t[101] & t[102] & ~t[103]) | (~t[81] & ~t[102] & t[82]) | (t[101] & t[102] & t[103]);
  assign t[81] = t[104] ^ x[8];
  assign t[82] = t[105] ^ x[9];
  assign t[83] = t[106] ^ x[15];
  assign t[84] = t[107] ^ x[16];
  assign t[85] = t[108] ^ x[22];
  assign t[86] = t[109] ^ x[23];
  assign t[87] = t[110] ^ x[29];
  assign t[88] = t[111] ^ x[30];
  assign t[89] = t[112] ^ x[31];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[113] ^ x[32];
  assign t[91] = t[114] ^ x[33];
  assign t[92] = t[115] ^ x[34];
  assign t[93] = t[116] ^ x[35];
  assign t[94] = t[117] ^ x[36];
  assign t[95] = t[118] ^ x[37];
  assign t[96] = t[119] ^ x[38];
  assign t[97] = t[120] ^ x[39];
  assign t[98] = t[121] ^ x[40];
  assign t[99] = t[122] ^ x[41];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind144(x, y);
 input [46:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[45];
  assign t[101] = t[125] ^ x[46];
  assign t[102] = (t[126] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & ~t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[127] & ~t[128] & ~t[131] & ~t[132]) | (~t[126] & t[127] & t[128] & t[129] & ~t[132]) | (~t[126] & t[127] & t[130] & t[131] & ~t[132]) | (t[126] & ~t[128] & ~t[130] & t[132]) | (~t[126] & t[128] & t[130] & t[132]);
  assign t[103] = (t[126] & t[127] & ~t[128] & t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[128] & ~t[129] & t[130] & ~t[131] & t[132]) | (~t[127] & t[128] & ~t[129] & ~t[130] & ~t[132]) | (~t[126] & t[128] & ~t[129] & ~t[130] & ~t[131]) | (~t[126] & ~t[127] & t[128] & ~t[131] & ~t[132]) | (~t[126] & t[128] & t[129] & ~t[130] & t[131]) | (t[128] & ~t[129] & t[131] & ~t[132]);
  assign t[104] = (t[133] & ~t[135] & ~t[136] & ~t[137] & ~t[138]) | (t[133] & ~t[134] & ~t[136] & ~t[137] & ~t[139]) | (t[133] & ~t[134] & ~t[135] & ~t[138] & ~t[139]) | (~t[133] & t[134] & t[135] & t[136] & ~t[139]) | (~t[133] & t[134] & t[137] & t[138] & ~t[139]) | (t[133] & ~t[135] & ~t[137] & t[139]) | (~t[133] & t[135] & t[137] & t[139]);
  assign t[105] = (t[133] & t[134] & ~t[135] & t[136] & ~t[137] & ~t[139]) | (t[133] & ~t[135] & ~t[136] & t[137] & ~t[138] & t[139]) | (~t[134] & t[135] & ~t[136] & ~t[137] & ~t[139]) | (~t[133] & t[135] & ~t[136] & ~t[137] & ~t[138]) | (~t[133] & ~t[134] & t[135] & ~t[138] & ~t[139]) | (~t[133] & t[135] & t[136] & ~t[137] & t[138]) | (t[135] & ~t[136] & t[138] & ~t[139]);
  assign t[106] = (t[140] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (t[140] & ~t[141] & ~t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[141] & ~t[142] & ~t[145] & ~t[146]) | (~t[140] & t[141] & t[142] & t[143] & ~t[146]) | (~t[140] & t[141] & t[144] & t[145] & ~t[146]) | (t[140] & ~t[142] & ~t[144] & t[146]) | (~t[140] & t[142] & t[144] & t[146]);
  assign t[107] = (t[140] & t[141] & ~t[142] & t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[142] & ~t[143] & t[144] & ~t[145] & t[146]) | (~t[141] & t[142] & ~t[143] & ~t[144] & ~t[146]) | (~t[140] & t[142] & ~t[143] & ~t[144] & ~t[145]) | (~t[140] & ~t[141] & t[142] & ~t[145] & ~t[146]) | (~t[140] & t[142] & t[143] & ~t[144] & t[145]) | (t[142] & ~t[143] & t[145] & ~t[146]);
  assign t[108] = (t[147] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (t[147] & ~t[148] & ~t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[148] & ~t[149] & ~t[152] & ~t[153]) | (~t[147] & t[148] & t[149] & t[150] & ~t[153]) | (~t[147] & t[148] & t[151] & t[152] & ~t[153]) | (t[147] & ~t[149] & ~t[151] & t[153]) | (~t[147] & t[149] & t[151] & t[153]);
  assign t[109] = (t[147] & t[148] & ~t[149] & t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[149] & ~t[150] & t[151] & ~t[152] & t[153]) | (~t[148] & t[149] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[148] & t[149] & ~t[152] & ~t[153]) | (~t[147] & t[149] & t[150] & ~t[151] & t[152]) | (t[149] & ~t[150] & t[152] & ~t[153]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[133] & t[134] & ~t[135] & ~t[137] & t[138] & ~t[139]) | (t[133] & t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[139]) | (~t[133] & ~t[135] & ~t[136] & t[137] & ~t[138]) | (~t[133] & ~t[134] & ~t[136] & t[137] & ~t[139]) | (~t[133] & ~t[135] & t[136] & t[137] & t[138]) | (t[136] & t[137] & ~t[138] & ~t[139]);
  assign t[111] = (t[134] & ~t[135] & ~t[136] & ~t[137] & ~t[138]) | (~t[133] & t[134] & ~t[136] & ~t[137] & ~t[139]) | (~t[133] & t[134] & ~t[135] & ~t[138] & ~t[139]) | (t[133] & ~t[134] & t[135] & t[136] & ~t[139]) | (t[133] & ~t[134] & t[137] & t[138] & ~t[139]) | (t[134] & ~t[136] & ~t[138] & t[139]) | (~t[134] & t[136] & t[138] & t[139]);
  assign t[112] = (t[133] & t[134] & t[135] & ~t[136] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[136] & ~t[137] & t[138] & t[139]) | (~t[134] & ~t[135] & t[136] & ~t[137] & ~t[138]) | (~t[133] & ~t[135] & t[136] & ~t[138] & ~t[139]) | (~t[133] & ~t[134] & t[136] & ~t[137] & ~t[139]) | (~t[134] & t[135] & t[136] & t[137] & ~t[138]) | (~t[135] & t[136] & t[137] & ~t[139]);
  assign t[113] = (t[133] & t[134] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[135] & ~t[136] & ~t[137] & t[138]) | (~t[133] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[133] & ~t[134] & ~t[135] & t[138] & ~t[139]) | (~t[134] & t[135] & ~t[136] & t[137] & t[138]) | (t[135] & ~t[137] & t[138] & ~t[139]);
  assign t[114] = (t[140] & t[141] & ~t[142] & ~t[144] & t[145] & ~t[146]) | (t[140] & t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[146]) | (~t[140] & ~t[142] & ~t[143] & t[144] & ~t[145]) | (~t[140] & ~t[141] & ~t[143] & t[144] & ~t[146]) | (~t[140] & ~t[142] & t[143] & t[144] & t[145]) | (t[143] & t[144] & ~t[145] & ~t[146]);
  assign t[115] = (t[141] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (~t[140] & t[141] & ~t[143] & ~t[144] & ~t[146]) | (~t[140] & t[141] & ~t[142] & ~t[145] & ~t[146]) | (t[140] & ~t[141] & t[142] & t[143] & ~t[146]) | (t[140] & ~t[141] & t[144] & t[145] & ~t[146]) | (t[141] & ~t[143] & ~t[145] & t[146]) | (~t[141] & t[143] & t[145] & t[146]);
  assign t[116] = (t[140] & t[141] & t[142] & ~t[143] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[143] & ~t[144] & t[145] & t[146]) | (~t[141] & ~t[142] & t[143] & ~t[144] & ~t[145]) | (~t[140] & ~t[142] & t[143] & ~t[145] & ~t[146]) | (~t[140] & ~t[141] & t[143] & ~t[144] & ~t[146]) | (~t[141] & t[142] & t[143] & t[144] & ~t[145]) | (~t[142] & t[143] & t[144] & ~t[146]);
  assign t[117] = (t[140] & t[141] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & ~t[143] & ~t[144] & t[145]) | (~t[140] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[140] & ~t[141] & ~t[142] & t[145] & ~t[146]) | (~t[141] & t[142] & ~t[143] & t[144] & t[145]) | (t[142] & ~t[144] & t[145] & ~t[146]);
  assign t[118] = (t[147] & t[148] & ~t[149] & ~t[151] & t[152] & ~t[153]) | (t[147] & t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[153]) | (~t[147] & ~t[149] & ~t[150] & t[151] & ~t[152]) | (~t[147] & ~t[148] & ~t[150] & t[151] & ~t[153]) | (~t[147] & ~t[149] & t[150] & t[151] & t[152]) | (t[150] & t[151] & ~t[152] & ~t[153]);
  assign t[119] = (t[148] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & t[148] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[148] & ~t[149] & ~t[152] & ~t[153]) | (t[147] & ~t[148] & t[149] & t[150] & ~t[153]) | (t[147] & ~t[148] & t[151] & t[152] & ~t[153]) | (t[148] & ~t[150] & ~t[152] & t[153]) | (~t[148] & t[150] & t[152] & t[153]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = (t[147] & t[148] & t[149] & ~t[150] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[150] & ~t[151] & t[152] & t[153]) | (~t[148] & ~t[149] & t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[149] & t[150] & ~t[152] & ~t[153]) | (~t[147] & ~t[148] & t[150] & ~t[151] & ~t[153]) | (~t[148] & t[149] & t[150] & t[151] & ~t[152]) | (~t[149] & t[150] & t[151] & ~t[153]);
  assign t[121] = (t[147] & t[148] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & ~t[150] & ~t[151] & t[152]) | (~t[147] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[147] & ~t[148] & ~t[149] & t[152] & ~t[153]) | (~t[148] & t[149] & ~t[150] & t[151] & t[152]) | (t[149] & ~t[151] & t[152] & ~t[153]);
  assign t[122] = (t[127] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (~t[126] & t[127] & ~t[129] & ~t[130] & ~t[132]) | (~t[126] & t[127] & ~t[128] & ~t[131] & ~t[132]) | (t[126] & ~t[127] & t[128] & t[129] & ~t[132]) | (t[126] & ~t[127] & t[130] & t[131] & ~t[132]) | (t[127] & ~t[129] & ~t[131] & t[132]) | (~t[127] & t[129] & t[131] & t[132]);
  assign t[123] = (t[126] & t[127] & t[128] & ~t[129] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[129] & ~t[130] & t[131] & t[132]) | (~t[127] & ~t[128] & t[129] & ~t[130] & ~t[131]) | (~t[126] & ~t[128] & t[129] & ~t[131] & ~t[132]) | (~t[126] & ~t[127] & t[129] & ~t[130] & ~t[132]) | (~t[127] & t[128] & t[129] & t[130] & ~t[131]) | (~t[128] & t[129] & t[130] & ~t[132]);
  assign t[124] = (t[126] & t[127] & ~t[128] & ~t[130] & t[131] & ~t[132]) | (t[126] & t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[132]) | (~t[126] & ~t[128] & ~t[129] & t[130] & ~t[131]) | (~t[126] & ~t[127] & ~t[129] & t[130] & ~t[132]) | (~t[126] & ~t[128] & t[129] & t[130] & t[131]) | (t[129] & t[130] & ~t[131] & ~t[132]);
  assign t[125] = (t[126] & t[127] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[126] & ~t[127] & ~t[128] & t[131] & ~t[132]) | (~t[127] & t[128] & ~t[129] & t[130] & t[131]) | (t[128] & ~t[130] & t[131] & ~t[132]);
  assign t[126] = t[154] ^ x[7];
  assign t[127] = t[155] ^ x[43];
  assign t[128] = t[156] ^ x[8];
  assign t[129] = t[157] ^ x[44];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[45];
  assign t[131] = t[159] ^ x[46];
  assign t[132] = t[160] ^ x[6];
  assign t[133] = t[161] ^ x[14];
  assign t[134] = t[162] ^ x[31];
  assign t[135] = t[163] ^ x[15];
  assign t[136] = t[164] ^ x[32];
  assign t[137] = t[165] ^ x[30];
  assign t[138] = t[166] ^ x[33];
  assign t[139] = t[167] ^ x[13];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[168] ^ x[21];
  assign t[141] = t[169] ^ x[35];
  assign t[142] = t[170] ^ x[22];
  assign t[143] = t[171] ^ x[36];
  assign t[144] = t[172] ^ x[34];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[20];
  assign t[147] = t[175] ^ x[28];
  assign t[148] = t[176] ^ x[39];
  assign t[149] = t[177] ^ x[29];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[178] ^ x[40];
  assign t[151] = t[179] ^ x[38];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[27];
  assign t[154] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[155] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[156] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[157] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[158] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[159] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[161] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[162] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[163] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[164] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[165] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[166] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[167] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[168] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[169] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[171] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[172] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[173] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[174] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[175] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[176] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[177] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[178] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[179] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[17] = t[65] ^ t[28];
  assign t[180] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[181] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[66] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[67] ^ t[38];
  assign t[26] = t[68] ^ t[69];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[69]);
  assign t[29] = ~(t[65] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[64]);
  assign t[30] = t[65] & t[42];
  assign t[31] = t[70] ^ t[71];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[71]);
  assign t[34] = ~(t[66] ^ t[33]);
  assign t[35] = t[66] & t[44];
  assign t[36] = t[72] ^ t[73];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[73]);
  assign t[39] = ~(t[67] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[67] & t[46];
  assign t[41] = t[65] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[66] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[67] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[69] ^ t[74];
  assign t[48] = t[65] ^ t[26];
  assign t[49] = t[71] ^ t[75];
  assign t[4] = ~t[7];
  assign t[50] = t[66] ^ t[31];
  assign t[51] = t[73] ^ t[76];
  assign t[52] = t[67] ^ t[36];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[77]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = ~(t[63]);
  assign t[61] = t[47] ^ t[15];
  assign t[62] = t[49] ^ t[19];
  assign t[63] = t[51] ^ t[23];
  assign t[64] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[67] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[68] = (t[80] & ~t[86]) | (~t[80] & t[86]);
  assign t[69] = (t[80] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[86]) | (~t[80] & ~t[88] & t[89]) | (t[87] & t[88] & t[86]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (t[82] & ~t[90]) | (~t[82] & t[90]);
  assign t[71] = (t[82] & ~t[92] & ~t[93]) | (~t[91] & t[92] & ~t[90]) | (~t[82] & ~t[92] & t[93]) | (t[91] & t[92] & t[90]);
  assign t[72] = (t[84] & ~t[94]) | (~t[84] & t[94]);
  assign t[73] = (t[84] & ~t[96] & ~t[97]) | (~t[95] & t[96] & ~t[94]) | (~t[84] & ~t[96] & t[97]) | (t[95] & t[96] & t[94]);
  assign t[74] = (t[80] & ~t[88] & ~t[86]) | (~t[87] & t[88] & ~t[89]) | (~t[80] & ~t[88] & t[86]) | (t[87] & t[88] & t[89]);
  assign t[75] = (t[82] & ~t[92] & ~t[90]) | (~t[91] & t[92] & ~t[93]) | (~t[82] & ~t[92] & t[90]) | (t[91] & t[92] & t[93]);
  assign t[76] = (t[84] & ~t[96] & ~t[94]) | (~t[95] & t[96] & ~t[97]) | (~t[84] & ~t[96] & t[94]) | (t[95] & t[96] & t[97]);
  assign t[77] = (t[78] & ~t[99] & ~t[101]) | (~t[98] & t[99] & ~t[100]) | (~t[78] & ~t[99] & t[101]) | (t[98] & t[99] & t[100]);
  assign t[78] = t[102] ^ x[7];
  assign t[79] = t[103] ^ x[8];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[104] ^ x[14];
  assign t[81] = t[105] ^ x[15];
  assign t[82] = t[106] ^ x[21];
  assign t[83] = t[107] ^ x[22];
  assign t[84] = t[108] ^ x[28];
  assign t[85] = t[109] ^ x[29];
  assign t[86] = t[110] ^ x[30];
  assign t[87] = t[111] ^ x[31];
  assign t[88] = t[112] ^ x[32];
  assign t[89] = t[113] ^ x[33];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[114] ^ x[34];
  assign t[91] = t[115] ^ x[35];
  assign t[92] = t[116] ^ x[36];
  assign t[93] = t[117] ^ x[37];
  assign t[94] = t[118] ^ x[38];
  assign t[95] = t[119] ^ x[39];
  assign t[96] = t[120] ^ x[40];
  assign t[97] = t[121] ^ x[41];
  assign t[98] = t[122] ^ x[43];
  assign t[99] = t[123] ^ x[44];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind145(x, y);
 input [46:0] x;
 output y;

 wire [178:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & t[124] & ~t[125] & t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[125] & ~t[126] & t[127] & ~t[128] & t[129]) | (~t[124] & t[125] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[124] & t[125] & ~t[128] & ~t[129]) | (~t[123] & t[125] & t[126] & ~t[127] & t[128]) | (t[125] & ~t[126] & t[128] & ~t[129]);
  assign t[101] = (t[130] & ~t[132] & ~t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[133] & ~t[134] & ~t[136]) | (t[130] & ~t[131] & ~t[132] & ~t[135] & ~t[136]) | (~t[130] & t[131] & t[132] & t[133] & ~t[136]) | (~t[130] & t[131] & t[134] & t[135] & ~t[136]) | (t[130] & ~t[132] & ~t[134] & t[136]) | (~t[130] & t[132] & t[134] & t[136]);
  assign t[102] = (t[130] & t[131] & ~t[132] & t[133] & ~t[134] & ~t[136]) | (t[130] & ~t[132] & ~t[133] & t[134] & ~t[135] & t[136]) | (~t[131] & t[132] & ~t[133] & ~t[134] & ~t[136]) | (~t[130] & t[132] & ~t[133] & ~t[134] & ~t[135]) | (~t[130] & ~t[131] & t[132] & ~t[135] & ~t[136]) | (~t[130] & t[132] & t[133] & ~t[134] & t[135]) | (t[132] & ~t[133] & t[135] & ~t[136]);
  assign t[103] = (t[137] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & ~t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[138] & ~t[139] & ~t[142] & ~t[143]) | (~t[137] & t[138] & t[139] & t[140] & ~t[143]) | (~t[137] & t[138] & t[141] & t[142] & ~t[143]) | (t[137] & ~t[139] & ~t[141] & t[143]) | (~t[137] & t[139] & t[141] & t[143]);
  assign t[104] = (t[137] & t[138] & ~t[139] & t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[139] & ~t[140] & t[141] & ~t[142] & t[143]) | (~t[138] & t[139] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[138] & t[139] & ~t[142] & ~t[143]) | (~t[137] & t[139] & t[140] & ~t[141] & t[142]) | (t[139] & ~t[140] & t[142] & ~t[143]);
  assign t[105] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[106] = (t[144] & t[145] & ~t[146] & t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[146] & ~t[147] & t[148] & ~t[149] & t[150]) | (~t[145] & t[146] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[145] & t[146] & ~t[149] & ~t[150]) | (~t[144] & t[146] & t[147] & ~t[148] & t[149]) | (t[146] & ~t[147] & t[149] & ~t[150]);
  assign t[107] = (t[130] & t[131] & ~t[132] & ~t[134] & t[135] & ~t[136]) | (t[130] & t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[136]) | (~t[130] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[130] & ~t[131] & ~t[133] & t[134] & ~t[136]) | (~t[130] & ~t[132] & t[133] & t[134] & t[135]) | (t[133] & t[134] & ~t[135] & ~t[136]);
  assign t[108] = (t[131] & ~t[132] & ~t[133] & ~t[134] & ~t[135]) | (~t[130] & t[131] & ~t[133] & ~t[134] & ~t[136]) | (~t[130] & t[131] & ~t[132] & ~t[135] & ~t[136]) | (t[130] & ~t[131] & t[132] & t[133] & ~t[136]) | (t[130] & ~t[131] & t[134] & t[135] & ~t[136]) | (t[131] & ~t[133] & ~t[135] & t[136]) | (~t[131] & t[133] & t[135] & t[136]);
  assign t[109] = (t[130] & t[131] & t[132] & ~t[133] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[133] & ~t[134] & t[135] & t[136]) | (~t[131] & ~t[132] & t[133] & ~t[134] & ~t[135]) | (~t[130] & ~t[132] & t[133] & ~t[135] & ~t[136]) | (~t[130] & ~t[131] & t[133] & ~t[134] & ~t[136]) | (~t[131] & t[132] & t[133] & t[134] & ~t[135]) | (~t[132] & t[133] & t[134] & ~t[136]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[130] & t[131] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[130] & ~t[131] & ~t[132] & t[135] & ~t[136]) | (~t[131] & t[132] & ~t[133] & t[134] & t[135]) | (t[132] & ~t[134] & t[135] & ~t[136]);
  assign t[111] = (t[137] & t[138] & ~t[139] & ~t[141] & t[142] & ~t[143]) | (t[137] & t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[143]) | (~t[137] & ~t[139] & ~t[140] & t[141] & ~t[142]) | (~t[137] & ~t[138] & ~t[140] & t[141] & ~t[143]) | (~t[137] & ~t[139] & t[140] & t[141] & t[142]) | (t[140] & t[141] & ~t[142] & ~t[143]);
  assign t[112] = (t[138] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & t[138] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[138] & ~t[139] & ~t[142] & ~t[143]) | (t[137] & ~t[138] & t[139] & t[140] & ~t[143]) | (t[137] & ~t[138] & t[141] & t[142] & ~t[143]) | (t[138] & ~t[140] & ~t[142] & t[143]) | (~t[138] & t[140] & t[142] & t[143]);
  assign t[113] = (t[137] & t[138] & t[139] & ~t[140] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[140] & ~t[141] & t[142] & t[143]) | (~t[138] & ~t[139] & t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[139] & t[140] & ~t[142] & ~t[143]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[143]) | (~t[138] & t[139] & t[140] & t[141] & ~t[142]) | (~t[139] & t[140] & t[141] & ~t[143]);
  assign t[114] = (t[137] & t[138] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[137] & ~t[138] & ~t[139] & t[142] & ~t[143]) | (~t[138] & t[139] & ~t[140] & t[141] & t[142]) | (t[139] & ~t[141] & t[142] & ~t[143]);
  assign t[115] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[116] = (t[145] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & t[145] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[145] & ~t[146] & ~t[149] & ~t[150]) | (t[144] & ~t[145] & t[146] & t[147] & ~t[150]) | (t[144] & ~t[145] & t[148] & t[149] & ~t[150]) | (t[145] & ~t[147] & ~t[149] & t[150]) | (~t[145] & t[147] & t[149] & t[150]);
  assign t[117] = (t[144] & t[145] & t[146] & ~t[147] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[147] & ~t[148] & t[149] & t[150]) | (~t[145] & ~t[146] & t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[146] & t[147] & ~t[149] & ~t[150]) | (~t[144] & ~t[145] & t[147] & ~t[148] & ~t[150]) | (~t[145] & t[146] & t[147] & t[148] & ~t[149]) | (~t[146] & t[147] & t[148] & ~t[150]);
  assign t[118] = (t[144] & t[145] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[144] & ~t[145] & ~t[146] & t[149] & ~t[150]) | (~t[145] & t[146] & ~t[147] & t[148] & t[149]) | (t[146] & ~t[148] & t[149] & ~t[150]);
  assign t[119] = (t[124] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & t[124] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[124] & ~t[125] & ~t[128] & ~t[129]) | (t[123] & ~t[124] & t[125] & t[126] & ~t[129]) | (t[123] & ~t[124] & t[127] & t[128] & ~t[129]) | (t[124] & ~t[126] & ~t[128] & t[129]) | (~t[124] & t[126] & t[128] & t[129]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = (t[123] & t[124] & t[125] & ~t[126] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[126] & ~t[127] & t[128] & t[129]) | (~t[124] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[125] & t[126] & ~t[128] & ~t[129]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[129]) | (~t[124] & t[125] & t[126] & t[127] & ~t[128]) | (~t[125] & t[126] & t[127] & ~t[129]);
  assign t[121] = (t[123] & t[124] & ~t[125] & ~t[127] & t[128] & ~t[129]) | (t[123] & t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[129]) | (~t[123] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[123] & ~t[124] & ~t[126] & t[127] & ~t[129]) | (~t[123] & ~t[125] & t[126] & t[127] & t[128]) | (t[126] & t[127] & ~t[128] & ~t[129]);
  assign t[122] = (t[123] & t[124] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[123] & ~t[124] & ~t[125] & t[128] & ~t[129]) | (~t[124] & t[125] & ~t[126] & t[127] & t[128]) | (t[125] & ~t[127] & t[128] & ~t[129]);
  assign t[123] = t[151] ^ x[7];
  assign t[124] = t[152] ^ x[43];
  assign t[125] = t[153] ^ x[8];
  assign t[126] = t[154] ^ x[44];
  assign t[127] = t[155] ^ x[45];
  assign t[128] = t[156] ^ x[46];
  assign t[129] = t[157] ^ x[6];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[14];
  assign t[131] = t[159] ^ x[31];
  assign t[132] = t[160] ^ x[15];
  assign t[133] = t[161] ^ x[32];
  assign t[134] = t[162] ^ x[30];
  assign t[135] = t[163] ^ x[33];
  assign t[136] = t[164] ^ x[13];
  assign t[137] = t[165] ^ x[21];
  assign t[138] = t[166] ^ x[35];
  assign t[139] = t[167] ^ x[22];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[168] ^ x[36];
  assign t[141] = t[169] ^ x[34];
  assign t[142] = t[170] ^ x[37];
  assign t[143] = t[171] ^ x[20];
  assign t[144] = t[172] ^ x[28];
  assign t[145] = t[173] ^ x[39];
  assign t[146] = t[174] ^ x[29];
  assign t[147] = t[175] ^ x[40];
  assign t[148] = t[176] ^ x[38];
  assign t[149] = t[177] ^ x[41];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[178] ^ x[27];
  assign t[151] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[152] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[153] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[154] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[155] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[156] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[157] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[158] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[159] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[161] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[162] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[163] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[164] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[165] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[166] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[167] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[168] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[169] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[171] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[172] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[173] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[174] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[175] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[176] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[177] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[178] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[17] = t[62] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[63] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[64] ^ t[38];
  assign t[26] = t[65] ^ t[66];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[66]);
  assign t[29] = ~(t[62] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[61]);
  assign t[30] = t[62] & t[42];
  assign t[31] = t[67] ^ t[68];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[68]);
  assign t[34] = ~(t[63] ^ t[33]);
  assign t[35] = t[63] & t[44];
  assign t[36] = t[69] ^ t[70];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[70]);
  assign t[39] = ~(t[64] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[64] & t[46];
  assign t[41] = t[62] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[63] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[64] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[66] ^ t[71];
  assign t[48] = t[62] ^ t[26];
  assign t[49] = t[68] ^ t[72];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ t[31];
  assign t[51] = t[70] ^ t[73];
  assign t[52] = t[64] ^ t[36];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[74]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[8]);
  assign t[59] = ~(t[10]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = ~(t[12]);
  assign t[61] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[62] = (t[77] & ~t[78]) | (~t[77] & t[78]);
  assign t[63] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[64] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[65] = (t[77] & ~t[83]) | (~t[77] & t[83]);
  assign t[66] = (t[77] & ~t[85] & ~t[86]) | (~t[84] & t[85] & ~t[83]) | (~t[77] & ~t[85] & t[86]) | (t[84] & t[85] & t[83]);
  assign t[67] = (t[79] & ~t[87]) | (~t[79] & t[87]);
  assign t[68] = (t[79] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[87]) | (~t[79] & ~t[89] & t[90]) | (t[88] & t[89] & t[87]);
  assign t[69] = (t[81] & ~t[91]) | (~t[81] & t[91]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (t[81] & ~t[93] & ~t[94]) | (~t[92] & t[93] & ~t[91]) | (~t[81] & ~t[93] & t[94]) | (t[92] & t[93] & t[91]);
  assign t[71] = (t[77] & ~t[85] & ~t[83]) | (~t[84] & t[85] & ~t[86]) | (~t[77] & ~t[85] & t[83]) | (t[84] & t[85] & t[86]);
  assign t[72] = (t[79] & ~t[89] & ~t[87]) | (~t[88] & t[89] & ~t[90]) | (~t[79] & ~t[89] & t[87]) | (t[88] & t[89] & t[90]);
  assign t[73] = (t[81] & ~t[93] & ~t[91]) | (~t[92] & t[93] & ~t[94]) | (~t[81] & ~t[93] & t[91]) | (t[92] & t[93] & t[94]);
  assign t[74] = (t[75] & ~t[96] & ~t[97]) | (~t[95] & t[96] & ~t[98]) | (~t[75] & ~t[96] & t[97]) | (t[95] & t[96] & t[98]);
  assign t[75] = t[99] ^ x[7];
  assign t[76] = t[100] ^ x[8];
  assign t[77] = t[101] ^ x[14];
  assign t[78] = t[102] ^ x[15];
  assign t[79] = t[103] ^ x[21];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[104] ^ x[22];
  assign t[81] = t[105] ^ x[28];
  assign t[82] = t[106] ^ x[29];
  assign t[83] = t[107] ^ x[30];
  assign t[84] = t[108] ^ x[31];
  assign t[85] = t[109] ^ x[32];
  assign t[86] = t[110] ^ x[33];
  assign t[87] = t[111] ^ x[34];
  assign t[88] = t[112] ^ x[35];
  assign t[89] = t[113] ^ x[36];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[114] ^ x[37];
  assign t[91] = t[115] ^ x[38];
  assign t[92] = t[116] ^ x[39];
  assign t[93] = t[117] ^ x[40];
  assign t[94] = t[118] ^ x[41];
  assign t[95] = t[119] ^ x[43];
  assign t[96] = t[120] ^ x[44];
  assign t[97] = t[121] ^ x[45];
  assign t[98] = t[122] ^ x[46];
  assign t[99] = (t[123] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[124] & ~t[125] & ~t[128] & ~t[129]) | (~t[123] & t[124] & t[125] & t[126] & ~t[129]) | (~t[123] & t[124] & t[127] & t[128] & ~t[129]) | (t[123] & ~t[125] & ~t[127] & t[129]) | (~t[123] & t[125] & t[127] & t[129]);
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind146(x, y);
 input [46:0] x;
 output y;

 wire [161:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[101] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[102] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[103] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[104] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[105] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[106] = t[134] ^ x[8];
  assign t[107] = t[135] ^ x[9];
  assign t[108] = t[136] ^ x[6];
  assign t[109] = t[137] ^ x[10];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[138] ^ x[11];
  assign t[111] = t[139] ^ x[12];
  assign t[112] = t[140] ^ x[7];
  assign t[113] = t[141] ^ x[18];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[43];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[17];
  assign t[11] = t[47] ^ t[48];
  assign t[120] = t[148] ^ x[28];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[44];
  assign t[123] = t[151] ^ x[30];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[27];
  assign t[127] = t[155] ^ x[38];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[45];
  assign t[12] = t[17] & t[18];
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[37];
  assign t[134] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[135] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[136] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[137] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[138] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[139] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[13] = t[49] ^ t[50];
  assign t[140] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[141] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[142] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[143] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[144] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[145] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[146] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[147] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[148] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[149] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[14] = t[19] & t[20];
  assign t[150] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[151] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[152] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[153] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[154] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[155] = (x[33] & ~x[34] & ~x[35]) | (~x[33] & x[34] & ~x[35]) | (~x[33] & ~x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[156] = (x[33] & ~x[34] & ~x[36]) | (~x[33] & x[34] & ~x[36]) | (~x[33] & ~x[34] & x[36]) | (x[33] & x[34] & x[36]);
  assign t[157] = (x[33] & ~x[35]) | (~x[33] & x[35]);
  assign t[158] = (x[33] & ~x[36]) | (~x[33] & x[36]);
  assign t[159] = (x[34] & ~x[35]) | (~x[34] & x[35]);
  assign t[15] = t[51] ^ t[52];
  assign t[160] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[161] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[47]);
  assign t[18] = ~(t[53] ^ t[17]);
  assign t[19] = ~(t[49]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[54] ^ t[19]);
  assign t[21] = ~(t[51]);
  assign t[22] = ~(t[55] ^ t[21]);
  assign t[23] = x[0] ? x[46] : t[24];
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~(t[27] ^ t[56]);
  assign t[26] = ~(t[28] ^ t[29]);
  assign t[27] = ~t[30];
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[4] ^ t[46]);
  assign t[30] = ~(t[33]);
  assign t[31] = t[34] ^ t[12];
  assign t[32] = t[35] ^ t[14];
  assign t[33] = t[36] ^ t[16];
  assign t[34] = t[37] ^ t[38];
  assign t[35] = t[39] ^ t[40];
  assign t[36] = t[41] ^ t[42];
  assign t[37] = t[57] ^ t[47];
  assign t[38] = t[17] & t[43];
  assign t[39] = t[58] ^ t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[19] & t[44];
  assign t[41] = t[59] ^ t[51];
  assign t[42] = t[21] & t[45];
  assign t[43] = t[53] ^ t[11];
  assign t[44] = t[54] ^ t[13];
  assign t[45] = t[55] ^ t[15];
  assign t[46] = (t[60] & ~t[62] & ~t[64]) | (~t[61] & t[62] & ~t[63]) | (~t[60] & ~t[62] & t[64]) | (t[61] & t[62] & t[63]);
  assign t[47] = (t[65] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[65] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[48] = (t[65] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[65] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[49] = (t[70] & ~t[72] & ~t[74]) | (~t[71] & t[72] & ~t[73]) | (~t[70] & ~t[72] & t[74]) | (t[71] & t[72] & t[73]);
  assign t[4] = ~t[7];
  assign t[50] = (t[70] & ~t[72] & ~t[73]) | (~t[71] & t[72] & ~t[74]) | (~t[70] & ~t[72] & t[73]) | (t[71] & t[72] & t[74]);
  assign t[51] = (t[75] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[75] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[52] = (t[75] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[75] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[53] = (t[65] & ~t[80]) | (~t[65] & t[80]);
  assign t[54] = (t[70] & ~t[81]) | (~t[70] & t[81]);
  assign t[55] = (t[75] & ~t[82]) | (~t[75] & t[82]);
  assign t[56] = (t[60] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[64]) | (~t[60] & ~t[62] & t[63]) | (t[61] & t[62] & t[64]);
  assign t[57] = (t[65] & ~t[68]) | (~t[65] & t[68]);
  assign t[58] = (t[70] & ~t[73]) | (~t[70] & t[73]);
  assign t[59] = (t[75] & ~t[78]) | (~t[75] & t[78]);
  assign t[5] = ~(t[8]);
  assign t[60] = t[83] ^ x[8];
  assign t[61] = t[84] ^ x[9];
  assign t[62] = t[85] ^ x[10];
  assign t[63] = t[86] ^ x[11];
  assign t[64] = t[87] ^ x[12];
  assign t[65] = t[88] ^ x[18];
  assign t[66] = t[89] ^ x[19];
  assign t[67] = t[90] ^ x[20];
  assign t[68] = t[91] ^ x[21];
  assign t[69] = t[92] ^ x[22];
  assign t[6] = ~(t[9]);
  assign t[70] = t[93] ^ x[28];
  assign t[71] = t[94] ^ x[29];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[31];
  assign t[74] = t[97] ^ x[32];
  assign t[75] = t[98] ^ x[38];
  assign t[76] = t[99] ^ x[39];
  assign t[77] = t[100] ^ x[40];
  assign t[78] = t[101] ^ x[41];
  assign t[79] = t[102] ^ x[42];
  assign t[7] = ~(t[10]);
  assign t[80] = t[103] ^ x[43];
  assign t[81] = t[104] ^ x[44];
  assign t[82] = t[105] ^ x[45];
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[85] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[86] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[89] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[92] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[93] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[94] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[95] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[97] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[98] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[99] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0] & ~t[23]) | (~t[0] & t[23]);
endmodule

module R2ind147(x, y);
 input [47:0] x;
 output y;

 wire [203:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[7];
  assign t[101] = t[125] ^ x[8];
  assign t[102] = t[126] ^ x[14];
  assign t[103] = t[127] ^ x[15];
  assign t[104] = t[128] ^ x[21];
  assign t[105] = t[129] ^ x[22];
  assign t[106] = t[130] ^ x[28];
  assign t[107] = t[131] ^ x[29];
  assign t[108] = t[132] ^ x[30];
  assign t[109] = t[133] ^ x[31];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[134] ^ x[32];
  assign t[111] = t[135] ^ x[33];
  assign t[112] = t[136] ^ x[34];
  assign t[113] = t[137] ^ x[35];
  assign t[114] = t[138] ^ x[36];
  assign t[115] = t[139] ^ x[37];
  assign t[116] = t[140] ^ x[38];
  assign t[117] = t[141] ^ x[39];
  assign t[118] = t[142] ^ x[40];
  assign t[119] = t[143] ^ x[41];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[144] ^ x[43];
  assign t[121] = t[145] ^ x[45];
  assign t[122] = t[146] ^ x[46];
  assign t[123] = t[147] ^ x[47];
  assign t[124] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[125] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[126] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[127] = (t[155] & t[156] & ~t[157] & t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[157] & ~t[158] & t[159] & ~t[160] & t[161]) | (~t[156] & t[157] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[156] & t[157] & ~t[160] & ~t[161]) | (~t[155] & t[157] & t[158] & ~t[159] & t[160]) | (t[157] & ~t[158] & t[160] & ~t[161]);
  assign t[128] = (t[162] & ~t[164] & ~t[165] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & ~t[165] & ~t[166] & ~t[168]) | (t[162] & ~t[163] & ~t[164] & ~t[167] & ~t[168]) | (~t[162] & t[163] & t[164] & t[165] & ~t[168]) | (~t[162] & t[163] & t[166] & t[167] & ~t[168]) | (t[162] & ~t[164] & ~t[166] & t[168]) | (~t[162] & t[164] & t[166] & t[168]);
  assign t[129] = (t[162] & t[163] & ~t[164] & t[165] & ~t[166] & ~t[168]) | (t[162] & ~t[164] & ~t[165] & t[166] & ~t[167] & t[168]) | (~t[163] & t[164] & ~t[165] & ~t[166] & ~t[168]) | (~t[162] & t[164] & ~t[165] & ~t[166] & ~t[167]) | (~t[162] & ~t[163] & t[164] & ~t[167] & ~t[168]) | (~t[162] & t[164] & t[165] & ~t[166] & t[167]) | (t[164] & ~t[165] & t[167] & ~t[168]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (t[169] & ~t[171] & ~t[172] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & ~t[172] & ~t[173] & ~t[175]) | (t[169] & ~t[170] & ~t[171] & ~t[174] & ~t[175]) | (~t[169] & t[170] & t[171] & t[172] & ~t[175]) | (~t[169] & t[170] & t[173] & t[174] & ~t[175]) | (t[169] & ~t[171] & ~t[173] & t[175]) | (~t[169] & t[171] & t[173] & t[175]);
  assign t[131] = (t[169] & t[170] & ~t[171] & t[172] & ~t[173] & ~t[175]) | (t[169] & ~t[171] & ~t[172] & t[173] & ~t[174] & t[175]) | (~t[170] & t[171] & ~t[172] & ~t[173] & ~t[175]) | (~t[169] & t[171] & ~t[172] & ~t[173] & ~t[174]) | (~t[169] & ~t[170] & t[171] & ~t[174] & ~t[175]) | (~t[169] & t[171] & t[172] & ~t[173] & t[174]) | (t[171] & ~t[172] & t[174] & ~t[175]);
  assign t[132] = (t[156] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & t[156] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[156] & ~t[157] & ~t[160] & ~t[161]) | (t[155] & ~t[156] & t[157] & t[158] & ~t[161]) | (t[155] & ~t[156] & t[159] & t[160] & ~t[161]) | (t[156] & ~t[158] & ~t[160] & t[161]) | (~t[156] & t[158] & t[160] & t[161]);
  assign t[133] = (t[155] & t[156] & t[157] & ~t[158] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & ~t[158] & ~t[159] & t[160] & t[161]) | (~t[156] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[157] & t[158] & ~t[160] & ~t[161]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[161]) | (~t[156] & t[157] & t[158] & t[159] & ~t[160]) | (~t[157] & t[158] & t[159] & ~t[161]);
  assign t[134] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[135] = (t[155] & t[156] & ~t[158] & t[159] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[158] & ~t[159] & t[160] & ~t[161]) | (~t[155] & ~t[156] & ~t[157] & t[160] & ~t[161]) | (~t[156] & t[157] & ~t[158] & t[159] & t[160]) | (t[157] & ~t[159] & t[160] & ~t[161]);
  assign t[136] = (t[163] & ~t[164] & ~t[165] & ~t[166] & ~t[167]) | (~t[162] & t[163] & ~t[165] & ~t[166] & ~t[168]) | (~t[162] & t[163] & ~t[164] & ~t[167] & ~t[168]) | (t[162] & ~t[163] & t[164] & t[165] & ~t[168]) | (t[162] & ~t[163] & t[166] & t[167] & ~t[168]) | (t[163] & ~t[165] & ~t[167] & t[168]) | (~t[163] & t[165] & t[167] & t[168]);
  assign t[137] = (t[162] & t[163] & t[164] & ~t[165] & ~t[167] & ~t[168]) | (t[163] & ~t[164] & ~t[165] & ~t[166] & t[167] & t[168]) | (~t[163] & ~t[164] & t[165] & ~t[166] & ~t[167]) | (~t[162] & ~t[164] & t[165] & ~t[167] & ~t[168]) | (~t[162] & ~t[163] & t[165] & ~t[166] & ~t[168]) | (~t[163] & t[164] & t[165] & t[166] & ~t[167]) | (~t[164] & t[165] & t[166] & ~t[168]);
  assign t[138] = (t[162] & t[163] & ~t[164] & ~t[166] & t[167] & ~t[168]) | (t[162] & t[164] & ~t[165] & ~t[166] & ~t[167] & t[168]) | (~t[163] & ~t[164] & t[166] & ~t[167] & ~t[168]) | (~t[162] & ~t[164] & ~t[165] & t[166] & ~t[167]) | (~t[162] & ~t[163] & ~t[165] & t[166] & ~t[168]) | (~t[162] & ~t[164] & t[165] & t[166] & t[167]) | (t[165] & t[166] & ~t[167] & ~t[168]);
  assign t[139] = (t[162] & t[163] & ~t[165] & t[166] & ~t[167] & ~t[168]) | (t[163] & ~t[164] & t[165] & ~t[166] & ~t[167] & t[168]) | (~t[163] & ~t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[165] & ~t[166] & t[167] & ~t[168]) | (~t[162] & ~t[163] & ~t[164] & t[167] & ~t[168]) | (~t[163] & t[164] & ~t[165] & t[166] & t[167]) | (t[164] & ~t[166] & t[167] & ~t[168]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (t[170] & ~t[171] & ~t[172] & ~t[173] & ~t[174]) | (~t[169] & t[170] & ~t[172] & ~t[173] & ~t[175]) | (~t[169] & t[170] & ~t[171] & ~t[174] & ~t[175]) | (t[169] & ~t[170] & t[171] & t[172] & ~t[175]) | (t[169] & ~t[170] & t[173] & t[174] & ~t[175]) | (t[170] & ~t[172] & ~t[174] & t[175]) | (~t[170] & t[172] & t[174] & t[175]);
  assign t[141] = (t[169] & t[170] & t[171] & ~t[172] & ~t[174] & ~t[175]) | (t[170] & ~t[171] & ~t[172] & ~t[173] & t[174] & t[175]) | (~t[170] & ~t[171] & t[172] & ~t[173] & ~t[174]) | (~t[169] & ~t[171] & t[172] & ~t[174] & ~t[175]) | (~t[169] & ~t[170] & t[172] & ~t[173] & ~t[175]) | (~t[170] & t[171] & t[172] & t[173] & ~t[174]) | (~t[171] & t[172] & t[173] & ~t[175]);
  assign t[142] = (t[169] & t[170] & ~t[171] & ~t[173] & t[174] & ~t[175]) | (t[169] & t[171] & ~t[172] & ~t[173] & ~t[174] & t[175]) | (~t[170] & ~t[171] & t[173] & ~t[174] & ~t[175]) | (~t[169] & ~t[171] & ~t[172] & t[173] & ~t[174]) | (~t[169] & ~t[170] & ~t[172] & t[173] & ~t[175]) | (~t[169] & ~t[171] & t[172] & t[173] & t[174]) | (t[172] & t[173] & ~t[174] & ~t[175]);
  assign t[143] = (t[169] & t[170] & ~t[172] & t[173] & ~t[174] & ~t[175]) | (t[170] & ~t[171] & t[172] & ~t[173] & ~t[174] & t[175]) | (~t[170] & ~t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[172] & ~t[173] & t[174] & ~t[175]) | (~t[169] & ~t[170] & ~t[171] & t[174] & ~t[175]) | (~t[170] & t[171] & ~t[172] & t[173] & t[174]) | (t[171] & ~t[173] & t[174] & ~t[175]);
  assign t[144] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[145] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[146] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[147] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[148] = t[176] ^ x[7];
  assign t[149] = t[177] ^ x[45];
  assign t[14] = t[86] & t[26];
  assign t[150] = t[178] ^ x[43];
  assign t[151] = t[179] ^ x[46];
  assign t[152] = t[180] ^ x[8];
  assign t[153] = t[181] ^ x[47];
  assign t[154] = t[182] ^ x[6];
  assign t[155] = t[183] ^ x[14];
  assign t[156] = t[184] ^ x[30];
  assign t[157] = t[185] ^ x[15];
  assign t[158] = t[186] ^ x[31];
  assign t[159] = t[187] ^ x[32];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[188] ^ x[33];
  assign t[161] = t[189] ^ x[13];
  assign t[162] = t[190] ^ x[21];
  assign t[163] = t[191] ^ x[34];
  assign t[164] = t[192] ^ x[22];
  assign t[165] = t[193] ^ x[35];
  assign t[166] = t[194] ^ x[36];
  assign t[167] = t[195] ^ x[37];
  assign t[168] = t[196] ^ x[20];
  assign t[169] = t[197] ^ x[28];
  assign t[16] = t[29] ^ t[27];
  assign t[170] = t[198] ^ x[38];
  assign t[171] = t[199] ^ x[29];
  assign t[172] = t[200] ^ x[39];
  assign t[173] = t[201] ^ x[40];
  assign t[174] = t[202] ^ x[41];
  assign t[175] = t[203] ^ x[27];
  assign t[176] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[177] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[178] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[179] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[181] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[182] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[183] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[184] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[185] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[186] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[187] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[188] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[189] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[18] = t[87] & t[31];
  assign t[190] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[191] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[192] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[193] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[194] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[195] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[196] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[197] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[198] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[199] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[201] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[202] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[203] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[88] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[89]);
  assign t[28] = ~(t[86] ^ t[27]);
  assign t[29] = t[90] ^ t[89];
  assign t[2] = ~(t[4] ^ t[85]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[91]);
  assign t[33] = ~(t[87] ^ t[32]);
  assign t[34] = t[92] ^ t[91];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[93]);
  assign t[38] = ~(t[88] ^ t[37]);
  assign t[39] = t[94] ^ t[93];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[86] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[86] ^ t[50];
  assign t[44] = t[87] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[87] ^ t[51];
  assign t[47] = t[88] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[88] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[89] ^ t[95];
  assign t[51] = t[91] ^ t[96];
  assign t[52] = t[93] ^ t[97];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[98]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62] ^ t[63]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[64] ^ t[65]);
  assign t[61] = ~(t[66] ^ t[67]);
  assign t[62] = t[68] ^ t[19];
  assign t[63] = t[10] ^ t[69];
  assign t[64] = t[70] ^ t[23];
  assign t[65] = t[12] ^ t[71];
  assign t[66] = t[72] ^ t[15];
  assign t[67] = t[8] ^ t[73];
  assign t[68] = t[34] ^ t[45];
  assign t[69] = t[87] ^ t[32];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[39] ^ t[48];
  assign t[71] = t[88] ^ t[37];
  assign t[72] = t[29] ^ t[42];
  assign t[73] = t[86] ^ t[27];
  assign t[74] = x[0] ? x[44] : t[75];
  assign t[75] = ~(t[76] ^ t[77]);
  assign t[76] = ~(t[78] ^ t[99]);
  assign t[77] = ~(t[79] ^ t[80]);
  assign t[78] = ~t[81];
  assign t[79] = ~(t[82]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[83]);
  assign t[81] = ~(t[84]);
  assign t[82] = t[50] ^ t[15];
  assign t[83] = t[51] ^ t[19];
  assign t[84] = t[52] ^ t[23];
  assign t[85] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[86] = (t[102] & ~t[103]) | (~t[102] & t[103]);
  assign t[87] = (t[104] & ~t[105]) | (~t[104] & t[105]);
  assign t[88] = (t[106] & ~t[107]) | (~t[106] & t[107]);
  assign t[89] = (t[102] & ~t[109] & ~t[111]) | (~t[108] & t[109] & ~t[110]) | (~t[102] & ~t[109] & t[111]) | (t[108] & t[109] & t[110]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (t[102] & ~t[110]) | (~t[102] & t[110]);
  assign t[91] = (t[104] & ~t[113] & ~t[115]) | (~t[112] & t[113] & ~t[114]) | (~t[104] & ~t[113] & t[115]) | (t[112] & t[113] & t[114]);
  assign t[92] = (t[104] & ~t[114]) | (~t[104] & t[114]);
  assign t[93] = (t[106] & ~t[117] & ~t[119]) | (~t[116] & t[117] & ~t[118]) | (~t[106] & ~t[117] & t[119]) | (t[116] & t[117] & t[118]);
  assign t[94] = (t[106] & ~t[118]) | (~t[106] & t[118]);
  assign t[95] = (t[102] & ~t[109] & ~t[110]) | (~t[108] & t[109] & ~t[111]) | (~t[102] & ~t[109] & t[110]) | (t[108] & t[109] & t[111]);
  assign t[96] = (t[104] & ~t[113] & ~t[114]) | (~t[112] & t[113] & ~t[115]) | (~t[104] & ~t[113] & t[114]) | (t[112] & t[113] & t[115]);
  assign t[97] = (t[106] & ~t[117] & ~t[118]) | (~t[116] & t[117] & ~t[119]) | (~t[106] & ~t[117] & t[118]) | (t[116] & t[117] & t[119]);
  assign t[98] = (t[100] & ~t[120]) | (~t[100] & t[120]);
  assign t[99] = (t[100] & ~t[122] & ~t[123]) | (~t[121] & t[122] & ~t[101]) | (~t[100] & ~t[122] & t[123]) | (t[121] & t[122] & t[101]);
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[74]) | (~t[0] & t[53] & ~t[74]) | (~t[0] & ~t[53] & t[74]) | (t[0] & t[53] & t[74]);
endmodule

module R2ind148(x, y);
 input [47:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[15];
  assign t[101] = t[125] ^ x[21];
  assign t[102] = t[126] ^ x[22];
  assign t[103] = t[127] ^ x[28];
  assign t[104] = t[128] ^ x[29];
  assign t[105] = t[129] ^ x[30];
  assign t[106] = t[130] ^ x[31];
  assign t[107] = t[131] ^ x[32];
  assign t[108] = t[132] ^ x[33];
  assign t[109] = t[133] ^ x[34];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[134] ^ x[35];
  assign t[111] = t[135] ^ x[36];
  assign t[112] = t[136] ^ x[37];
  assign t[113] = t[137] ^ x[38];
  assign t[114] = t[138] ^ x[39];
  assign t[115] = t[139] ^ x[40];
  assign t[116] = t[140] ^ x[41];
  assign t[117] = t[141] ^ x[43];
  assign t[118] = t[142] ^ x[45];
  assign t[119] = t[143] ^ x[46];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[144] ^ x[47];
  assign t[121] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[122] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[123] = (t[152] & ~t[154] & ~t[155] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & ~t[155] & ~t[156] & ~t[158]) | (t[152] & ~t[153] & ~t[154] & ~t[157] & ~t[158]) | (~t[152] & t[153] & t[154] & t[155] & ~t[158]) | (~t[152] & t[153] & t[156] & t[157] & ~t[158]) | (t[152] & ~t[154] & ~t[156] & t[158]) | (~t[152] & t[154] & t[156] & t[158]);
  assign t[124] = (t[152] & t[153] & ~t[154] & t[155] & ~t[156] & ~t[158]) | (t[152] & ~t[154] & ~t[155] & t[156] & ~t[157] & t[158]) | (~t[153] & t[154] & ~t[155] & ~t[156] & ~t[158]) | (~t[152] & t[154] & ~t[155] & ~t[156] & ~t[157]) | (~t[152] & ~t[153] & t[154] & ~t[157] & ~t[158]) | (~t[152] & t[154] & t[155] & ~t[156] & t[157]) | (t[154] & ~t[155] & t[157] & ~t[158]);
  assign t[125] = (t[159] & ~t[161] & ~t[162] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & ~t[162] & ~t[163] & ~t[165]) | (t[159] & ~t[160] & ~t[161] & ~t[164] & ~t[165]) | (~t[159] & t[160] & t[161] & t[162] & ~t[165]) | (~t[159] & t[160] & t[163] & t[164] & ~t[165]) | (t[159] & ~t[161] & ~t[163] & t[165]) | (~t[159] & t[161] & t[163] & t[165]);
  assign t[126] = (t[159] & t[160] & ~t[161] & t[162] & ~t[163] & ~t[165]) | (t[159] & ~t[161] & ~t[162] & t[163] & ~t[164] & t[165]) | (~t[160] & t[161] & ~t[162] & ~t[163] & ~t[165]) | (~t[159] & t[161] & ~t[162] & ~t[163] & ~t[164]) | (~t[159] & ~t[160] & t[161] & ~t[164] & ~t[165]) | (~t[159] & t[161] & t[162] & ~t[163] & t[164]) | (t[161] & ~t[162] & t[164] & ~t[165]);
  assign t[127] = (t[166] & ~t[168] & ~t[169] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & ~t[169] & ~t[170] & ~t[172]) | (t[166] & ~t[167] & ~t[168] & ~t[171] & ~t[172]) | (~t[166] & t[167] & t[168] & t[169] & ~t[172]) | (~t[166] & t[167] & t[170] & t[171] & ~t[172]) | (t[166] & ~t[168] & ~t[170] & t[172]) | (~t[166] & t[168] & t[170] & t[172]);
  assign t[128] = (t[166] & t[167] & ~t[168] & t[169] & ~t[170] & ~t[172]) | (t[166] & ~t[168] & ~t[169] & t[170] & ~t[171] & t[172]) | (~t[167] & t[168] & ~t[169] & ~t[170] & ~t[172]) | (~t[166] & t[168] & ~t[169] & ~t[170] & ~t[171]) | (~t[166] & ~t[167] & t[168] & ~t[171] & ~t[172]) | (~t[166] & t[168] & t[169] & ~t[170] & t[171]) | (t[168] & ~t[169] & t[171] & ~t[172]);
  assign t[129] = (t[153] & ~t[154] & ~t[155] & ~t[156] & ~t[157]) | (~t[152] & t[153] & ~t[155] & ~t[156] & ~t[158]) | (~t[152] & t[153] & ~t[154] & ~t[157] & ~t[158]) | (t[152] & ~t[153] & t[154] & t[155] & ~t[158]) | (t[152] & ~t[153] & t[156] & t[157] & ~t[158]) | (t[153] & ~t[155] & ~t[157] & t[158]) | (~t[153] & t[155] & t[157] & t[158]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (t[152] & t[153] & t[154] & ~t[155] & ~t[157] & ~t[158]) | (t[153] & ~t[154] & ~t[155] & ~t[156] & t[157] & t[158]) | (~t[153] & ~t[154] & t[155] & ~t[156] & ~t[157]) | (~t[152] & ~t[154] & t[155] & ~t[157] & ~t[158]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[158]) | (~t[153] & t[154] & t[155] & t[156] & ~t[157]) | (~t[154] & t[155] & t[156] & ~t[158]);
  assign t[131] = (t[152] & t[153] & ~t[154] & ~t[156] & t[157] & ~t[158]) | (t[152] & t[154] & ~t[155] & ~t[156] & ~t[157] & t[158]) | (~t[153] & ~t[154] & t[156] & ~t[157] & ~t[158]) | (~t[152] & ~t[154] & ~t[155] & t[156] & ~t[157]) | (~t[152] & ~t[153] & ~t[155] & t[156] & ~t[158]) | (~t[152] & ~t[154] & t[155] & t[156] & t[157]) | (t[155] & t[156] & ~t[157] & ~t[158]);
  assign t[132] = (t[152] & t[153] & ~t[155] & t[156] & ~t[157] & ~t[158]) | (t[153] & ~t[154] & t[155] & ~t[156] & ~t[157] & t[158]) | (~t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[155] & ~t[156] & t[157] & ~t[158]) | (~t[152] & ~t[153] & ~t[154] & t[157] & ~t[158]) | (~t[153] & t[154] & ~t[155] & t[156] & t[157]) | (t[154] & ~t[156] & t[157] & ~t[158]);
  assign t[133] = (t[160] & ~t[161] & ~t[162] & ~t[163] & ~t[164]) | (~t[159] & t[160] & ~t[162] & ~t[163] & ~t[165]) | (~t[159] & t[160] & ~t[161] & ~t[164] & ~t[165]) | (t[159] & ~t[160] & t[161] & t[162] & ~t[165]) | (t[159] & ~t[160] & t[163] & t[164] & ~t[165]) | (t[160] & ~t[162] & ~t[164] & t[165]) | (~t[160] & t[162] & t[164] & t[165]);
  assign t[134] = (t[159] & t[160] & t[161] & ~t[162] & ~t[164] & ~t[165]) | (t[160] & ~t[161] & ~t[162] & ~t[163] & t[164] & t[165]) | (~t[160] & ~t[161] & t[162] & ~t[163] & ~t[164]) | (~t[159] & ~t[161] & t[162] & ~t[164] & ~t[165]) | (~t[159] & ~t[160] & t[162] & ~t[163] & ~t[165]) | (~t[160] & t[161] & t[162] & t[163] & ~t[164]) | (~t[161] & t[162] & t[163] & ~t[165]);
  assign t[135] = (t[159] & t[160] & ~t[161] & ~t[163] & t[164] & ~t[165]) | (t[159] & t[161] & ~t[162] & ~t[163] & ~t[164] & t[165]) | (~t[160] & ~t[161] & t[163] & ~t[164] & ~t[165]) | (~t[159] & ~t[161] & ~t[162] & t[163] & ~t[164]) | (~t[159] & ~t[160] & ~t[162] & t[163] & ~t[165]) | (~t[159] & ~t[161] & t[162] & t[163] & t[164]) | (t[162] & t[163] & ~t[164] & ~t[165]);
  assign t[136] = (t[159] & t[160] & ~t[162] & t[163] & ~t[164] & ~t[165]) | (t[160] & ~t[161] & t[162] & ~t[163] & ~t[164] & t[165]) | (~t[160] & ~t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[162] & ~t[163] & t[164] & ~t[165]) | (~t[159] & ~t[160] & ~t[161] & t[164] & ~t[165]) | (~t[160] & t[161] & ~t[162] & t[163] & t[164]) | (t[161] & ~t[163] & t[164] & ~t[165]);
  assign t[137] = (t[167] & ~t[168] & ~t[169] & ~t[170] & ~t[171]) | (~t[166] & t[167] & ~t[169] & ~t[170] & ~t[172]) | (~t[166] & t[167] & ~t[168] & ~t[171] & ~t[172]) | (t[166] & ~t[167] & t[168] & t[169] & ~t[172]) | (t[166] & ~t[167] & t[170] & t[171] & ~t[172]) | (t[167] & ~t[169] & ~t[171] & t[172]) | (~t[167] & t[169] & t[171] & t[172]);
  assign t[138] = (t[166] & t[167] & t[168] & ~t[169] & ~t[171] & ~t[172]) | (t[167] & ~t[168] & ~t[169] & ~t[170] & t[171] & t[172]) | (~t[167] & ~t[168] & t[169] & ~t[170] & ~t[171]) | (~t[166] & ~t[168] & t[169] & ~t[171] & ~t[172]) | (~t[166] & ~t[167] & t[169] & ~t[170] & ~t[172]) | (~t[167] & t[168] & t[169] & t[170] & ~t[171]) | (~t[168] & t[169] & t[170] & ~t[172]);
  assign t[139] = (t[166] & t[167] & ~t[168] & ~t[170] & t[171] & ~t[172]) | (t[166] & t[168] & ~t[169] & ~t[170] & ~t[171] & t[172]) | (~t[167] & ~t[168] & t[170] & ~t[171] & ~t[172]) | (~t[166] & ~t[168] & ~t[169] & t[170] & ~t[171]) | (~t[166] & ~t[167] & ~t[169] & t[170] & ~t[172]) | (~t[166] & ~t[168] & t[169] & t[170] & t[171]) | (t[169] & t[170] & ~t[171] & ~t[172]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (t[166] & t[167] & ~t[169] & t[170] & ~t[171] & ~t[172]) | (t[167] & ~t[168] & t[169] & ~t[170] & ~t[171] & t[172]) | (~t[167] & ~t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[169] & ~t[170] & t[171] & ~t[172]) | (~t[166] & ~t[167] & ~t[168] & t[171] & ~t[172]) | (~t[167] & t[168] & ~t[169] & t[170] & t[171]) | (t[168] & ~t[170] & t[171] & ~t[172]);
  assign t[141] = (t[145] & t[146] & ~t[147] & t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[147] & ~t[148] & t[149] & ~t[150] & t[151]) | (~t[146] & t[147] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[146] & t[147] & ~t[150] & ~t[151]) | (~t[145] & t[147] & t[148] & ~t[149] & t[150]) | (t[147] & ~t[148] & t[150] & ~t[151]);
  assign t[142] = (t[146] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & t[146] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[146] & ~t[147] & ~t[150] & ~t[151]) | (t[145] & ~t[146] & t[147] & t[148] & ~t[151]) | (t[145] & ~t[146] & t[149] & t[150] & ~t[151]) | (t[146] & ~t[148] & ~t[150] & t[151]) | (~t[146] & t[148] & t[150] & t[151]);
  assign t[143] = (t[145] & t[146] & t[147] & ~t[148] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & ~t[148] & ~t[149] & t[150] & t[151]) | (~t[146] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[147] & t[148] & ~t[150] & ~t[151]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[151]) | (~t[146] & t[147] & t[148] & t[149] & ~t[150]) | (~t[147] & t[148] & t[149] & ~t[151]);
  assign t[144] = (t[145] & t[146] & ~t[148] & t[149] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[148] & ~t[149] & t[150] & ~t[151]) | (~t[145] & ~t[146] & ~t[147] & t[150] & ~t[151]) | (~t[146] & t[147] & ~t[148] & t[149] & t[150]) | (t[147] & ~t[149] & t[150] & ~t[151]);
  assign t[145] = t[173] ^ x[7];
  assign t[146] = t[174] ^ x[45];
  assign t[147] = t[175] ^ x[43];
  assign t[148] = t[176] ^ x[46];
  assign t[149] = t[177] ^ x[8];
  assign t[14] = t[83] & t[26];
  assign t[150] = t[178] ^ x[47];
  assign t[151] = t[179] ^ x[6];
  assign t[152] = t[180] ^ x[14];
  assign t[153] = t[181] ^ x[30];
  assign t[154] = t[182] ^ x[15];
  assign t[155] = t[183] ^ x[31];
  assign t[156] = t[184] ^ x[32];
  assign t[157] = t[185] ^ x[33];
  assign t[158] = t[186] ^ x[13];
  assign t[159] = t[187] ^ x[21];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[188] ^ x[34];
  assign t[161] = t[189] ^ x[22];
  assign t[162] = t[190] ^ x[35];
  assign t[163] = t[191] ^ x[36];
  assign t[164] = t[192] ^ x[37];
  assign t[165] = t[193] ^ x[20];
  assign t[166] = t[194] ^ x[28];
  assign t[167] = t[195] ^ x[38];
  assign t[168] = t[196] ^ x[29];
  assign t[169] = t[197] ^ x[39];
  assign t[16] = t[29] ^ t[27];
  assign t[170] = t[198] ^ x[40];
  assign t[171] = t[199] ^ x[41];
  assign t[172] = t[200] ^ x[27];
  assign t[173] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[174] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[175] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[176] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[177] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[178] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[179] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[181] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[182] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[183] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[184] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[185] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[186] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[187] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[188] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[189] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[18] = t[84] & t[31];
  assign t[190] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[191] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[192] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[193] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[194] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[195] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[196] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[197] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[198] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[199] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[85] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[86]);
  assign t[28] = ~(t[83] ^ t[27]);
  assign t[29] = t[87] ^ t[86];
  assign t[2] = ~(t[4] ^ t[82]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[88]);
  assign t[33] = ~(t[84] ^ t[32]);
  assign t[34] = t[89] ^ t[88];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[90]);
  assign t[38] = ~(t[85] ^ t[37]);
  assign t[39] = t[91] ^ t[90];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[83] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[83] ^ t[50];
  assign t[44] = t[84] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[84] ^ t[51];
  assign t[47] = t[85] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[85] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[86] ^ t[92];
  assign t[51] = t[88] ^ t[93];
  assign t[52] = t[90] ^ t[94];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[95]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62] ^ t[63]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[64] ^ t[65]);
  assign t[61] = ~(t[66] ^ t[67]);
  assign t[62] = t[68] ^ t[19];
  assign t[63] = t[10] ^ t[69];
  assign t[64] = t[70] ^ t[23];
  assign t[65] = t[12] ^ t[71];
  assign t[66] = t[72] ^ t[15];
  assign t[67] = t[8] ^ t[73];
  assign t[68] = t[34] ^ t[45];
  assign t[69] = t[84] ^ t[32];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[39] ^ t[48];
  assign t[71] = t[85] ^ t[37];
  assign t[72] = t[29] ^ t[42];
  assign t[73] = t[83] ^ t[27];
  assign t[74] = x[0] ? x[44] : t[75];
  assign t[75] = ~(t[76] ^ t[77]);
  assign t[76] = ~(t[78] ^ t[96]);
  assign t[77] = ~(t[79] ^ t[80]);
  assign t[78] = ~t[81];
  assign t[79] = ~(t[66]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[62]);
  assign t[81] = ~(t[64]);
  assign t[82] = (t[97] & ~t[98]) | (~t[97] & t[98]);
  assign t[83] = (t[99] & ~t[100]) | (~t[99] & t[100]);
  assign t[84] = (t[101] & ~t[102]) | (~t[101] & t[102]);
  assign t[85] = (t[103] & ~t[104]) | (~t[103] & t[104]);
  assign t[86] = (t[99] & ~t[106] & ~t[108]) | (~t[105] & t[106] & ~t[107]) | (~t[99] & ~t[106] & t[108]) | (t[105] & t[106] & t[107]);
  assign t[87] = (t[99] & ~t[107]) | (~t[99] & t[107]);
  assign t[88] = (t[101] & ~t[110] & ~t[112]) | (~t[109] & t[110] & ~t[111]) | (~t[101] & ~t[110] & t[112]) | (t[109] & t[110] & t[111]);
  assign t[89] = (t[101] & ~t[111]) | (~t[101] & t[111]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (t[103] & ~t[114] & ~t[116]) | (~t[113] & t[114] & ~t[115]) | (~t[103] & ~t[114] & t[116]) | (t[113] & t[114] & t[115]);
  assign t[91] = (t[103] & ~t[115]) | (~t[103] & t[115]);
  assign t[92] = (t[99] & ~t[106] & ~t[107]) | (~t[105] & t[106] & ~t[108]) | (~t[99] & ~t[106] & t[107]) | (t[105] & t[106] & t[108]);
  assign t[93] = (t[101] & ~t[110] & ~t[111]) | (~t[109] & t[110] & ~t[112]) | (~t[101] & ~t[110] & t[111]) | (t[109] & t[110] & t[112]);
  assign t[94] = (t[103] & ~t[114] & ~t[115]) | (~t[113] & t[114] & ~t[116]) | (~t[103] & ~t[114] & t[115]) | (t[113] & t[114] & t[116]);
  assign t[95] = (t[97] & ~t[117]) | (~t[97] & t[117]);
  assign t[96] = (t[97] & ~t[119] & ~t[98]) | (~t[118] & t[119] & ~t[120]) | (~t[97] & ~t[119] & t[98]) | (t[118] & t[119] & t[120]);
  assign t[97] = t[121] ^ x[7];
  assign t[98] = t[122] ^ x[8];
  assign t[99] = t[123] ^ x[14];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[74]) | (~t[0] & t[53] & ~t[74]) | (~t[0] & ~t[53] & t[74]) | (t[0] & t[53] & t[74]);
endmodule

module R2ind149(x, y);
 input [46:0] x;
 output y;

 wire [179:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[123] ^ x[46];
  assign t[101] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[102] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[103] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[104] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[105] = (t[138] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[139] & ~t[140] & ~t[143] & ~t[144]) | (~t[138] & t[139] & t[140] & t[141] & ~t[144]) | (~t[138] & t[139] & t[142] & t[143] & ~t[144]) | (t[138] & ~t[140] & ~t[142] & t[144]) | (~t[138] & t[140] & t[142] & t[144]);
  assign t[106] = (t[138] & t[139] & ~t[140] & t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[140] & ~t[141] & t[142] & ~t[143] & t[144]) | (~t[139] & t[140] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[139] & t[140] & ~t[143] & ~t[144]) | (~t[138] & t[140] & t[141] & ~t[142] & t[143]) | (t[140] & ~t[141] & t[143] & ~t[144]);
  assign t[107] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[108] = (t[145] & t[146] & ~t[147] & t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[147] & ~t[148] & t[149] & ~t[150] & t[151]) | (~t[146] & t[147] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[146] & t[147] & ~t[150] & ~t[151]) | (~t[145] & t[147] & t[148] & ~t[149] & t[150]) | (t[147] & ~t[148] & t[150] & ~t[151]);
  assign t[109] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[111] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[112] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[113] = (t[139] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & t[139] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[139] & ~t[140] & ~t[143] & ~t[144]) | (t[138] & ~t[139] & t[140] & t[141] & ~t[144]) | (t[138] & ~t[139] & t[142] & t[143] & ~t[144]) | (t[139] & ~t[141] & ~t[143] & t[144]) | (~t[139] & t[141] & t[143] & t[144]);
  assign t[114] = (t[138] & t[139] & t[140] & ~t[141] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & ~t[141] & ~t[142] & t[143] & t[144]) | (~t[139] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[140] & t[141] & ~t[143] & ~t[144]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[144]) | (~t[139] & t[140] & t[141] & t[142] & ~t[143]) | (~t[140] & t[141] & t[142] & ~t[144]);
  assign t[115] = (t[138] & t[139] & ~t[140] & ~t[142] & t[143] & ~t[144]) | (t[138] & t[140] & ~t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & t[142] & ~t[143] & ~t[144]) | (~t[138] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[138] & ~t[139] & ~t[141] & t[142] & ~t[144]) | (~t[138] & ~t[140] & t[141] & t[142] & t[143]) | (t[141] & t[142] & ~t[143] & ~t[144]);
  assign t[116] = (t[138] & t[139] & ~t[141] & t[142] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[141] & ~t[142] & t[143] & ~t[144]) | (~t[138] & ~t[139] & ~t[140] & t[143] & ~t[144]) | (~t[139] & t[140] & ~t[141] & t[142] & t[143]) | (t[140] & ~t[142] & t[143] & ~t[144]);
  assign t[117] = (t[146] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & t[146] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[146] & ~t[147] & ~t[150] & ~t[151]) | (t[145] & ~t[146] & t[147] & t[148] & ~t[151]) | (t[145] & ~t[146] & t[149] & t[150] & ~t[151]) | (t[146] & ~t[148] & ~t[150] & t[151]) | (~t[146] & t[148] & t[150] & t[151]);
  assign t[118] = (t[145] & t[146] & t[147] & ~t[148] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & ~t[148] & ~t[149] & t[150] & t[151]) | (~t[146] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[147] & t[148] & ~t[150] & ~t[151]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[151]) | (~t[146] & t[147] & t[148] & t[149] & ~t[150]) | (~t[147] & t[148] & t[149] & ~t[151]);
  assign t[119] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[145] & t[146] & ~t[148] & t[149] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[148] & ~t[149] & t[150] & ~t[151]) | (~t[145] & ~t[146] & ~t[147] & t[150] & ~t[151]) | (~t[146] & t[147] & ~t[148] & t[149] & t[150]) | (t[147] & ~t[149] & t[150] & ~t[151]);
  assign t[121] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[122] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[123] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[124] = t[152] ^ x[8];
  assign t[125] = t[153] ^ x[44];
  assign t[126] = t[154] ^ x[6];
  assign t[127] = t[155] ^ x[45];
  assign t[128] = t[156] ^ x[9];
  assign t[129] = t[157] ^ x[46];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[7];
  assign t[131] = t[159] ^ x[15];
  assign t[132] = t[160] ^ x[31];
  assign t[133] = t[161] ^ x[16];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = t[163] ^ x[33];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[14];
  assign t[138] = t[166] ^ x[22];
  assign t[139] = t[167] ^ x[35];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[168] ^ x[23];
  assign t[141] = t[169] ^ x[36];
  assign t[142] = t[170] ^ x[37];
  assign t[143] = t[171] ^ x[38];
  assign t[144] = t[172] ^ x[21];
  assign t[145] = t[173] ^ x[29];
  assign t[146] = t[174] ^ x[39];
  assign t[147] = t[175] ^ x[30];
  assign t[148] = t[176] ^ x[40];
  assign t[149] = t[177] ^ x[41];
  assign t[14] = t[65] & t[26];
  assign t[150] = t[178] ^ x[42];
  assign t[151] = t[179] ^ x[28];
  assign t[152] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[153] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[154] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[155] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[156] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[157] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[158] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[159] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[161] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[162] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[163] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[164] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[165] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[166] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[167] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[168] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[169] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[171] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[172] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[173] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[174] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[175] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[176] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[177] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[178] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[179] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[66] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[67] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[65] ^ t[27]);
  assign t[29] = t[69] ^ t[68];
  assign t[2] = ~(t[4] ^ t[64]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[70]);
  assign t[33] = ~(t[66] ^ t[32]);
  assign t[34] = t[71] ^ t[70];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[72]);
  assign t[38] = ~(t[67] ^ t[37]);
  assign t[39] = t[73] ^ t[72];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[65] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[65] ^ t[50];
  assign t[44] = t[66] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[66] ^ t[51];
  assign t[47] = t[67] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[67] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[68] ^ t[74];
  assign t[51] = t[70] ^ t[75];
  assign t[52] = t[72] ^ t[76];
  assign t[53] = x[0] ? x[43] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[77]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = t[50] ^ t[15];
  assign t[62] = t[51] ^ t[19];
  assign t[63] = t[52] ^ t[23];
  assign t[64] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[67] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[68] = (t[80] & ~t[87] & ~t[89]) | (~t[86] & t[87] & ~t[88]) | (~t[80] & ~t[87] & t[89]) | (t[86] & t[87] & t[88]);
  assign t[69] = (t[80] & ~t[88]) | (~t[80] & t[88]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[82] & ~t[91] & ~t[93]) | (~t[90] & t[91] & ~t[92]) | (~t[82] & ~t[91] & t[93]) | (t[90] & t[91] & t[92]);
  assign t[71] = (t[82] & ~t[92]) | (~t[82] & t[92]);
  assign t[72] = (t[84] & ~t[95] & ~t[97]) | (~t[94] & t[95] & ~t[96]) | (~t[84] & ~t[95] & t[97]) | (t[94] & t[95] & t[96]);
  assign t[73] = (t[84] & ~t[96]) | (~t[84] & t[96]);
  assign t[74] = (t[80] & ~t[87] & ~t[88]) | (~t[86] & t[87] & ~t[89]) | (~t[80] & ~t[87] & t[88]) | (t[86] & t[87] & t[89]);
  assign t[75] = (t[82] & ~t[91] & ~t[92]) | (~t[90] & t[91] & ~t[93]) | (~t[82] & ~t[91] & t[92]) | (t[90] & t[91] & t[93]);
  assign t[76] = (t[84] & ~t[95] & ~t[96]) | (~t[94] & t[95] & ~t[97]) | (~t[84] & ~t[95] & t[96]) | (t[94] & t[95] & t[97]);
  assign t[77] = (t[78] & ~t[99] & ~t[100]) | (~t[98] & t[99] & ~t[79]) | (~t[78] & ~t[99] & t[100]) | (t[98] & t[99] & t[79]);
  assign t[78] = t[101] ^ x[8];
  assign t[79] = t[102] ^ x[9];
  assign t[7] = t[12] ^ t[13];
  assign t[80] = t[103] ^ x[15];
  assign t[81] = t[104] ^ x[16];
  assign t[82] = t[105] ^ x[22];
  assign t[83] = t[106] ^ x[23];
  assign t[84] = t[107] ^ x[29];
  assign t[85] = t[108] ^ x[30];
  assign t[86] = t[109] ^ x[31];
  assign t[87] = t[110] ^ x[32];
  assign t[88] = t[111] ^ x[33];
  assign t[89] = t[112] ^ x[34];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[113] ^ x[35];
  assign t[91] = t[114] ^ x[36];
  assign t[92] = t[115] ^ x[37];
  assign t[93] = t[116] ^ x[38];
  assign t[94] = t[117] ^ x[39];
  assign t[95] = t[118] ^ x[40];
  assign t[96] = t[119] ^ x[41];
  assign t[97] = t[120] ^ x[42];
  assign t[98] = t[121] ^ x[44];
  assign t[99] = t[122] ^ x[45];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind150(x, y);
 input [46:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[123] ^ x[42];
  assign t[101] = t[124] ^ x[44];
  assign t[102] = t[125] ^ x[45];
  assign t[103] = t[126] ^ x[46];
  assign t[104] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[105] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[106] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[107] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[108] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[109] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[111] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[112] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[113] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[114] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[115] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[116] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[117] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[118] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[119] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[121] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[122] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[123] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[124] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[125] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[126] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[127] = t[155] ^ x[8];
  assign t[128] = t[156] ^ x[44];
  assign t[129] = t[157] ^ x[6];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[45];
  assign t[131] = t[159] ^ x[9];
  assign t[132] = t[160] ^ x[46];
  assign t[133] = t[161] ^ x[7];
  assign t[134] = t[162] ^ x[15];
  assign t[135] = t[163] ^ x[31];
  assign t[136] = t[164] ^ x[16];
  assign t[137] = t[165] ^ x[32];
  assign t[138] = t[166] ^ x[33];
  assign t[139] = t[167] ^ x[34];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[168] ^ x[14];
  assign t[141] = t[169] ^ x[22];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[23];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[21];
  assign t[148] = t[176] ^ x[29];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = t[68] & t[26];
  assign t[150] = t[178] ^ x[30];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[28];
  assign t[155] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[156] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[157] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[158] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[159] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[161] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[162] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[163] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[164] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[165] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[166] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[167] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[168] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[169] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[171] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[172] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[173] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[174] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[175] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[176] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[177] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[178] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[179] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[181] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[182] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[18] = t[69] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[70] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[71]);
  assign t[28] = ~(t[68] ^ t[27]);
  assign t[29] = t[72] ^ t[71];
  assign t[2] = ~(t[4] ^ t[67]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[73]);
  assign t[33] = ~(t[69] ^ t[32]);
  assign t[34] = t[74] ^ t[73];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[75]);
  assign t[38] = ~(t[70] ^ t[37]);
  assign t[39] = t[76] ^ t[75];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[68] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[68] ^ t[50];
  assign t[44] = t[69] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[69] ^ t[51];
  assign t[47] = t[70] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[70] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[71] ^ t[77];
  assign t[51] = t[73] ^ t[78];
  assign t[52] = t[75] ^ t[79];
  assign t[53] = x[0] ? x[43] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[80]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = t[64] ^ t[15];
  assign t[62] = t[65] ^ t[19];
  assign t[63] = t[66] ^ t[23];
  assign t[64] = t[29] ^ t[42];
  assign t[65] = t[34] ^ t[45];
  assign t[66] = t[39] ^ t[48];
  assign t[67] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[68] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[69] = (t[85] & ~t[86]) | (~t[85] & t[86]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[87] & ~t[88]) | (~t[87] & t[88]);
  assign t[71] = (t[83] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[83] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[72] = (t[83] & ~t[91]) | (~t[83] & t[91]);
  assign t[73] = (t[85] & ~t[94] & ~t[96]) | (~t[93] & t[94] & ~t[95]) | (~t[85] & ~t[94] & t[96]) | (t[93] & t[94] & t[95]);
  assign t[74] = (t[85] & ~t[95]) | (~t[85] & t[95]);
  assign t[75] = (t[87] & ~t[98] & ~t[100]) | (~t[97] & t[98] & ~t[99]) | (~t[87] & ~t[98] & t[100]) | (t[97] & t[98] & t[99]);
  assign t[76] = (t[87] & ~t[99]) | (~t[87] & t[99]);
  assign t[77] = (t[83] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[83] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[78] = (t[85] & ~t[94] & ~t[95]) | (~t[93] & t[94] & ~t[96]) | (~t[85] & ~t[94] & t[95]) | (t[93] & t[94] & t[96]);
  assign t[79] = (t[87] & ~t[98] & ~t[99]) | (~t[97] & t[98] & ~t[100]) | (~t[87] & ~t[98] & t[99]) | (t[97] & t[98] & t[100]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[81] & ~t[102] & ~t[82]) | (~t[101] & t[102] & ~t[103]) | (~t[81] & ~t[102] & t[82]) | (t[101] & t[102] & t[103]);
  assign t[81] = t[104] ^ x[8];
  assign t[82] = t[105] ^ x[9];
  assign t[83] = t[106] ^ x[15];
  assign t[84] = t[107] ^ x[16];
  assign t[85] = t[108] ^ x[22];
  assign t[86] = t[109] ^ x[23];
  assign t[87] = t[110] ^ x[29];
  assign t[88] = t[111] ^ x[30];
  assign t[89] = t[112] ^ x[31];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[113] ^ x[32];
  assign t[91] = t[114] ^ x[33];
  assign t[92] = t[115] ^ x[34];
  assign t[93] = t[116] ^ x[35];
  assign t[94] = t[117] ^ x[36];
  assign t[95] = t[118] ^ x[37];
  assign t[96] = t[119] ^ x[38];
  assign t[97] = t[120] ^ x[39];
  assign t[98] = t[121] ^ x[40];
  assign t[99] = t[122] ^ x[41];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind151(x, y);
 input [46:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[44];
  assign t[101] = t[125] ^ x[45];
  assign t[102] = t[126] ^ x[46];
  assign t[103] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[104] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[105] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[106] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[107] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[108] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[109] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[10] = t[17] ^ t[18];
  assign t[110] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[111] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[112] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[113] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[114] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[115] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[116] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[117] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[118] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[119] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[121] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[122] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[123] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[124] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[125] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[126] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[127] = t[155] ^ x[7];
  assign t[128] = t[156] ^ x[43];
  assign t[129] = t[157] ^ x[8];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[158] ^ x[44];
  assign t[131] = t[159] ^ x[45];
  assign t[132] = t[160] ^ x[46];
  assign t[133] = t[161] ^ x[6];
  assign t[134] = t[162] ^ x[14];
  assign t[135] = t[163] ^ x[31];
  assign t[136] = t[164] ^ x[15];
  assign t[137] = t[165] ^ x[32];
  assign t[138] = t[166] ^ x[30];
  assign t[139] = t[167] ^ x[33];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[168] ^ x[13];
  assign t[141] = t[169] ^ x[21];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[22];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[34];
  assign t[146] = t[174] ^ x[37];
  assign t[147] = t[175] ^ x[20];
  assign t[148] = t[176] ^ x[28];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[178] ^ x[29];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[38];
  assign t[153] = t[181] ^ x[41];
  assign t[154] = t[182] ^ x[27];
  assign t[155] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[156] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[157] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[158] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[159] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[15] = t[27] ^ t[28];
  assign t[160] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[161] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[162] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[163] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[164] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[165] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[166] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[167] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[168] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[169] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[16] = t[29] & t[30];
  assign t[170] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[171] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[172] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[173] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[174] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[175] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[176] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[177] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[178] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[179] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[17] = t[31] ^ t[16];
  assign t[180] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[181] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[182] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[18] = t[66] ^ t[29];
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[67] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[68] ^ t[39];
  assign t[27] = t[69] ^ t[70];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[70]);
  assign t[2] = ~(t[4] ^ t[65]);
  assign t[30] = ~(t[66] ^ t[29]);
  assign t[31] = t[66] & t[43];
  assign t[32] = t[71] ^ t[72];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[72]);
  assign t[35] = ~(t[67] ^ t[34]);
  assign t[36] = t[67] & t[45];
  assign t[37] = t[73] ^ t[74];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[74]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[68] ^ t[39]);
  assign t[41] = t[68] & t[47];
  assign t[42] = t[66] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[67] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[68] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[70] ^ t[75];
  assign t[49] = t[66] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[72] ^ t[76];
  assign t[51] = t[67] ^ t[32];
  assign t[52] = t[74] ^ t[77];
  assign t[53] = t[68] ^ t[37];
  assign t[54] = x[0] ? x[42] : t[55];
  assign t[55] = ~(t[56] ^ t[57]);
  assign t[56] = ~(t[58] ^ t[78]);
  assign t[57] = ~(t[59] ^ t[60]);
  assign t[58] = ~t[61];
  assign t[59] = ~(t[62]);
  assign t[5] = ~(t[8]);
  assign t[60] = ~(t[63]);
  assign t[61] = ~(t[64]);
  assign t[62] = t[52] ^ t[24];
  assign t[63] = t[48] ^ t[16];
  assign t[64] = t[50] ^ t[20];
  assign t[65] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[66] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[67] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[68] = (t[85] & ~t[86]) | (~t[85] & t[86]);
  assign t[69] = (t[81] & ~t[87]) | (~t[81] & t[87]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[81] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[87]) | (~t[81] & ~t[89] & t[90]) | (t[88] & t[89] & t[87]);
  assign t[71] = (t[83] & ~t[91]) | (~t[83] & t[91]);
  assign t[72] = (t[83] & ~t[93] & ~t[94]) | (~t[92] & t[93] & ~t[91]) | (~t[83] & ~t[93] & t[94]) | (t[92] & t[93] & t[91]);
  assign t[73] = (t[85] & ~t[95]) | (~t[85] & t[95]);
  assign t[74] = (t[85] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[95]) | (~t[85] & ~t[97] & t[98]) | (t[96] & t[97] & t[95]);
  assign t[75] = (t[81] & ~t[89] & ~t[87]) | (~t[88] & t[89] & ~t[90]) | (~t[81] & ~t[89] & t[87]) | (t[88] & t[89] & t[90]);
  assign t[76] = (t[83] & ~t[93] & ~t[91]) | (~t[92] & t[93] & ~t[94]) | (~t[83] & ~t[93] & t[91]) | (t[92] & t[93] & t[94]);
  assign t[77] = (t[85] & ~t[97] & ~t[95]) | (~t[96] & t[97] & ~t[98]) | (~t[85] & ~t[97] & t[95]) | (t[96] & t[97] & t[98]);
  assign t[78] = (t[79] & ~t[100] & ~t[102]) | (~t[99] & t[100] & ~t[101]) | (~t[79] & ~t[100] & t[102]) | (t[99] & t[100] & t[101]);
  assign t[79] = t[103] ^ x[7];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = t[104] ^ x[8];
  assign t[81] = t[105] ^ x[14];
  assign t[82] = t[106] ^ x[15];
  assign t[83] = t[107] ^ x[21];
  assign t[84] = t[108] ^ x[22];
  assign t[85] = t[109] ^ x[28];
  assign t[86] = t[110] ^ x[29];
  assign t[87] = t[111] ^ x[30];
  assign t[88] = t[112] ^ x[31];
  assign t[89] = t[113] ^ x[32];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = t[114] ^ x[33];
  assign t[91] = t[115] ^ x[34];
  assign t[92] = t[116] ^ x[35];
  assign t[93] = t[117] ^ x[36];
  assign t[94] = t[118] ^ x[37];
  assign t[95] = t[119] ^ x[38];
  assign t[96] = t[120] ^ x[39];
  assign t[97] = t[121] ^ x[40];
  assign t[98] = t[122] ^ x[41];
  assign t[99] = t[123] ^ x[43];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0] & ~t[54]) | (~t[0] & t[54]);
endmodule

module R2ind152(x, y);
 input [46:0] x;
 output y;

 wire [179:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[101] = (t[124] & t[125] & ~t[126] & t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[126] & ~t[127] & t[128] & ~t[129] & t[130]) | (~t[125] & t[126] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[125] & t[126] & ~t[129] & ~t[130]) | (~t[124] & t[126] & t[127] & ~t[128] & t[129]) | (t[126] & ~t[127] & t[129] & ~t[130]);
  assign t[102] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[103] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[104] = (t[138] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[139] & ~t[140] & ~t[143] & ~t[144]) | (~t[138] & t[139] & t[140] & t[141] & ~t[144]) | (~t[138] & t[139] & t[142] & t[143] & ~t[144]) | (t[138] & ~t[140] & ~t[142] & t[144]) | (~t[138] & t[140] & t[142] & t[144]);
  assign t[105] = (t[138] & t[139] & ~t[140] & t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[140] & ~t[141] & t[142] & ~t[143] & t[144]) | (~t[139] & t[140] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[139] & t[140] & ~t[143] & ~t[144]) | (~t[138] & t[140] & t[141] & ~t[142] & t[143]) | (t[140] & ~t[141] & t[143] & ~t[144]);
  assign t[106] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[107] = (t[145] & t[146] & ~t[147] & t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[147] & ~t[148] & t[149] & ~t[150] & t[151]) | (~t[146] & t[147] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[146] & t[147] & ~t[150] & ~t[151]) | (~t[145] & t[147] & t[148] & ~t[149] & t[150]) | (t[147] & ~t[148] & t[150] & ~t[151]);
  assign t[108] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[109] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[10] = t[17] ^ t[18];
  assign t[110] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[111] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[112] = (t[138] & t[139] & ~t[140] & ~t[142] & t[143] & ~t[144]) | (t[138] & t[140] & ~t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & t[142] & ~t[143] & ~t[144]) | (~t[138] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[138] & ~t[139] & ~t[141] & t[142] & ~t[144]) | (~t[138] & ~t[140] & t[141] & t[142] & t[143]) | (t[141] & t[142] & ~t[143] & ~t[144]);
  assign t[113] = (t[139] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & t[139] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[139] & ~t[140] & ~t[143] & ~t[144]) | (t[138] & ~t[139] & t[140] & t[141] & ~t[144]) | (t[138] & ~t[139] & t[142] & t[143] & ~t[144]) | (t[139] & ~t[141] & ~t[143] & t[144]) | (~t[139] & t[141] & t[143] & t[144]);
  assign t[114] = (t[138] & t[139] & t[140] & ~t[141] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & ~t[141] & ~t[142] & t[143] & t[144]) | (~t[139] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[140] & t[141] & ~t[143] & ~t[144]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[144]) | (~t[139] & t[140] & t[141] & t[142] & ~t[143]) | (~t[140] & t[141] & t[142] & ~t[144]);
  assign t[115] = (t[138] & t[139] & ~t[141] & t[142] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[141] & ~t[142] & t[143] & ~t[144]) | (~t[138] & ~t[139] & ~t[140] & t[143] & ~t[144]) | (~t[139] & t[140] & ~t[141] & t[142] & t[143]) | (t[140] & ~t[142] & t[143] & ~t[144]);
  assign t[116] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[117] = (t[146] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & t[146] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[146] & ~t[147] & ~t[150] & ~t[151]) | (t[145] & ~t[146] & t[147] & t[148] & ~t[151]) | (t[145] & ~t[146] & t[149] & t[150] & ~t[151]) | (t[146] & ~t[148] & ~t[150] & t[151]) | (~t[146] & t[148] & t[150] & t[151]);
  assign t[118] = (t[145] & t[146] & t[147] & ~t[148] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & ~t[148] & ~t[149] & t[150] & t[151]) | (~t[146] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[147] & t[148] & ~t[150] & ~t[151]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[151]) | (~t[146] & t[147] & t[148] & t[149] & ~t[150]) | (~t[147] & t[148] & t[149] & ~t[151]);
  assign t[119] = (t[145] & t[146] & ~t[148] & t[149] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[148] & ~t[149] & t[150] & ~t[151]) | (~t[145] & ~t[146] & ~t[147] & t[150] & ~t[151]) | (~t[146] & t[147] & ~t[148] & t[149] & t[150]) | (t[147] & ~t[149] & t[150] & ~t[151]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[121] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[122] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[123] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[124] = t[152] ^ x[7];
  assign t[125] = t[153] ^ x[43];
  assign t[126] = t[154] ^ x[8];
  assign t[127] = t[155] ^ x[44];
  assign t[128] = t[156] ^ x[45];
  assign t[129] = t[157] ^ x[46];
  assign t[12] = t[21] ^ t[22];
  assign t[130] = t[158] ^ x[6];
  assign t[131] = t[159] ^ x[14];
  assign t[132] = t[160] ^ x[31];
  assign t[133] = t[161] ^ x[15];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = t[163] ^ x[30];
  assign t[136] = t[164] ^ x[33];
  assign t[137] = t[165] ^ x[13];
  assign t[138] = t[166] ^ x[21];
  assign t[139] = t[167] ^ x[35];
  assign t[13] = t[23] ^ t[24];
  assign t[140] = t[168] ^ x[22];
  assign t[141] = t[169] ^ x[36];
  assign t[142] = t[170] ^ x[34];
  assign t[143] = t[171] ^ x[37];
  assign t[144] = t[172] ^ x[20];
  assign t[145] = t[173] ^ x[28];
  assign t[146] = t[174] ^ x[39];
  assign t[147] = t[175] ^ x[29];
  assign t[148] = t[176] ^ x[40];
  assign t[149] = t[177] ^ x[38];
  assign t[14] = t[25] ^ t[26];
  assign t[150] = t[178] ^ x[41];
  assign t[151] = t[179] ^ x[27];
  assign t[152] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[153] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[154] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[155] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[156] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[157] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[158] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[159] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[15] = t[27] ^ t[28];
  assign t[160] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[161] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[162] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[163] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[164] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[165] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[166] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[167] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[168] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[169] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[16] = t[29] & t[30];
  assign t[170] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[171] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[172] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[173] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[174] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[175] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[176] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[177] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[178] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[179] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[17] = t[31] ^ t[16];
  assign t[18] = t[63] ^ t[29];
  assign t[19] = t[32] ^ t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] & t[35];
  assign t[21] = t[36] ^ t[20];
  assign t[22] = t[64] ^ t[34];
  assign t[23] = t[37] ^ t[38];
  assign t[24] = t[39] & t[40];
  assign t[25] = t[41] ^ t[24];
  assign t[26] = t[65] ^ t[39];
  assign t[27] = t[66] ^ t[67];
  assign t[28] = t[29] & t[42];
  assign t[29] = ~(t[67]);
  assign t[2] = ~(t[4] ^ t[62]);
  assign t[30] = ~(t[63] ^ t[29]);
  assign t[31] = t[63] & t[43];
  assign t[32] = t[68] ^ t[69];
  assign t[33] = t[34] & t[44];
  assign t[34] = ~(t[69]);
  assign t[35] = ~(t[64] ^ t[34]);
  assign t[36] = t[64] & t[45];
  assign t[37] = t[70] ^ t[71];
  assign t[38] = t[39] & t[46];
  assign t[39] = ~(t[71]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[65] ^ t[39]);
  assign t[41] = t[65] & t[47];
  assign t[42] = t[63] ^ t[48];
  assign t[43] = t[49] ^ t[28];
  assign t[44] = t[64] ^ t[50];
  assign t[45] = t[51] ^ t[33];
  assign t[46] = t[65] ^ t[52];
  assign t[47] = t[53] ^ t[38];
  assign t[48] = t[67] ^ t[72];
  assign t[49] = t[63] ^ t[27];
  assign t[4] = ~t[7];
  assign t[50] = t[69] ^ t[73];
  assign t[51] = t[64] ^ t[32];
  assign t[52] = t[71] ^ t[74];
  assign t[53] = t[65] ^ t[37];
  assign t[54] = x[0] ? x[42] : t[55];
  assign t[55] = ~(t[56] ^ t[57]);
  assign t[56] = ~(t[58] ^ t[75]);
  assign t[57] = ~(t[59] ^ t[60]);
  assign t[58] = ~t[61];
  assign t[59] = ~(t[13]);
  assign t[5] = ~(t[8]);
  assign t[60] = ~(t[9]);
  assign t[61] = ~(t[11]);
  assign t[62] = (t[76] & ~t[77]) | (~t[76] & t[77]);
  assign t[63] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[64] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[65] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[66] = (t[78] & ~t[84]) | (~t[78] & t[84]);
  assign t[67] = (t[78] & ~t[86] & ~t[87]) | (~t[85] & t[86] & ~t[84]) | (~t[78] & ~t[86] & t[87]) | (t[85] & t[86] & t[84]);
  assign t[68] = (t[80] & ~t[88]) | (~t[80] & t[88]);
  assign t[69] = (t[80] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[88]) | (~t[80] & ~t[90] & t[91]) | (t[89] & t[90] & t[88]);
  assign t[6] = ~(t[9] ^ t[10]);
  assign t[70] = (t[82] & ~t[92]) | (~t[82] & t[92]);
  assign t[71] = (t[82] & ~t[94] & ~t[95]) | (~t[93] & t[94] & ~t[92]) | (~t[82] & ~t[94] & t[95]) | (t[93] & t[94] & t[92]);
  assign t[72] = (t[78] & ~t[86] & ~t[84]) | (~t[85] & t[86] & ~t[87]) | (~t[78] & ~t[86] & t[84]) | (t[85] & t[86] & t[87]);
  assign t[73] = (t[80] & ~t[90] & ~t[88]) | (~t[89] & t[90] & ~t[91]) | (~t[80] & ~t[90] & t[88]) | (t[89] & t[90] & t[91]);
  assign t[74] = (t[82] & ~t[94] & ~t[92]) | (~t[93] & t[94] & ~t[95]) | (~t[82] & ~t[94] & t[92]) | (t[93] & t[94] & t[95]);
  assign t[75] = (t[76] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[99]) | (~t[76] & ~t[97] & t[98]) | (t[96] & t[97] & t[99]);
  assign t[76] = t[100] ^ x[7];
  assign t[77] = t[101] ^ x[8];
  assign t[78] = t[102] ^ x[14];
  assign t[79] = t[103] ^ x[15];
  assign t[7] = ~(t[11] ^ t[12]);
  assign t[80] = t[104] ^ x[21];
  assign t[81] = t[105] ^ x[22];
  assign t[82] = t[106] ^ x[28];
  assign t[83] = t[107] ^ x[29];
  assign t[84] = t[108] ^ x[30];
  assign t[85] = t[109] ^ x[31];
  assign t[86] = t[110] ^ x[32];
  assign t[87] = t[111] ^ x[33];
  assign t[88] = t[112] ^ x[34];
  assign t[89] = t[113] ^ x[35];
  assign t[8] = ~(t[13] ^ t[14]);
  assign t[90] = t[114] ^ x[36];
  assign t[91] = t[115] ^ x[37];
  assign t[92] = t[116] ^ x[38];
  assign t[93] = t[117] ^ x[39];
  assign t[94] = t[118] ^ x[40];
  assign t[95] = t[119] ^ x[41];
  assign t[96] = t[120] ^ x[43];
  assign t[97] = t[121] ^ x[44];
  assign t[98] = t[122] ^ x[45];
  assign t[99] = t[123] ^ x[46];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0] & ~t[54]) | (~t[0] & t[54]);
endmodule

module R2ind153(x, y);
 input [46:0] x;
 output y;

 wire [161:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[101] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[102] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[103] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[104] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[105] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[106] = t[134] ^ x[8];
  assign t[107] = t[135] ^ x[9];
  assign t[108] = t[136] ^ x[6];
  assign t[109] = t[137] ^ x[10];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[138] ^ x[11];
  assign t[111] = t[139] ^ x[12];
  assign t[112] = t[140] ^ x[7];
  assign t[113] = t[141] ^ x[18];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[43];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[17];
  assign t[11] = t[47] ^ t[48];
  assign t[120] = t[148] ^ x[28];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[44];
  assign t[123] = t[151] ^ x[30];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[27];
  assign t[127] = t[155] ^ x[38];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[45];
  assign t[12] = t[17] & t[18];
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[37];
  assign t[134] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[135] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[136] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[137] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[138] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[139] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[13] = t[49] ^ t[50];
  assign t[140] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[141] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[142] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[143] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[144] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[145] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[146] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[147] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[148] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[149] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[14] = t[19] & t[20];
  assign t[150] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[151] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[152] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[153] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[154] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[155] = (x[33] & ~x[34] & ~x[35]) | (~x[33] & x[34] & ~x[35]) | (~x[33] & ~x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[156] = (x[33] & ~x[34] & ~x[36]) | (~x[33] & x[34] & ~x[36]) | (~x[33] & ~x[34] & x[36]) | (x[33] & x[34] & x[36]);
  assign t[157] = (x[33] & ~x[35]) | (~x[33] & x[35]);
  assign t[158] = (x[33] & ~x[36]) | (~x[33] & x[36]);
  assign t[159] = (x[34] & ~x[35]) | (~x[34] & x[35]);
  assign t[15] = t[51] ^ t[52];
  assign t[160] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[161] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[47]);
  assign t[18] = ~(t[53] ^ t[17]);
  assign t[19] = ~(t[49]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[54] ^ t[19]);
  assign t[21] = ~(t[51]);
  assign t[22] = ~(t[55] ^ t[21]);
  assign t[23] = x[0] ? x[46] : t[24];
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~(t[27] ^ t[56]);
  assign t[26] = ~(t[28] ^ t[29]);
  assign t[27] = ~t[30];
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[4] ^ t[46]);
  assign t[30] = ~(t[33]);
  assign t[31] = t[34] ^ t[12];
  assign t[32] = t[35] ^ t[14];
  assign t[33] = t[36] ^ t[16];
  assign t[34] = t[37] ^ t[38];
  assign t[35] = t[39] ^ t[40];
  assign t[36] = t[41] ^ t[42];
  assign t[37] = t[57] ^ t[47];
  assign t[38] = t[17] & t[43];
  assign t[39] = t[58] ^ t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[19] & t[44];
  assign t[41] = t[59] ^ t[51];
  assign t[42] = t[21] & t[45];
  assign t[43] = t[53] ^ t[11];
  assign t[44] = t[54] ^ t[13];
  assign t[45] = t[55] ^ t[15];
  assign t[46] = (t[60] & ~t[62] & ~t[64]) | (~t[61] & t[62] & ~t[63]) | (~t[60] & ~t[62] & t[64]) | (t[61] & t[62] & t[63]);
  assign t[47] = (t[65] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[65] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[48] = (t[65] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[65] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[49] = (t[70] & ~t[72] & ~t[74]) | (~t[71] & t[72] & ~t[73]) | (~t[70] & ~t[72] & t[74]) | (t[71] & t[72] & t[73]);
  assign t[4] = ~t[7];
  assign t[50] = (t[70] & ~t[72] & ~t[73]) | (~t[71] & t[72] & ~t[74]) | (~t[70] & ~t[72] & t[73]) | (t[71] & t[72] & t[74]);
  assign t[51] = (t[75] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[75] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[52] = (t[75] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[75] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[53] = (t[65] & ~t[80]) | (~t[65] & t[80]);
  assign t[54] = (t[70] & ~t[81]) | (~t[70] & t[81]);
  assign t[55] = (t[75] & ~t[82]) | (~t[75] & t[82]);
  assign t[56] = (t[60] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[64]) | (~t[60] & ~t[62] & t[63]) | (t[61] & t[62] & t[64]);
  assign t[57] = (t[65] & ~t[68]) | (~t[65] & t[68]);
  assign t[58] = (t[70] & ~t[73]) | (~t[70] & t[73]);
  assign t[59] = (t[75] & ~t[78]) | (~t[75] & t[78]);
  assign t[5] = ~(t[8]);
  assign t[60] = t[83] ^ x[8];
  assign t[61] = t[84] ^ x[9];
  assign t[62] = t[85] ^ x[10];
  assign t[63] = t[86] ^ x[11];
  assign t[64] = t[87] ^ x[12];
  assign t[65] = t[88] ^ x[18];
  assign t[66] = t[89] ^ x[19];
  assign t[67] = t[90] ^ x[20];
  assign t[68] = t[91] ^ x[21];
  assign t[69] = t[92] ^ x[22];
  assign t[6] = ~(t[9]);
  assign t[70] = t[93] ^ x[28];
  assign t[71] = t[94] ^ x[29];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[31];
  assign t[74] = t[97] ^ x[32];
  assign t[75] = t[98] ^ x[38];
  assign t[76] = t[99] ^ x[39];
  assign t[77] = t[100] ^ x[40];
  assign t[78] = t[101] ^ x[41];
  assign t[79] = t[102] ^ x[42];
  assign t[7] = ~(t[10]);
  assign t[80] = t[103] ^ x[43];
  assign t[81] = t[104] ^ x[44];
  assign t[82] = t[105] ^ x[45];
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[85] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[86] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[89] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[92] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[93] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[94] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[95] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[97] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[98] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[99] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0] & ~t[23]) | (~t[0] & t[23]);
endmodule

module R2ind154(x, y);
 input [47:0] x;
 output y;

 wire [202:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[8];
  assign t[101] = t[125] ^ x[14];
  assign t[102] = t[126] ^ x[15];
  assign t[103] = t[127] ^ x[21];
  assign t[104] = t[128] ^ x[22];
  assign t[105] = t[129] ^ x[28];
  assign t[106] = t[130] ^ x[29];
  assign t[107] = t[131] ^ x[30];
  assign t[108] = t[132] ^ x[31];
  assign t[109] = t[133] ^ x[32];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[134] ^ x[33];
  assign t[111] = t[135] ^ x[34];
  assign t[112] = t[136] ^ x[35];
  assign t[113] = t[137] ^ x[36];
  assign t[114] = t[138] ^ x[37];
  assign t[115] = t[139] ^ x[38];
  assign t[116] = t[140] ^ x[39];
  assign t[117] = t[141] ^ x[40];
  assign t[118] = t[142] ^ x[41];
  assign t[119] = t[143] ^ x[43];
  assign t[11] = t[20] & t[21];
  assign t[120] = t[144] ^ x[45];
  assign t[121] = t[145] ^ x[46];
  assign t[122] = t[146] ^ x[47];
  assign t[123] = (t[147] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (t[147] & ~t[148] & ~t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[148] & ~t[149] & ~t[152] & ~t[153]) | (~t[147] & t[148] & t[149] & t[150] & ~t[153]) | (~t[147] & t[148] & t[151] & t[152] & ~t[153]) | (t[147] & ~t[149] & ~t[151] & t[153]) | (~t[147] & t[149] & t[151] & t[153]);
  assign t[124] = (t[147] & t[148] & ~t[149] & ~t[151] & t[152] & ~t[153]) | (t[147] & t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[153]) | (~t[147] & ~t[149] & ~t[150] & t[151] & ~t[152]) | (~t[147] & ~t[148] & ~t[150] & t[151] & ~t[153]) | (~t[147] & ~t[149] & t[150] & t[151] & t[152]) | (t[150] & t[151] & ~t[152] & ~t[153]);
  assign t[125] = (t[154] & ~t[156] & ~t[157] & ~t[158] & ~t[159]) | (t[154] & ~t[155] & ~t[157] & ~t[158] & ~t[160]) | (t[154] & ~t[155] & ~t[156] & ~t[159] & ~t[160]) | (~t[154] & t[155] & t[156] & t[157] & ~t[160]) | (~t[154] & t[155] & t[158] & t[159] & ~t[160]) | (t[154] & ~t[156] & ~t[158] & t[160]) | (~t[154] & t[156] & t[158] & t[160]);
  assign t[126] = (t[154] & t[155] & ~t[156] & t[157] & ~t[158] & ~t[160]) | (t[154] & ~t[156] & ~t[157] & t[158] & ~t[159] & t[160]) | (~t[155] & t[156] & ~t[157] & ~t[158] & ~t[160]) | (~t[154] & t[156] & ~t[157] & ~t[158] & ~t[159]) | (~t[154] & ~t[155] & t[156] & ~t[159] & ~t[160]) | (~t[154] & t[156] & t[157] & ~t[158] & t[159]) | (t[156] & ~t[157] & t[159] & ~t[160]);
  assign t[127] = (t[161] & ~t[163] & ~t[164] & ~t[165] & ~t[166]) | (t[161] & ~t[162] & ~t[164] & ~t[165] & ~t[167]) | (t[161] & ~t[162] & ~t[163] & ~t[166] & ~t[167]) | (~t[161] & t[162] & t[163] & t[164] & ~t[167]) | (~t[161] & t[162] & t[165] & t[166] & ~t[167]) | (t[161] & ~t[163] & ~t[165] & t[167]) | (~t[161] & t[163] & t[165] & t[167]);
  assign t[128] = (t[161] & t[162] & ~t[163] & t[164] & ~t[165] & ~t[167]) | (t[161] & ~t[163] & ~t[164] & t[165] & ~t[166] & t[167]) | (~t[162] & t[163] & ~t[164] & ~t[165] & ~t[167]) | (~t[161] & t[163] & ~t[164] & ~t[165] & ~t[166]) | (~t[161] & ~t[162] & t[163] & ~t[166] & ~t[167]) | (~t[161] & t[163] & t[164] & ~t[165] & t[166]) | (t[163] & ~t[164] & t[166] & ~t[167]);
  assign t[129] = (t[168] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (t[168] & ~t[169] & ~t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[169] & ~t[170] & ~t[173] & ~t[174]) | (~t[168] & t[169] & t[170] & t[171] & ~t[174]) | (~t[168] & t[169] & t[172] & t[173] & ~t[174]) | (t[168] & ~t[170] & ~t[172] & t[174]) | (~t[168] & t[170] & t[172] & t[174]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (t[168] & t[169] & ~t[170] & t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[170] & ~t[171] & t[172] & ~t[173] & t[174]) | (~t[169] & t[170] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[169] & t[170] & ~t[173] & ~t[174]) | (~t[168] & t[170] & t[171] & ~t[172] & t[173]) | (t[170] & ~t[171] & t[173] & ~t[174]);
  assign t[131] = (t[155] & ~t[156] & ~t[157] & ~t[158] & ~t[159]) | (~t[154] & t[155] & ~t[157] & ~t[158] & ~t[160]) | (~t[154] & t[155] & ~t[156] & ~t[159] & ~t[160]) | (t[154] & ~t[155] & t[156] & t[157] & ~t[160]) | (t[154] & ~t[155] & t[158] & t[159] & ~t[160]) | (t[155] & ~t[157] & ~t[159] & t[160]) | (~t[155] & t[157] & t[159] & t[160]);
  assign t[132] = (t[154] & t[155] & t[156] & ~t[157] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[157] & ~t[158] & t[159] & t[160]) | (~t[155] & ~t[156] & t[157] & ~t[158] & ~t[159]) | (~t[154] & ~t[156] & t[157] & ~t[159] & ~t[160]) | (~t[154] & ~t[155] & t[157] & ~t[158] & ~t[160]) | (~t[155] & t[156] & t[157] & t[158] & ~t[159]) | (~t[156] & t[157] & t[158] & ~t[160]);
  assign t[133] = (t[154] & t[155] & ~t[156] & ~t[158] & t[159] & ~t[160]) | (t[154] & t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[160]) | (~t[154] & ~t[156] & ~t[157] & t[158] & ~t[159]) | (~t[154] & ~t[155] & ~t[157] & t[158] & ~t[160]) | (~t[154] & ~t[156] & t[157] & t[158] & t[159]) | (t[157] & t[158] & ~t[159] & ~t[160]);
  assign t[134] = (t[154] & t[155] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[156] & ~t[157] & ~t[158] & t[159]) | (~t[154] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[154] & ~t[155] & ~t[156] & t[159] & ~t[160]) | (~t[155] & t[156] & ~t[157] & t[158] & t[159]) | (t[156] & ~t[158] & t[159] & ~t[160]);
  assign t[135] = (t[162] & ~t[163] & ~t[164] & ~t[165] & ~t[166]) | (~t[161] & t[162] & ~t[164] & ~t[165] & ~t[167]) | (~t[161] & t[162] & ~t[163] & ~t[166] & ~t[167]) | (t[161] & ~t[162] & t[163] & t[164] & ~t[167]) | (t[161] & ~t[162] & t[165] & t[166] & ~t[167]) | (t[162] & ~t[164] & ~t[166] & t[167]) | (~t[162] & t[164] & t[166] & t[167]);
  assign t[136] = (t[161] & t[162] & t[163] & ~t[164] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & ~t[164] & ~t[165] & t[166] & t[167]) | (~t[162] & ~t[163] & t[164] & ~t[165] & ~t[166]) | (~t[161] & ~t[163] & t[164] & ~t[166] & ~t[167]) | (~t[161] & ~t[162] & t[164] & ~t[165] & ~t[167]) | (~t[162] & t[163] & t[164] & t[165] & ~t[166]) | (~t[163] & t[164] & t[165] & ~t[167]);
  assign t[137] = (t[161] & t[162] & ~t[163] & ~t[165] & t[166] & ~t[167]) | (t[161] & t[163] & ~t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[163] & t[165] & ~t[166] & ~t[167]) | (~t[161] & ~t[163] & ~t[164] & t[165] & ~t[166]) | (~t[161] & ~t[162] & ~t[164] & t[165] & ~t[167]) | (~t[161] & ~t[163] & t[164] & t[165] & t[166]) | (t[164] & t[165] & ~t[166] & ~t[167]);
  assign t[138] = (t[161] & t[162] & ~t[164] & t[165] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[163] & ~t[164] & ~t[165] & t[166]) | (~t[161] & ~t[164] & ~t[165] & t[166] & ~t[167]) | (~t[161] & ~t[162] & ~t[163] & t[166] & ~t[167]) | (~t[162] & t[163] & ~t[164] & t[165] & t[166]) | (t[163] & ~t[165] & t[166] & ~t[167]);
  assign t[139] = (t[169] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & t[169] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[169] & ~t[170] & ~t[173] & ~t[174]) | (t[168] & ~t[169] & t[170] & t[171] & ~t[174]) | (t[168] & ~t[169] & t[172] & t[173] & ~t[174]) | (t[169] & ~t[171] & ~t[173] & t[174]) | (~t[169] & t[171] & t[173] & t[174]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (t[168] & t[169] & t[170] & ~t[171] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & ~t[171] & ~t[172] & t[173] & t[174]) | (~t[169] & ~t[170] & t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[170] & t[171] & ~t[173] & ~t[174]) | (~t[168] & ~t[169] & t[171] & ~t[172] & ~t[174]) | (~t[169] & t[170] & t[171] & t[172] & ~t[173]) | (~t[170] & t[171] & t[172] & ~t[174]);
  assign t[141] = (t[168] & t[169] & ~t[170] & ~t[172] & t[173] & ~t[174]) | (t[168] & t[170] & ~t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & t[172] & ~t[173] & ~t[174]) | (~t[168] & ~t[170] & ~t[171] & t[172] & ~t[173]) | (~t[168] & ~t[169] & ~t[171] & t[172] & ~t[174]) | (~t[168] & ~t[170] & t[171] & t[172] & t[173]) | (t[171] & t[172] & ~t[173] & ~t[174]);
  assign t[142] = (t[168] & t[169] & ~t[171] & t[172] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & ~t[171] & ~t[172] & t[173]) | (~t[168] & ~t[171] & ~t[172] & t[173] & ~t[174]) | (~t[168] & ~t[169] & ~t[170] & t[173] & ~t[174]) | (~t[169] & t[170] & ~t[171] & t[172] & t[173]) | (t[170] & ~t[172] & t[173] & ~t[174]);
  assign t[143] = (t[147] & t[148] & ~t[149] & t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[149] & ~t[150] & t[151] & ~t[152] & t[153]) | (~t[148] & t[149] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[148] & t[149] & ~t[152] & ~t[153]) | (~t[147] & t[149] & t[150] & ~t[151] & t[152]) | (t[149] & ~t[150] & t[152] & ~t[153]);
  assign t[144] = (t[148] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & t[148] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[148] & ~t[149] & ~t[152] & ~t[153]) | (t[147] & ~t[148] & t[149] & t[150] & ~t[153]) | (t[147] & ~t[148] & t[151] & t[152] & ~t[153]) | (t[148] & ~t[150] & ~t[152] & t[153]) | (~t[148] & t[150] & t[152] & t[153]);
  assign t[145] = (t[147] & t[148] & t[149] & ~t[150] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[150] & ~t[151] & t[152] & t[153]) | (~t[148] & ~t[149] & t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[149] & t[150] & ~t[152] & ~t[153]) | (~t[147] & ~t[148] & t[150] & ~t[151] & ~t[153]) | (~t[148] & t[149] & t[150] & t[151] & ~t[152]) | (~t[149] & t[150] & t[151] & ~t[153]);
  assign t[146] = (t[147] & t[148] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & ~t[150] & ~t[151] & t[152]) | (~t[147] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[147] & ~t[148] & ~t[149] & t[152] & ~t[153]) | (~t[148] & t[149] & ~t[150] & t[151] & t[152]) | (t[149] & ~t[151] & t[152] & ~t[153]);
  assign t[147] = t[175] ^ x[7];
  assign t[148] = t[176] ^ x[45];
  assign t[149] = t[177] ^ x[43];
  assign t[14] = t[85] & t[26];
  assign t[150] = t[178] ^ x[46];
  assign t[151] = t[179] ^ x[8];
  assign t[152] = t[180] ^ x[47];
  assign t[153] = t[181] ^ x[6];
  assign t[154] = t[182] ^ x[14];
  assign t[155] = t[183] ^ x[30];
  assign t[156] = t[184] ^ x[15];
  assign t[157] = t[185] ^ x[31];
  assign t[158] = t[186] ^ x[32];
  assign t[159] = t[187] ^ x[33];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[188] ^ x[13];
  assign t[161] = t[189] ^ x[21];
  assign t[162] = t[190] ^ x[34];
  assign t[163] = t[191] ^ x[22];
  assign t[164] = t[192] ^ x[35];
  assign t[165] = t[193] ^ x[36];
  assign t[166] = t[194] ^ x[37];
  assign t[167] = t[195] ^ x[20];
  assign t[168] = t[196] ^ x[28];
  assign t[169] = t[197] ^ x[38];
  assign t[16] = t[29] ^ t[27];
  assign t[170] = t[198] ^ x[29];
  assign t[171] = t[199] ^ x[39];
  assign t[172] = t[200] ^ x[40];
  assign t[173] = t[201] ^ x[41];
  assign t[174] = t[202] ^ x[27];
  assign t[175] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[176] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[177] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[178] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[179] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[181] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[182] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[183] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[184] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[185] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[186] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[187] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[188] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[189] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[18] = t[86] & t[31];
  assign t[190] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[191] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[192] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[193] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[194] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[195] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[196] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[197] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[198] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[199] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[201] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[202] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[87] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[88]);
  assign t[28] = ~(t[85] ^ t[27]);
  assign t[29] = t[89] ^ t[88];
  assign t[2] = ~(t[4] ^ t[84]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[90]);
  assign t[33] = ~(t[86] ^ t[32]);
  assign t[34] = t[91] ^ t[90];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[92]);
  assign t[38] = ~(t[87] ^ t[37]);
  assign t[39] = t[93] ^ t[92];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[85] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[85] ^ t[50];
  assign t[44] = t[86] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[86] ^ t[51];
  assign t[47] = t[87] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[87] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[88] ^ t[94];
  assign t[51] = t[90] ^ t[95];
  assign t[52] = t[92] ^ t[96];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[97]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61] ^ t[62]);
  assign t[59] = ~(t[63] ^ t[64]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[65] ^ t[66]);
  assign t[61] = t[67] ^ t[15];
  assign t[62] = t[8] ^ t[68];
  assign t[63] = t[69] ^ t[19];
  assign t[64] = t[10] ^ t[70];
  assign t[65] = t[71] ^ t[23];
  assign t[66] = t[12] ^ t[72];
  assign t[67] = t[29] ^ t[42];
  assign t[68] = t[85] ^ t[27];
  assign t[69] = t[34] ^ t[45];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[86] ^ t[32];
  assign t[71] = t[39] ^ t[48];
  assign t[72] = t[87] ^ t[37];
  assign t[73] = x[0] ? x[44] : t[74];
  assign t[74] = ~(t[75] ^ t[76]);
  assign t[75] = ~(t[77] ^ t[98]);
  assign t[76] = ~(t[78] ^ t[79]);
  assign t[77] = ~t[80];
  assign t[78] = ~(t[81]);
  assign t[79] = ~(t[82]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[83]);
  assign t[81] = t[50] ^ t[15];
  assign t[82] = t[51] ^ t[19];
  assign t[83] = t[52] ^ t[23];
  assign t[84] = (t[99] & ~t[100]) | (~t[99] & t[100]);
  assign t[85] = (t[101] & ~t[102]) | (~t[101] & t[102]);
  assign t[86] = (t[103] & ~t[104]) | (~t[103] & t[104]);
  assign t[87] = (t[105] & ~t[106]) | (~t[105] & t[106]);
  assign t[88] = (t[101] & ~t[108] & ~t[110]) | (~t[107] & t[108] & ~t[109]) | (~t[101] & ~t[108] & t[110]) | (t[107] & t[108] & t[109]);
  assign t[89] = (t[101] & ~t[109]) | (~t[101] & t[109]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (t[103] & ~t[112] & ~t[114]) | (~t[111] & t[112] & ~t[113]) | (~t[103] & ~t[112] & t[114]) | (t[111] & t[112] & t[113]);
  assign t[91] = (t[103] & ~t[113]) | (~t[103] & t[113]);
  assign t[92] = (t[105] & ~t[116] & ~t[118]) | (~t[115] & t[116] & ~t[117]) | (~t[105] & ~t[116] & t[118]) | (t[115] & t[116] & t[117]);
  assign t[93] = (t[105] & ~t[117]) | (~t[105] & t[117]);
  assign t[94] = (t[101] & ~t[108] & ~t[109]) | (~t[107] & t[108] & ~t[110]) | (~t[101] & ~t[108] & t[109]) | (t[107] & t[108] & t[110]);
  assign t[95] = (t[103] & ~t[112] & ~t[113]) | (~t[111] & t[112] & ~t[114]) | (~t[103] & ~t[112] & t[113]) | (t[111] & t[112] & t[114]);
  assign t[96] = (t[105] & ~t[116] & ~t[117]) | (~t[115] & t[116] & ~t[118]) | (~t[105] & ~t[116] & t[117]) | (t[115] & t[116] & t[118]);
  assign t[97] = (t[99] & ~t[119]) | (~t[99] & t[119]);
  assign t[98] = (t[99] & ~t[121] & ~t[122]) | (~t[120] & t[121] & ~t[100]) | (~t[99] & ~t[121] & t[122]) | (t[120] & t[121] & t[100]);
  assign t[99] = t[123] ^ x[7];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[73]) | (~t[0] & t[53] & ~t[73]) | (~t[0] & ~t[53] & t[73]) | (t[0] & t[53] & t[73]);
endmodule

module R2ind155(x, y);
 input [47:0] x;
 output y;

 wire [199:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[21];
  assign t[101] = t[125] ^ x[22];
  assign t[102] = t[126] ^ x[28];
  assign t[103] = t[127] ^ x[29];
  assign t[104] = t[128] ^ x[30];
  assign t[105] = t[129] ^ x[31];
  assign t[106] = t[130] ^ x[32];
  assign t[107] = t[131] ^ x[33];
  assign t[108] = t[132] ^ x[34];
  assign t[109] = t[133] ^ x[35];
  assign t[10] = t[18] ^ t[19];
  assign t[110] = t[134] ^ x[36];
  assign t[111] = t[135] ^ x[37];
  assign t[112] = t[136] ^ x[38];
  assign t[113] = t[137] ^ x[39];
  assign t[114] = t[138] ^ x[40];
  assign t[115] = t[139] ^ x[41];
  assign t[116] = t[140] ^ x[43];
  assign t[117] = t[141] ^ x[45];
  assign t[118] = t[142] ^ x[46];
  assign t[119] = t[143] ^ x[47];
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[121] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[122] = (t[151] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & ~t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[152] & ~t[153] & ~t[156] & ~t[157]) | (~t[151] & t[152] & t[153] & t[154] & ~t[157]) | (~t[151] & t[152] & t[155] & t[156] & ~t[157]) | (t[151] & ~t[153] & ~t[155] & t[157]) | (~t[151] & t[153] & t[155] & t[157]);
  assign t[123] = (t[151] & t[152] & ~t[153] & t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[153] & ~t[154] & t[155] & ~t[156] & t[157]) | (~t[152] & t[153] & ~t[154] & ~t[155] & ~t[157]) | (~t[151] & t[153] & ~t[154] & ~t[155] & ~t[156]) | (~t[151] & ~t[152] & t[153] & ~t[156] & ~t[157]) | (~t[151] & t[153] & t[154] & ~t[155] & t[156]) | (t[153] & ~t[154] & t[156] & ~t[157]);
  assign t[124] = (t[158] & ~t[160] & ~t[161] & ~t[162] & ~t[163]) | (t[158] & ~t[159] & ~t[161] & ~t[162] & ~t[164]) | (t[158] & ~t[159] & ~t[160] & ~t[163] & ~t[164]) | (~t[158] & t[159] & t[160] & t[161] & ~t[164]) | (~t[158] & t[159] & t[162] & t[163] & ~t[164]) | (t[158] & ~t[160] & ~t[162] & t[164]) | (~t[158] & t[160] & t[162] & t[164]);
  assign t[125] = (t[158] & t[159] & ~t[160] & t[161] & ~t[162] & ~t[164]) | (t[158] & ~t[160] & ~t[161] & t[162] & ~t[163] & t[164]) | (~t[159] & t[160] & ~t[161] & ~t[162] & ~t[164]) | (~t[158] & t[160] & ~t[161] & ~t[162] & ~t[163]) | (~t[158] & ~t[159] & t[160] & ~t[163] & ~t[164]) | (~t[158] & t[160] & t[161] & ~t[162] & t[163]) | (t[160] & ~t[161] & t[163] & ~t[164]);
  assign t[126] = (t[165] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (t[165] & ~t[166] & ~t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[166] & ~t[167] & ~t[170] & ~t[171]) | (~t[165] & t[166] & t[167] & t[168] & ~t[171]) | (~t[165] & t[166] & t[169] & t[170] & ~t[171]) | (t[165] & ~t[167] & ~t[169] & t[171]) | (~t[165] & t[167] & t[169] & t[171]);
  assign t[127] = (t[165] & t[166] & ~t[167] & t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[167] & ~t[168] & t[169] & ~t[170] & t[171]) | (~t[166] & t[167] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[166] & t[167] & ~t[170] & ~t[171]) | (~t[165] & t[167] & t[168] & ~t[169] & t[170]) | (t[167] & ~t[168] & t[170] & ~t[171]);
  assign t[128] = (t[152] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (~t[151] & t[152] & ~t[154] & ~t[155] & ~t[157]) | (~t[151] & t[152] & ~t[153] & ~t[156] & ~t[157]) | (t[151] & ~t[152] & t[153] & t[154] & ~t[157]) | (t[151] & ~t[152] & t[155] & t[156] & ~t[157]) | (t[152] & ~t[154] & ~t[156] & t[157]) | (~t[152] & t[154] & t[156] & t[157]);
  assign t[129] = (t[151] & t[152] & t[153] & ~t[154] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & ~t[154] & ~t[155] & t[156] & t[157]) | (~t[152] & ~t[153] & t[154] & ~t[155] & ~t[156]) | (~t[151] & ~t[153] & t[154] & ~t[156] & ~t[157]) | (~t[151] & ~t[152] & t[154] & ~t[155] & ~t[157]) | (~t[152] & t[153] & t[154] & t[155] & ~t[156]) | (~t[153] & t[154] & t[155] & ~t[157]);
  assign t[12] = t[22] ^ t[23];
  assign t[130] = (t[151] & t[152] & ~t[153] & ~t[155] & t[156] & ~t[157]) | (t[151] & t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[157]) | (~t[151] & ~t[153] & ~t[154] & t[155] & ~t[156]) | (~t[151] & ~t[152] & ~t[154] & t[155] & ~t[157]) | (~t[151] & ~t[153] & t[154] & t[155] & t[156]) | (t[154] & t[155] & ~t[156] & ~t[157]);
  assign t[131] = (t[151] & t[152] & ~t[154] & t[155] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & ~t[154] & ~t[155] & t[156]) | (~t[151] & ~t[154] & ~t[155] & t[156] & ~t[157]) | (~t[151] & ~t[152] & ~t[153] & t[156] & ~t[157]) | (~t[152] & t[153] & ~t[154] & t[155] & t[156]) | (t[153] & ~t[155] & t[156] & ~t[157]);
  assign t[132] = (t[159] & ~t[160] & ~t[161] & ~t[162] & ~t[163]) | (~t[158] & t[159] & ~t[161] & ~t[162] & ~t[164]) | (~t[158] & t[159] & ~t[160] & ~t[163] & ~t[164]) | (t[158] & ~t[159] & t[160] & t[161] & ~t[164]) | (t[158] & ~t[159] & t[162] & t[163] & ~t[164]) | (t[159] & ~t[161] & ~t[163] & t[164]) | (~t[159] & t[161] & t[163] & t[164]);
  assign t[133] = (t[158] & t[159] & t[160] & ~t[161] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & ~t[161] & ~t[162] & t[163] & t[164]) | (~t[159] & ~t[160] & t[161] & ~t[162] & ~t[163]) | (~t[158] & ~t[160] & t[161] & ~t[163] & ~t[164]) | (~t[158] & ~t[159] & t[161] & ~t[162] & ~t[164]) | (~t[159] & t[160] & t[161] & t[162] & ~t[163]) | (~t[160] & t[161] & t[162] & ~t[164]);
  assign t[134] = (t[158] & t[159] & ~t[160] & ~t[162] & t[163] & ~t[164]) | (t[158] & t[160] & ~t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[160] & t[162] & ~t[163] & ~t[164]) | (~t[158] & ~t[160] & ~t[161] & t[162] & ~t[163]) | (~t[158] & ~t[159] & ~t[161] & t[162] & ~t[164]) | (~t[158] & ~t[160] & t[161] & t[162] & t[163]) | (t[161] & t[162] & ~t[163] & ~t[164]);
  assign t[135] = (t[158] & t[159] & ~t[161] & t[162] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[160] & ~t[161] & ~t[162] & t[163]) | (~t[158] & ~t[161] & ~t[162] & t[163] & ~t[164]) | (~t[158] & ~t[159] & ~t[160] & t[163] & ~t[164]) | (~t[159] & t[160] & ~t[161] & t[162] & t[163]) | (t[160] & ~t[162] & t[163] & ~t[164]);
  assign t[136] = (t[166] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & t[166] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[166] & ~t[167] & ~t[170] & ~t[171]) | (t[165] & ~t[166] & t[167] & t[168] & ~t[171]) | (t[165] & ~t[166] & t[169] & t[170] & ~t[171]) | (t[166] & ~t[168] & ~t[170] & t[171]) | (~t[166] & t[168] & t[170] & t[171]);
  assign t[137] = (t[165] & t[166] & t[167] & ~t[168] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & ~t[168] & ~t[169] & t[170] & t[171]) | (~t[166] & ~t[167] & t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[167] & t[168] & ~t[170] & ~t[171]) | (~t[165] & ~t[166] & t[168] & ~t[169] & ~t[171]) | (~t[166] & t[167] & t[168] & t[169] & ~t[170]) | (~t[167] & t[168] & t[169] & ~t[171]);
  assign t[138] = (t[165] & t[166] & ~t[167] & ~t[169] & t[170] & ~t[171]) | (t[165] & t[167] & ~t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & t[169] & ~t[170] & ~t[171]) | (~t[165] & ~t[167] & ~t[168] & t[169] & ~t[170]) | (~t[165] & ~t[166] & ~t[168] & t[169] & ~t[171]) | (~t[165] & ~t[167] & t[168] & t[169] & t[170]) | (t[168] & t[169] & ~t[170] & ~t[171]);
  assign t[139] = (t[165] & t[166] & ~t[168] & t[169] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & ~t[168] & ~t[169] & t[170]) | (~t[165] & ~t[168] & ~t[169] & t[170] & ~t[171]) | (~t[165] & ~t[166] & ~t[167] & t[170] & ~t[171]) | (~t[166] & t[167] & ~t[168] & t[169] & t[170]) | (t[167] & ~t[169] & t[170] & ~t[171]);
  assign t[13] = t[24] & t[25];
  assign t[140] = (t[144] & t[145] & ~t[146] & t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[146] & ~t[147] & t[148] & ~t[149] & t[150]) | (~t[145] & t[146] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[145] & t[146] & ~t[149] & ~t[150]) | (~t[144] & t[146] & t[147] & ~t[148] & t[149]) | (t[146] & ~t[147] & t[149] & ~t[150]);
  assign t[141] = (t[145] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & t[145] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[145] & ~t[146] & ~t[149] & ~t[150]) | (t[144] & ~t[145] & t[146] & t[147] & ~t[150]) | (t[144] & ~t[145] & t[148] & t[149] & ~t[150]) | (t[145] & ~t[147] & ~t[149] & t[150]) | (~t[145] & t[147] & t[149] & t[150]);
  assign t[142] = (t[144] & t[145] & t[146] & ~t[147] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[147] & ~t[148] & t[149] & t[150]) | (~t[145] & ~t[146] & t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[146] & t[147] & ~t[149] & ~t[150]) | (~t[144] & ~t[145] & t[147] & ~t[148] & ~t[150]) | (~t[145] & t[146] & t[147] & t[148] & ~t[149]) | (~t[146] & t[147] & t[148] & ~t[150]);
  assign t[143] = (t[144] & t[145] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[144] & ~t[145] & ~t[146] & t[149] & ~t[150]) | (~t[145] & t[146] & ~t[147] & t[148] & t[149]) | (t[146] & ~t[148] & t[149] & ~t[150]);
  assign t[144] = t[172] ^ x[7];
  assign t[145] = t[173] ^ x[45];
  assign t[146] = t[174] ^ x[43];
  assign t[147] = t[175] ^ x[46];
  assign t[148] = t[176] ^ x[8];
  assign t[149] = t[177] ^ x[47];
  assign t[14] = t[82] & t[26];
  assign t[150] = t[178] ^ x[6];
  assign t[151] = t[179] ^ x[14];
  assign t[152] = t[180] ^ x[30];
  assign t[153] = t[181] ^ x[15];
  assign t[154] = t[182] ^ x[31];
  assign t[155] = t[183] ^ x[32];
  assign t[156] = t[184] ^ x[33];
  assign t[157] = t[185] ^ x[13];
  assign t[158] = t[186] ^ x[21];
  assign t[159] = t[187] ^ x[34];
  assign t[15] = t[27] & t[28];
  assign t[160] = t[188] ^ x[22];
  assign t[161] = t[189] ^ x[35];
  assign t[162] = t[190] ^ x[36];
  assign t[163] = t[191] ^ x[37];
  assign t[164] = t[192] ^ x[20];
  assign t[165] = t[193] ^ x[28];
  assign t[166] = t[194] ^ x[38];
  assign t[167] = t[195] ^ x[29];
  assign t[168] = t[196] ^ x[39];
  assign t[169] = t[197] ^ x[40];
  assign t[16] = t[29] ^ t[27];
  assign t[170] = t[198] ^ x[41];
  assign t[171] = t[199] ^ x[27];
  assign t[172] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[173] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[174] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[175] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[176] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[177] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[178] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[179] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[181] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[182] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[183] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[184] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[185] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[186] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[187] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[188] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[189] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[18] = t[83] & t[31];
  assign t[190] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[191] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[192] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[193] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[194] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[195] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[196] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[197] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[198] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[199] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[84] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[85]);
  assign t[28] = ~(t[82] ^ t[27]);
  assign t[29] = t[86] ^ t[85];
  assign t[2] = ~(t[4] ^ t[81]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[87]);
  assign t[33] = ~(t[83] ^ t[32]);
  assign t[34] = t[88] ^ t[87];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[89]);
  assign t[38] = ~(t[84] ^ t[37]);
  assign t[39] = t[90] ^ t[89];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[82] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[82] ^ t[50];
  assign t[44] = t[83] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[83] ^ t[51];
  assign t[47] = t[84] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[84] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[85] ^ t[91];
  assign t[51] = t[87] ^ t[92];
  assign t[52] = t[89] ^ t[93];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[94]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61] ^ t[62]);
  assign t[59] = ~(t[63] ^ t[64]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[65] ^ t[66]);
  assign t[61] = t[67] ^ t[15];
  assign t[62] = t[8] ^ t[68];
  assign t[63] = t[69] ^ t[19];
  assign t[64] = t[10] ^ t[70];
  assign t[65] = t[71] ^ t[23];
  assign t[66] = t[12] ^ t[72];
  assign t[67] = t[29] ^ t[42];
  assign t[68] = t[82] ^ t[27];
  assign t[69] = t[34] ^ t[45];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[83] ^ t[32];
  assign t[71] = t[39] ^ t[48];
  assign t[72] = t[84] ^ t[37];
  assign t[73] = x[0] ? x[44] : t[74];
  assign t[74] = ~(t[75] ^ t[76]);
  assign t[75] = ~(t[77] ^ t[95]);
  assign t[76] = ~(t[78] ^ t[79]);
  assign t[77] = ~t[80];
  assign t[78] = ~(t[61]);
  assign t[79] = ~(t[63]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = ~(t[65]);
  assign t[81] = (t[96] & ~t[97]) | (~t[96] & t[97]);
  assign t[82] = (t[98] & ~t[99]) | (~t[98] & t[99]);
  assign t[83] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[84] = (t[102] & ~t[103]) | (~t[102] & t[103]);
  assign t[85] = (t[98] & ~t[105] & ~t[107]) | (~t[104] & t[105] & ~t[106]) | (~t[98] & ~t[105] & t[107]) | (t[104] & t[105] & t[106]);
  assign t[86] = (t[98] & ~t[106]) | (~t[98] & t[106]);
  assign t[87] = (t[100] & ~t[109] & ~t[111]) | (~t[108] & t[109] & ~t[110]) | (~t[100] & ~t[109] & t[111]) | (t[108] & t[109] & t[110]);
  assign t[88] = (t[100] & ~t[110]) | (~t[100] & t[110]);
  assign t[89] = (t[102] & ~t[113] & ~t[115]) | (~t[112] & t[113] & ~t[114]) | (~t[102] & ~t[113] & t[115]) | (t[112] & t[113] & t[114]);
  assign t[8] = t[14] ^ t[15];
  assign t[90] = (t[102] & ~t[114]) | (~t[102] & t[114]);
  assign t[91] = (t[98] & ~t[105] & ~t[106]) | (~t[104] & t[105] & ~t[107]) | (~t[98] & ~t[105] & t[106]) | (t[104] & t[105] & t[107]);
  assign t[92] = (t[100] & ~t[109] & ~t[110]) | (~t[108] & t[109] & ~t[111]) | (~t[100] & ~t[109] & t[110]) | (t[108] & t[109] & t[111]);
  assign t[93] = (t[102] & ~t[113] & ~t[114]) | (~t[112] & t[113] & ~t[115]) | (~t[102] & ~t[113] & t[114]) | (t[112] & t[113] & t[115]);
  assign t[94] = (t[96] & ~t[116]) | (~t[96] & t[116]);
  assign t[95] = (t[96] & ~t[118] & ~t[97]) | (~t[117] & t[118] & ~t[119]) | (~t[96] & ~t[118] & t[97]) | (t[117] & t[118] & t[119]);
  assign t[96] = t[120] ^ x[7];
  assign t[97] = t[121] ^ x[8];
  assign t[98] = t[122] ^ x[14];
  assign t[99] = t[123] ^ x[15];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53] & ~t[73]) | (~t[0] & t[53] & ~t[73]) | (~t[0] & ~t[53] & t[73]) | (t[0] & t[53] & t[73]);
endmodule

module R2ind156(x, y);
 input [46:0] x;
 output y;

 wire [179:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[123] ^ x[46];
  assign t[101] = (t[124] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[127] & ~t[128] & ~t[130]) | (t[124] & ~t[125] & ~t[126] & ~t[129] & ~t[130]) | (~t[124] & t[125] & t[126] & t[127] & ~t[130]) | (~t[124] & t[125] & t[128] & t[129] & ~t[130]) | (t[124] & ~t[126] & ~t[128] & t[130]) | (~t[124] & t[126] & t[128] & t[130]);
  assign t[102] = (t[124] & t[125] & ~t[126] & ~t[128] & t[129] & ~t[130]) | (t[124] & t[126] & ~t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & t[128] & ~t[129] & ~t[130]) | (~t[124] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[124] & ~t[125] & ~t[127] & t[128] & ~t[130]) | (~t[124] & ~t[126] & t[127] & t[128] & t[129]) | (t[127] & t[128] & ~t[129] & ~t[130]);
  assign t[103] = (t[131] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[132] & ~t[133] & ~t[136] & ~t[137]) | (~t[131] & t[132] & t[133] & t[134] & ~t[137]) | (~t[131] & t[132] & t[135] & t[136] & ~t[137]) | (t[131] & ~t[133] & ~t[135] & t[137]) | (~t[131] & t[133] & t[135] & t[137]);
  assign t[104] = (t[131] & t[132] & ~t[133] & t[134] & ~t[135] & ~t[137]) | (t[131] & ~t[133] & ~t[134] & t[135] & ~t[136] & t[137]) | (~t[132] & t[133] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[132] & t[133] & ~t[136] & ~t[137]) | (~t[131] & t[133] & t[134] & ~t[135] & t[136]) | (t[133] & ~t[134] & t[136] & ~t[137]);
  assign t[105] = (t[138] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[139] & ~t[140] & ~t[143] & ~t[144]) | (~t[138] & t[139] & t[140] & t[141] & ~t[144]) | (~t[138] & t[139] & t[142] & t[143] & ~t[144]) | (t[138] & ~t[140] & ~t[142] & t[144]) | (~t[138] & t[140] & t[142] & t[144]);
  assign t[106] = (t[138] & t[139] & ~t[140] & t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[140] & ~t[141] & t[142] & ~t[143] & t[144]) | (~t[139] & t[140] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[139] & t[140] & ~t[143] & ~t[144]) | (~t[138] & t[140] & t[141] & ~t[142] & t[143]) | (t[140] & ~t[141] & t[143] & ~t[144]);
  assign t[107] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[108] = (t[145] & t[146] & ~t[147] & t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[147] & ~t[148] & t[149] & ~t[150] & t[151]) | (~t[146] & t[147] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[146] & t[147] & ~t[150] & ~t[151]) | (~t[145] & t[147] & t[148] & ~t[149] & t[150]) | (t[147] & ~t[148] & t[150] & ~t[151]);
  assign t[109] = (t[132] & ~t[133] & ~t[134] & ~t[135] & ~t[136]) | (~t[131] & t[132] & ~t[134] & ~t[135] & ~t[137]) | (~t[131] & t[132] & ~t[133] & ~t[136] & ~t[137]) | (t[131] & ~t[132] & t[133] & t[134] & ~t[137]) | (t[131] & ~t[132] & t[135] & t[136] & ~t[137]) | (t[132] & ~t[134] & ~t[136] & t[137]) | (~t[132] & t[134] & t[136] & t[137]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[131] & t[132] & t[133] & ~t[134] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & ~t[134] & ~t[135] & t[136] & t[137]) | (~t[132] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (~t[131] & ~t[133] & t[134] & ~t[136] & ~t[137]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[137]) | (~t[132] & t[133] & t[134] & t[135] & ~t[136]) | (~t[133] & t[134] & t[135] & ~t[137]);
  assign t[111] = (t[131] & t[132] & ~t[133] & ~t[135] & t[136] & ~t[137]) | (t[131] & t[133] & ~t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & t[135] & ~t[136] & ~t[137]) | (~t[131] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[131] & ~t[132] & ~t[134] & t[135] & ~t[137]) | (~t[131] & ~t[133] & t[134] & t[135] & t[136]) | (t[134] & t[135] & ~t[136] & ~t[137]);
  assign t[112] = (t[131] & t[132] & ~t[134] & t[135] & ~t[136] & ~t[137]) | (t[132] & ~t[133] & t[134] & ~t[135] & ~t[136] & t[137]) | (~t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[134] & ~t[135] & t[136] & ~t[137]) | (~t[131] & ~t[132] & ~t[133] & t[136] & ~t[137]) | (~t[132] & t[133] & ~t[134] & t[135] & t[136]) | (t[133] & ~t[135] & t[136] & ~t[137]);
  assign t[113] = (t[139] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & t[139] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[139] & ~t[140] & ~t[143] & ~t[144]) | (t[138] & ~t[139] & t[140] & t[141] & ~t[144]) | (t[138] & ~t[139] & t[142] & t[143] & ~t[144]) | (t[139] & ~t[141] & ~t[143] & t[144]) | (~t[139] & t[141] & t[143] & t[144]);
  assign t[114] = (t[138] & t[139] & t[140] & ~t[141] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & ~t[141] & ~t[142] & t[143] & t[144]) | (~t[139] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[140] & t[141] & ~t[143] & ~t[144]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[144]) | (~t[139] & t[140] & t[141] & t[142] & ~t[143]) | (~t[140] & t[141] & t[142] & ~t[144]);
  assign t[115] = (t[138] & t[139] & ~t[140] & ~t[142] & t[143] & ~t[144]) | (t[138] & t[140] & ~t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & t[142] & ~t[143] & ~t[144]) | (~t[138] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[138] & ~t[139] & ~t[141] & t[142] & ~t[144]) | (~t[138] & ~t[140] & t[141] & t[142] & t[143]) | (t[141] & t[142] & ~t[143] & ~t[144]);
  assign t[116] = (t[138] & t[139] & ~t[141] & t[142] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[141] & ~t[142] & t[143] & ~t[144]) | (~t[138] & ~t[139] & ~t[140] & t[143] & ~t[144]) | (~t[139] & t[140] & ~t[141] & t[142] & t[143]) | (t[140] & ~t[142] & t[143] & ~t[144]);
  assign t[117] = (t[146] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (~t[145] & t[146] & ~t[148] & ~t[149] & ~t[151]) | (~t[145] & t[146] & ~t[147] & ~t[150] & ~t[151]) | (t[145] & ~t[146] & t[147] & t[148] & ~t[151]) | (t[145] & ~t[146] & t[149] & t[150] & ~t[151]) | (t[146] & ~t[148] & ~t[150] & t[151]) | (~t[146] & t[148] & t[150] & t[151]);
  assign t[118] = (t[145] & t[146] & t[147] & ~t[148] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & ~t[148] & ~t[149] & t[150] & t[151]) | (~t[146] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (~t[145] & ~t[147] & t[148] & ~t[150] & ~t[151]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[151]) | (~t[146] & t[147] & t[148] & t[149] & ~t[150]) | (~t[147] & t[148] & t[149] & ~t[151]);
  assign t[119] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[145] & t[146] & ~t[148] & t[149] & ~t[150] & ~t[151]) | (t[146] & ~t[147] & t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[148] & ~t[149] & t[150] & ~t[151]) | (~t[145] & ~t[146] & ~t[147] & t[150] & ~t[151]) | (~t[146] & t[147] & ~t[148] & t[149] & t[150]) | (t[147] & ~t[149] & t[150] & ~t[151]);
  assign t[121] = (t[125] & ~t[126] & ~t[127] & ~t[128] & ~t[129]) | (~t[124] & t[125] & ~t[127] & ~t[128] & ~t[130]) | (~t[124] & t[125] & ~t[126] & ~t[129] & ~t[130]) | (t[124] & ~t[125] & t[126] & t[127] & ~t[130]) | (t[124] & ~t[125] & t[128] & t[129] & ~t[130]) | (t[125] & ~t[127] & ~t[129] & t[130]) | (~t[125] & t[127] & t[129] & t[130]);
  assign t[122] = (t[124] & t[125] & t[126] & ~t[127] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & ~t[127] & ~t[128] & t[129] & t[130]) | (~t[125] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (~t[124] & ~t[126] & t[127] & ~t[129] & ~t[130]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[130]) | (~t[125] & t[126] & t[127] & t[128] & ~t[129]) | (~t[126] & t[127] & t[128] & ~t[130]);
  assign t[123] = (t[124] & t[125] & ~t[127] & t[128] & ~t[129] & ~t[130]) | (t[125] & ~t[126] & t[127] & ~t[128] & ~t[129] & t[130]) | (~t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[127] & ~t[128] & t[129] & ~t[130]) | (~t[124] & ~t[125] & ~t[126] & t[129] & ~t[130]) | (~t[125] & t[126] & ~t[127] & t[128] & t[129]) | (t[126] & ~t[128] & t[129] & ~t[130]);
  assign t[124] = t[152] ^ x[8];
  assign t[125] = t[153] ^ x[44];
  assign t[126] = t[154] ^ x[6];
  assign t[127] = t[155] ^ x[45];
  assign t[128] = t[156] ^ x[9];
  assign t[129] = t[157] ^ x[46];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[7];
  assign t[131] = t[159] ^ x[15];
  assign t[132] = t[160] ^ x[31];
  assign t[133] = t[161] ^ x[16];
  assign t[134] = t[162] ^ x[32];
  assign t[135] = t[163] ^ x[33];
  assign t[136] = t[164] ^ x[34];
  assign t[137] = t[165] ^ x[14];
  assign t[138] = t[166] ^ x[22];
  assign t[139] = t[167] ^ x[35];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[168] ^ x[23];
  assign t[141] = t[169] ^ x[36];
  assign t[142] = t[170] ^ x[37];
  assign t[143] = t[171] ^ x[38];
  assign t[144] = t[172] ^ x[21];
  assign t[145] = t[173] ^ x[29];
  assign t[146] = t[174] ^ x[39];
  assign t[147] = t[175] ^ x[30];
  assign t[148] = t[176] ^ x[40];
  assign t[149] = t[177] ^ x[41];
  assign t[14] = t[65] & t[26];
  assign t[150] = t[178] ^ x[42];
  assign t[151] = t[179] ^ x[28];
  assign t[152] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[153] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[154] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[155] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[156] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[157] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[158] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[159] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[161] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[162] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[163] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[164] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[165] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[166] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[167] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[168] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[169] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[171] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[172] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[173] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[174] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[175] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[176] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[177] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[178] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[179] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[17] = t[30] ^ t[15];
  assign t[18] = t[66] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[67] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[68]);
  assign t[28] = ~(t[65] ^ t[27]);
  assign t[29] = t[69] ^ t[68];
  assign t[2] = ~(t[4] ^ t[64]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[70]);
  assign t[33] = ~(t[66] ^ t[32]);
  assign t[34] = t[71] ^ t[70];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[72]);
  assign t[38] = ~(t[67] ^ t[37]);
  assign t[39] = t[73] ^ t[72];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[65] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[65] ^ t[50];
  assign t[44] = t[66] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[66] ^ t[51];
  assign t[47] = t[67] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[67] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[68] ^ t[74];
  assign t[51] = t[70] ^ t[75];
  assign t[52] = t[72] ^ t[76];
  assign t[53] = x[0] ? x[43] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[77]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = t[50] ^ t[15];
  assign t[62] = t[51] ^ t[19];
  assign t[63] = t[52] ^ t[23];
  assign t[64] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[67] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[68] = (t[80] & ~t[87] & ~t[89]) | (~t[86] & t[87] & ~t[88]) | (~t[80] & ~t[87] & t[89]) | (t[86] & t[87] & t[88]);
  assign t[69] = (t[80] & ~t[88]) | (~t[80] & t[88]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[82] & ~t[91] & ~t[93]) | (~t[90] & t[91] & ~t[92]) | (~t[82] & ~t[91] & t[93]) | (t[90] & t[91] & t[92]);
  assign t[71] = (t[82] & ~t[92]) | (~t[82] & t[92]);
  assign t[72] = (t[84] & ~t[95] & ~t[97]) | (~t[94] & t[95] & ~t[96]) | (~t[84] & ~t[95] & t[97]) | (t[94] & t[95] & t[96]);
  assign t[73] = (t[84] & ~t[96]) | (~t[84] & t[96]);
  assign t[74] = (t[80] & ~t[87] & ~t[88]) | (~t[86] & t[87] & ~t[89]) | (~t[80] & ~t[87] & t[88]) | (t[86] & t[87] & t[89]);
  assign t[75] = (t[82] & ~t[91] & ~t[92]) | (~t[90] & t[91] & ~t[93]) | (~t[82] & ~t[91] & t[92]) | (t[90] & t[91] & t[93]);
  assign t[76] = (t[84] & ~t[95] & ~t[96]) | (~t[94] & t[95] & ~t[97]) | (~t[84] & ~t[95] & t[96]) | (t[94] & t[95] & t[97]);
  assign t[77] = (t[78] & ~t[99] & ~t[100]) | (~t[98] & t[99] & ~t[79]) | (~t[78] & ~t[99] & t[100]) | (t[98] & t[99] & t[79]);
  assign t[78] = t[101] ^ x[8];
  assign t[79] = t[102] ^ x[9];
  assign t[7] = t[12] ^ t[13];
  assign t[80] = t[103] ^ x[15];
  assign t[81] = t[104] ^ x[16];
  assign t[82] = t[105] ^ x[22];
  assign t[83] = t[106] ^ x[23];
  assign t[84] = t[107] ^ x[29];
  assign t[85] = t[108] ^ x[30];
  assign t[86] = t[109] ^ x[31];
  assign t[87] = t[110] ^ x[32];
  assign t[88] = t[111] ^ x[33];
  assign t[89] = t[112] ^ x[34];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[113] ^ x[35];
  assign t[91] = t[114] ^ x[36];
  assign t[92] = t[115] ^ x[37];
  assign t[93] = t[116] ^ x[38];
  assign t[94] = t[117] ^ x[39];
  assign t[95] = t[118] ^ x[40];
  assign t[96] = t[119] ^ x[41];
  assign t[97] = t[120] ^ x[42];
  assign t[98] = t[121] ^ x[44];
  assign t[99] = t[122] ^ x[45];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind157(x, y);
 input [46:0] x;
 output y;

 wire [182:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[123] ^ x[42];
  assign t[101] = t[124] ^ x[44];
  assign t[102] = t[125] ^ x[45];
  assign t[103] = t[126] ^ x[46];
  assign t[104] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[105] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[106] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[107] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[108] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[109] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[111] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[112] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[113] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[114] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[115] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[116] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[117] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[118] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[119] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[11] = t[20] & t[21];
  assign t[120] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[121] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[122] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[123] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[124] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[125] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[126] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[127] = t[155] ^ x[8];
  assign t[128] = t[156] ^ x[44];
  assign t[129] = t[157] ^ x[6];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[45];
  assign t[131] = t[159] ^ x[9];
  assign t[132] = t[160] ^ x[46];
  assign t[133] = t[161] ^ x[7];
  assign t[134] = t[162] ^ x[15];
  assign t[135] = t[163] ^ x[31];
  assign t[136] = t[164] ^ x[16];
  assign t[137] = t[165] ^ x[32];
  assign t[138] = t[166] ^ x[33];
  assign t[139] = t[167] ^ x[34];
  assign t[13] = t[24] & t[25];
  assign t[140] = t[168] ^ x[14];
  assign t[141] = t[169] ^ x[22];
  assign t[142] = t[170] ^ x[35];
  assign t[143] = t[171] ^ x[23];
  assign t[144] = t[172] ^ x[36];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[38];
  assign t[147] = t[175] ^ x[21];
  assign t[148] = t[176] ^ x[29];
  assign t[149] = t[177] ^ x[39];
  assign t[14] = t[68] & t[26];
  assign t[150] = t[178] ^ x[30];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[42];
  assign t[154] = t[182] ^ x[28];
  assign t[155] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[156] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[157] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[158] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[159] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[15] = t[27] & t[28];
  assign t[160] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[161] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[162] = (x[10] & ~x[11] & ~x[12]) | (~x[10] & x[11] & ~x[12]) | (~x[10] & ~x[11] & x[12]) | (x[10] & x[11] & x[12]);
  assign t[163] = (x[10] & ~x[11] & ~x[13]) | (~x[10] & x[11] & ~x[13]) | (~x[10] & ~x[11] & x[13]) | (x[10] & x[11] & x[13]);
  assign t[164] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[165] = (x[10] & ~x[13]) | (~x[10] & x[13]);
  assign t[166] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[167] = (x[11] & ~x[13]) | (~x[11] & x[13]);
  assign t[168] = (x[12] & ~x[13]) | (~x[12] & x[13]);
  assign t[169] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[16] = t[29] ^ t[27];
  assign t[170] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[171] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[172] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[173] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[174] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[175] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[176] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[177] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[178] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[179] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[17] = t[30] ^ t[15];
  assign t[180] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[181] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[182] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[18] = t[69] & t[31];
  assign t[19] = t[32] & t[33];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[34] ^ t[32];
  assign t[21] = t[35] ^ t[19];
  assign t[22] = t[70] & t[36];
  assign t[23] = t[37] & t[38];
  assign t[24] = t[39] ^ t[37];
  assign t[25] = t[40] ^ t[23];
  assign t[26] = t[41] ^ t[42];
  assign t[27] = ~(t[71]);
  assign t[28] = ~(t[68] ^ t[27]);
  assign t[29] = t[72] ^ t[71];
  assign t[2] = ~(t[4] ^ t[67]);
  assign t[30] = ~(t[43] ^ t[16]);
  assign t[31] = t[44] ^ t[45];
  assign t[32] = ~(t[73]);
  assign t[33] = ~(t[69] ^ t[32]);
  assign t[34] = t[74] ^ t[73];
  assign t[35] = ~(t[46] ^ t[20]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = ~(t[75]);
  assign t[38] = ~(t[70] ^ t[37]);
  assign t[39] = t[76] ^ t[75];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = ~(t[49] ^ t[24]);
  assign t[41] = t[68] ^ t[29];
  assign t[42] = t[27] & t[43];
  assign t[43] = t[68] ^ t[50];
  assign t[44] = t[69] ^ t[34];
  assign t[45] = t[32] & t[46];
  assign t[46] = t[69] ^ t[51];
  assign t[47] = t[70] ^ t[39];
  assign t[48] = t[37] & t[49];
  assign t[49] = t[70] ^ t[52];
  assign t[4] = ~t[7];
  assign t[50] = t[71] ^ t[77];
  assign t[51] = t[73] ^ t[78];
  assign t[52] = t[75] ^ t[79];
  assign t[53] = x[0] ? x[43] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[80]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = t[64] ^ t[15];
  assign t[62] = t[65] ^ t[19];
  assign t[63] = t[66] ^ t[23];
  assign t[64] = t[29] ^ t[42];
  assign t[65] = t[34] ^ t[45];
  assign t[66] = t[39] ^ t[48];
  assign t[67] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[68] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[69] = (t[85] & ~t[86]) | (~t[85] & t[86]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[87] & ~t[88]) | (~t[87] & t[88]);
  assign t[71] = (t[83] & ~t[90] & ~t[92]) | (~t[89] & t[90] & ~t[91]) | (~t[83] & ~t[90] & t[92]) | (t[89] & t[90] & t[91]);
  assign t[72] = (t[83] & ~t[91]) | (~t[83] & t[91]);
  assign t[73] = (t[85] & ~t[94] & ~t[96]) | (~t[93] & t[94] & ~t[95]) | (~t[85] & ~t[94] & t[96]) | (t[93] & t[94] & t[95]);
  assign t[74] = (t[85] & ~t[95]) | (~t[85] & t[95]);
  assign t[75] = (t[87] & ~t[98] & ~t[100]) | (~t[97] & t[98] & ~t[99]) | (~t[87] & ~t[98] & t[100]) | (t[97] & t[98] & t[99]);
  assign t[76] = (t[87] & ~t[99]) | (~t[87] & t[99]);
  assign t[77] = (t[83] & ~t[90] & ~t[91]) | (~t[89] & t[90] & ~t[92]) | (~t[83] & ~t[90] & t[91]) | (t[89] & t[90] & t[92]);
  assign t[78] = (t[85] & ~t[94] & ~t[95]) | (~t[93] & t[94] & ~t[96]) | (~t[85] & ~t[94] & t[95]) | (t[93] & t[94] & t[96]);
  assign t[79] = (t[87] & ~t[98] & ~t[99]) | (~t[97] & t[98] & ~t[100]) | (~t[87] & ~t[98] & t[99]) | (t[97] & t[98] & t[100]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (t[81] & ~t[102] & ~t[82]) | (~t[101] & t[102] & ~t[103]) | (~t[81] & ~t[102] & t[82]) | (t[101] & t[102] & t[103]);
  assign t[81] = t[104] ^ x[8];
  assign t[82] = t[105] ^ x[9];
  assign t[83] = t[106] ^ x[15];
  assign t[84] = t[107] ^ x[16];
  assign t[85] = t[108] ^ x[22];
  assign t[86] = t[109] ^ x[23];
  assign t[87] = t[110] ^ x[29];
  assign t[88] = t[111] ^ x[30];
  assign t[89] = t[112] ^ x[31];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[113] ^ x[32];
  assign t[91] = t[114] ^ x[33];
  assign t[92] = t[115] ^ x[34];
  assign t[93] = t[116] ^ x[35];
  assign t[94] = t[117] ^ x[36];
  assign t[95] = t[118] ^ x[37];
  assign t[96] = t[119] ^ x[38];
  assign t[97] = t[120] ^ x[39];
  assign t[98] = t[121] ^ x[40];
  assign t[99] = t[122] ^ x[41];
  assign t[9] = t[16] & t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind158(x, y);
 input [46:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[124] ^ x[45];
  assign t[101] = t[125] ^ x[46];
  assign t[102] = (t[126] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (t[126] & ~t[127] & ~t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[127] & ~t[128] & ~t[131] & ~t[132]) | (~t[126] & t[127] & t[128] & t[129] & ~t[132]) | (~t[126] & t[127] & t[130] & t[131] & ~t[132]) | (t[126] & ~t[128] & ~t[130] & t[132]) | (~t[126] & t[128] & t[130] & t[132]);
  assign t[103] = (t[126] & t[127] & ~t[128] & t[129] & ~t[130] & ~t[132]) | (t[126] & ~t[128] & ~t[129] & t[130] & ~t[131] & t[132]) | (~t[127] & t[128] & ~t[129] & ~t[130] & ~t[132]) | (~t[126] & t[128] & ~t[129] & ~t[130] & ~t[131]) | (~t[126] & ~t[127] & t[128] & ~t[131] & ~t[132]) | (~t[126] & t[128] & t[129] & ~t[130] & t[131]) | (t[128] & ~t[129] & t[131] & ~t[132]);
  assign t[104] = (t[133] & ~t[135] & ~t[136] & ~t[137] & ~t[138]) | (t[133] & ~t[134] & ~t[136] & ~t[137] & ~t[139]) | (t[133] & ~t[134] & ~t[135] & ~t[138] & ~t[139]) | (~t[133] & t[134] & t[135] & t[136] & ~t[139]) | (~t[133] & t[134] & t[137] & t[138] & ~t[139]) | (t[133] & ~t[135] & ~t[137] & t[139]) | (~t[133] & t[135] & t[137] & t[139]);
  assign t[105] = (t[133] & t[134] & ~t[135] & t[136] & ~t[137] & ~t[139]) | (t[133] & ~t[135] & ~t[136] & t[137] & ~t[138] & t[139]) | (~t[134] & t[135] & ~t[136] & ~t[137] & ~t[139]) | (~t[133] & t[135] & ~t[136] & ~t[137] & ~t[138]) | (~t[133] & ~t[134] & t[135] & ~t[138] & ~t[139]) | (~t[133] & t[135] & t[136] & ~t[137] & t[138]) | (t[135] & ~t[136] & t[138] & ~t[139]);
  assign t[106] = (t[140] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (t[140] & ~t[141] & ~t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[141] & ~t[142] & ~t[145] & ~t[146]) | (~t[140] & t[141] & t[142] & t[143] & ~t[146]) | (~t[140] & t[141] & t[144] & t[145] & ~t[146]) | (t[140] & ~t[142] & ~t[144] & t[146]) | (~t[140] & t[142] & t[144] & t[146]);
  assign t[107] = (t[140] & t[141] & ~t[142] & t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[142] & ~t[143] & t[144] & ~t[145] & t[146]) | (~t[141] & t[142] & ~t[143] & ~t[144] & ~t[146]) | (~t[140] & t[142] & ~t[143] & ~t[144] & ~t[145]) | (~t[140] & ~t[141] & t[142] & ~t[145] & ~t[146]) | (~t[140] & t[142] & t[143] & ~t[144] & t[145]) | (t[142] & ~t[143] & t[145] & ~t[146]);
  assign t[108] = (t[147] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (t[147] & ~t[148] & ~t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[148] & ~t[149] & ~t[152] & ~t[153]) | (~t[147] & t[148] & t[149] & t[150] & ~t[153]) | (~t[147] & t[148] & t[151] & t[152] & ~t[153]) | (t[147] & ~t[149] & ~t[151] & t[153]) | (~t[147] & t[149] & t[151] & t[153]);
  assign t[109] = (t[147] & t[148] & ~t[149] & t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[149] & ~t[150] & t[151] & ~t[152] & t[153]) | (~t[148] & t[149] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[148] & t[149] & ~t[152] & ~t[153]) | (~t[147] & t[149] & t[150] & ~t[151] & t[152]) | (t[149] & ~t[150] & t[152] & ~t[153]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[133] & t[134] & ~t[135] & ~t[137] & t[138] & ~t[139]) | (t[133] & t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[139]) | (~t[133] & ~t[135] & ~t[136] & t[137] & ~t[138]) | (~t[133] & ~t[134] & ~t[136] & t[137] & ~t[139]) | (~t[133] & ~t[135] & t[136] & t[137] & t[138]) | (t[136] & t[137] & ~t[138] & ~t[139]);
  assign t[111] = (t[134] & ~t[135] & ~t[136] & ~t[137] & ~t[138]) | (~t[133] & t[134] & ~t[136] & ~t[137] & ~t[139]) | (~t[133] & t[134] & ~t[135] & ~t[138] & ~t[139]) | (t[133] & ~t[134] & t[135] & t[136] & ~t[139]) | (t[133] & ~t[134] & t[137] & t[138] & ~t[139]) | (t[134] & ~t[136] & ~t[138] & t[139]) | (~t[134] & t[136] & t[138] & t[139]);
  assign t[112] = (t[133] & t[134] & t[135] & ~t[136] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[136] & ~t[137] & t[138] & t[139]) | (~t[134] & ~t[135] & t[136] & ~t[137] & ~t[138]) | (~t[133] & ~t[135] & t[136] & ~t[138] & ~t[139]) | (~t[133] & ~t[134] & t[136] & ~t[137] & ~t[139]) | (~t[134] & t[135] & t[136] & t[137] & ~t[138]) | (~t[135] & t[136] & t[137] & ~t[139]);
  assign t[113] = (t[133] & t[134] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[135] & ~t[136] & ~t[137] & t[138]) | (~t[133] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[133] & ~t[134] & ~t[135] & t[138] & ~t[139]) | (~t[134] & t[135] & ~t[136] & t[137] & t[138]) | (t[135] & ~t[137] & t[138] & ~t[139]);
  assign t[114] = (t[140] & t[141] & ~t[142] & ~t[144] & t[145] & ~t[146]) | (t[140] & t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[146]) | (~t[140] & ~t[142] & ~t[143] & t[144] & ~t[145]) | (~t[140] & ~t[141] & ~t[143] & t[144] & ~t[146]) | (~t[140] & ~t[142] & t[143] & t[144] & t[145]) | (t[143] & t[144] & ~t[145] & ~t[146]);
  assign t[115] = (t[141] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (~t[140] & t[141] & ~t[143] & ~t[144] & ~t[146]) | (~t[140] & t[141] & ~t[142] & ~t[145] & ~t[146]) | (t[140] & ~t[141] & t[142] & t[143] & ~t[146]) | (t[140] & ~t[141] & t[144] & t[145] & ~t[146]) | (t[141] & ~t[143] & ~t[145] & t[146]) | (~t[141] & t[143] & t[145] & t[146]);
  assign t[116] = (t[140] & t[141] & t[142] & ~t[143] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[143] & ~t[144] & t[145] & t[146]) | (~t[141] & ~t[142] & t[143] & ~t[144] & ~t[145]) | (~t[140] & ~t[142] & t[143] & ~t[145] & ~t[146]) | (~t[140] & ~t[141] & t[143] & ~t[144] & ~t[146]) | (~t[141] & t[142] & t[143] & t[144] & ~t[145]) | (~t[142] & t[143] & t[144] & ~t[146]);
  assign t[117] = (t[140] & t[141] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & ~t[143] & ~t[144] & t[145]) | (~t[140] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[140] & ~t[141] & ~t[142] & t[145] & ~t[146]) | (~t[141] & t[142] & ~t[143] & t[144] & t[145]) | (t[142] & ~t[144] & t[145] & ~t[146]);
  assign t[118] = (t[147] & t[148] & ~t[149] & ~t[151] & t[152] & ~t[153]) | (t[147] & t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[153]) | (~t[147] & ~t[149] & ~t[150] & t[151] & ~t[152]) | (~t[147] & ~t[148] & ~t[150] & t[151] & ~t[153]) | (~t[147] & ~t[149] & t[150] & t[151] & t[152]) | (t[150] & t[151] & ~t[152] & ~t[153]);
  assign t[119] = (t[148] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (~t[147] & t[148] & ~t[150] & ~t[151] & ~t[153]) | (~t[147] & t[148] & ~t[149] & ~t[152] & ~t[153]) | (t[147] & ~t[148] & t[149] & t[150] & ~t[153]) | (t[147] & ~t[148] & t[151] & t[152] & ~t[153]) | (t[148] & ~t[150] & ~t[152] & t[153]) | (~t[148] & t[150] & t[152] & t[153]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = (t[147] & t[148] & t[149] & ~t[150] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[150] & ~t[151] & t[152] & t[153]) | (~t[148] & ~t[149] & t[150] & ~t[151] & ~t[152]) | (~t[147] & ~t[149] & t[150] & ~t[152] & ~t[153]) | (~t[147] & ~t[148] & t[150] & ~t[151] & ~t[153]) | (~t[148] & t[149] & t[150] & t[151] & ~t[152]) | (~t[149] & t[150] & t[151] & ~t[153]);
  assign t[121] = (t[147] & t[148] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & ~t[150] & ~t[151] & t[152]) | (~t[147] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[147] & ~t[148] & ~t[149] & t[152] & ~t[153]) | (~t[148] & t[149] & ~t[150] & t[151] & t[152]) | (t[149] & ~t[151] & t[152] & ~t[153]);
  assign t[122] = (t[127] & ~t[128] & ~t[129] & ~t[130] & ~t[131]) | (~t[126] & t[127] & ~t[129] & ~t[130] & ~t[132]) | (~t[126] & t[127] & ~t[128] & ~t[131] & ~t[132]) | (t[126] & ~t[127] & t[128] & t[129] & ~t[132]) | (t[126] & ~t[127] & t[130] & t[131] & ~t[132]) | (t[127] & ~t[129] & ~t[131] & t[132]) | (~t[127] & t[129] & t[131] & t[132]);
  assign t[123] = (t[126] & t[127] & t[128] & ~t[129] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[129] & ~t[130] & t[131] & t[132]) | (~t[127] & ~t[128] & t[129] & ~t[130] & ~t[131]) | (~t[126] & ~t[128] & t[129] & ~t[131] & ~t[132]) | (~t[126] & ~t[127] & t[129] & ~t[130] & ~t[132]) | (~t[127] & t[128] & t[129] & t[130] & ~t[131]) | (~t[128] & t[129] & t[130] & ~t[132]);
  assign t[124] = (t[126] & t[127] & ~t[128] & ~t[130] & t[131] & ~t[132]) | (t[126] & t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[132]) | (~t[126] & ~t[128] & ~t[129] & t[130] & ~t[131]) | (~t[126] & ~t[127] & ~t[129] & t[130] & ~t[132]) | (~t[126] & ~t[128] & t[129] & t[130] & t[131]) | (t[129] & t[130] & ~t[131] & ~t[132]);
  assign t[125] = (t[126] & t[127] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[128] & ~t[129] & ~t[130] & t[131]) | (~t[126] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[126] & ~t[127] & ~t[128] & t[131] & ~t[132]) | (~t[127] & t[128] & ~t[129] & t[130] & t[131]) | (t[128] & ~t[130] & t[131] & ~t[132]);
  assign t[126] = t[154] ^ x[7];
  assign t[127] = t[155] ^ x[43];
  assign t[128] = t[156] ^ x[8];
  assign t[129] = t[157] ^ x[44];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[45];
  assign t[131] = t[159] ^ x[46];
  assign t[132] = t[160] ^ x[6];
  assign t[133] = t[161] ^ x[14];
  assign t[134] = t[162] ^ x[31];
  assign t[135] = t[163] ^ x[15];
  assign t[136] = t[164] ^ x[32];
  assign t[137] = t[165] ^ x[30];
  assign t[138] = t[166] ^ x[33];
  assign t[139] = t[167] ^ x[13];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[168] ^ x[21];
  assign t[141] = t[169] ^ x[35];
  assign t[142] = t[170] ^ x[22];
  assign t[143] = t[171] ^ x[36];
  assign t[144] = t[172] ^ x[34];
  assign t[145] = t[173] ^ x[37];
  assign t[146] = t[174] ^ x[20];
  assign t[147] = t[175] ^ x[28];
  assign t[148] = t[176] ^ x[39];
  assign t[149] = t[177] ^ x[29];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[178] ^ x[40];
  assign t[151] = t[179] ^ x[38];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[27];
  assign t[154] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[155] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[156] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[157] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[158] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[159] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[161] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[162] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[163] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[164] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[165] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[166] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[167] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[168] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[169] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[171] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[172] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[173] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[174] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[175] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[176] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[177] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[178] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[179] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[17] = t[65] ^ t[28];
  assign t[180] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[181] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[66] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[67] ^ t[38];
  assign t[26] = t[68] ^ t[69];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[69]);
  assign t[29] = ~(t[65] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[64]);
  assign t[30] = t[65] & t[42];
  assign t[31] = t[70] ^ t[71];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[71]);
  assign t[34] = ~(t[66] ^ t[33]);
  assign t[35] = t[66] & t[44];
  assign t[36] = t[72] ^ t[73];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[73]);
  assign t[39] = ~(t[67] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[67] & t[46];
  assign t[41] = t[65] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[66] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[67] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[69] ^ t[74];
  assign t[48] = t[65] ^ t[26];
  assign t[49] = t[71] ^ t[75];
  assign t[4] = ~t[7];
  assign t[50] = t[66] ^ t[31];
  assign t[51] = t[73] ^ t[76];
  assign t[52] = t[67] ^ t[36];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[77]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[61]);
  assign t[59] = ~(t[62]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = ~(t[63]);
  assign t[61] = t[47] ^ t[15];
  assign t[62] = t[49] ^ t[19];
  assign t[63] = t[51] ^ t[23];
  assign t[64] = (t[78] & ~t[79]) | (~t[78] & t[79]);
  assign t[65] = (t[80] & ~t[81]) | (~t[80] & t[81]);
  assign t[66] = (t[82] & ~t[83]) | (~t[82] & t[83]);
  assign t[67] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[68] = (t[80] & ~t[86]) | (~t[80] & t[86]);
  assign t[69] = (t[80] & ~t[88] & ~t[89]) | (~t[87] & t[88] & ~t[86]) | (~t[80] & ~t[88] & t[89]) | (t[87] & t[88] & t[86]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (t[82] & ~t[90]) | (~t[82] & t[90]);
  assign t[71] = (t[82] & ~t[92] & ~t[93]) | (~t[91] & t[92] & ~t[90]) | (~t[82] & ~t[92] & t[93]) | (t[91] & t[92] & t[90]);
  assign t[72] = (t[84] & ~t[94]) | (~t[84] & t[94]);
  assign t[73] = (t[84] & ~t[96] & ~t[97]) | (~t[95] & t[96] & ~t[94]) | (~t[84] & ~t[96] & t[97]) | (t[95] & t[96] & t[94]);
  assign t[74] = (t[80] & ~t[88] & ~t[86]) | (~t[87] & t[88] & ~t[89]) | (~t[80] & ~t[88] & t[86]) | (t[87] & t[88] & t[89]);
  assign t[75] = (t[82] & ~t[92] & ~t[90]) | (~t[91] & t[92] & ~t[93]) | (~t[82] & ~t[92] & t[90]) | (t[91] & t[92] & t[93]);
  assign t[76] = (t[84] & ~t[96] & ~t[94]) | (~t[95] & t[96] & ~t[97]) | (~t[84] & ~t[96] & t[94]) | (t[95] & t[96] & t[97]);
  assign t[77] = (t[78] & ~t[99] & ~t[101]) | (~t[98] & t[99] & ~t[100]) | (~t[78] & ~t[99] & t[101]) | (t[98] & t[99] & t[100]);
  assign t[78] = t[102] ^ x[7];
  assign t[79] = t[103] ^ x[8];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[104] ^ x[14];
  assign t[81] = t[105] ^ x[15];
  assign t[82] = t[106] ^ x[21];
  assign t[83] = t[107] ^ x[22];
  assign t[84] = t[108] ^ x[28];
  assign t[85] = t[109] ^ x[29];
  assign t[86] = t[110] ^ x[30];
  assign t[87] = t[111] ^ x[31];
  assign t[88] = t[112] ^ x[32];
  assign t[89] = t[113] ^ x[33];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[114] ^ x[34];
  assign t[91] = t[115] ^ x[35];
  assign t[92] = t[116] ^ x[36];
  assign t[93] = t[117] ^ x[37];
  assign t[94] = t[118] ^ x[38];
  assign t[95] = t[119] ^ x[39];
  assign t[96] = t[120] ^ x[40];
  assign t[97] = t[121] ^ x[41];
  assign t[98] = t[122] ^ x[43];
  assign t[99] = t[123] ^ x[44];
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind159(x, y);
 input [46:0] x;
 output y;

 wire [178:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[123] & t[124] & ~t[125] & t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[125] & ~t[126] & t[127] & ~t[128] & t[129]) | (~t[124] & t[125] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[124] & t[125] & ~t[128] & ~t[129]) | (~t[123] & t[125] & t[126] & ~t[127] & t[128]) | (t[125] & ~t[126] & t[128] & ~t[129]);
  assign t[101] = (t[130] & ~t[132] & ~t[133] & ~t[134] & ~t[135]) | (t[130] & ~t[131] & ~t[133] & ~t[134] & ~t[136]) | (t[130] & ~t[131] & ~t[132] & ~t[135] & ~t[136]) | (~t[130] & t[131] & t[132] & t[133] & ~t[136]) | (~t[130] & t[131] & t[134] & t[135] & ~t[136]) | (t[130] & ~t[132] & ~t[134] & t[136]) | (~t[130] & t[132] & t[134] & t[136]);
  assign t[102] = (t[130] & t[131] & ~t[132] & t[133] & ~t[134] & ~t[136]) | (t[130] & ~t[132] & ~t[133] & t[134] & ~t[135] & t[136]) | (~t[131] & t[132] & ~t[133] & ~t[134] & ~t[136]) | (~t[130] & t[132] & ~t[133] & ~t[134] & ~t[135]) | (~t[130] & ~t[131] & t[132] & ~t[135] & ~t[136]) | (~t[130] & t[132] & t[133] & ~t[134] & t[135]) | (t[132] & ~t[133] & t[135] & ~t[136]);
  assign t[103] = (t[137] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & ~t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[138] & ~t[139] & ~t[142] & ~t[143]) | (~t[137] & t[138] & t[139] & t[140] & ~t[143]) | (~t[137] & t[138] & t[141] & t[142] & ~t[143]) | (t[137] & ~t[139] & ~t[141] & t[143]) | (~t[137] & t[139] & t[141] & t[143]);
  assign t[104] = (t[137] & t[138] & ~t[139] & t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[139] & ~t[140] & t[141] & ~t[142] & t[143]) | (~t[138] & t[139] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[138] & t[139] & ~t[142] & ~t[143]) | (~t[137] & t[139] & t[140] & ~t[141] & t[142]) | (t[139] & ~t[140] & t[142] & ~t[143]);
  assign t[105] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[106] = (t[144] & t[145] & ~t[146] & t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[146] & ~t[147] & t[148] & ~t[149] & t[150]) | (~t[145] & t[146] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[145] & t[146] & ~t[149] & ~t[150]) | (~t[144] & t[146] & t[147] & ~t[148] & t[149]) | (t[146] & ~t[147] & t[149] & ~t[150]);
  assign t[107] = (t[130] & t[131] & ~t[132] & ~t[134] & t[135] & ~t[136]) | (t[130] & t[132] & ~t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[132] & t[134] & ~t[135] & ~t[136]) | (~t[130] & ~t[132] & ~t[133] & t[134] & ~t[135]) | (~t[130] & ~t[131] & ~t[133] & t[134] & ~t[136]) | (~t[130] & ~t[132] & t[133] & t[134] & t[135]) | (t[133] & t[134] & ~t[135] & ~t[136]);
  assign t[108] = (t[131] & ~t[132] & ~t[133] & ~t[134] & ~t[135]) | (~t[130] & t[131] & ~t[133] & ~t[134] & ~t[136]) | (~t[130] & t[131] & ~t[132] & ~t[135] & ~t[136]) | (t[130] & ~t[131] & t[132] & t[133] & ~t[136]) | (t[130] & ~t[131] & t[134] & t[135] & ~t[136]) | (t[131] & ~t[133] & ~t[135] & t[136]) | (~t[131] & t[133] & t[135] & t[136]);
  assign t[109] = (t[130] & t[131] & t[132] & ~t[133] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & ~t[133] & ~t[134] & t[135] & t[136]) | (~t[131] & ~t[132] & t[133] & ~t[134] & ~t[135]) | (~t[130] & ~t[132] & t[133] & ~t[135] & ~t[136]) | (~t[130] & ~t[131] & t[133] & ~t[134] & ~t[136]) | (~t[131] & t[132] & t[133] & t[134] & ~t[135]) | (~t[132] & t[133] & t[134] & ~t[136]);
  assign t[10] = t[18] ^ t[19];
  assign t[110] = (t[130] & t[131] & ~t[133] & t[134] & ~t[135] & ~t[136]) | (t[131] & ~t[132] & t[133] & ~t[134] & ~t[135] & t[136]) | (~t[131] & ~t[132] & ~t[133] & ~t[134] & t[135]) | (~t[130] & ~t[133] & ~t[134] & t[135] & ~t[136]) | (~t[130] & ~t[131] & ~t[132] & t[135] & ~t[136]) | (~t[131] & t[132] & ~t[133] & t[134] & t[135]) | (t[132] & ~t[134] & t[135] & ~t[136]);
  assign t[111] = (t[137] & t[138] & ~t[139] & ~t[141] & t[142] & ~t[143]) | (t[137] & t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[143]) | (~t[137] & ~t[139] & ~t[140] & t[141] & ~t[142]) | (~t[137] & ~t[138] & ~t[140] & t[141] & ~t[143]) | (~t[137] & ~t[139] & t[140] & t[141] & t[142]) | (t[140] & t[141] & ~t[142] & ~t[143]);
  assign t[112] = (t[138] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & t[138] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[138] & ~t[139] & ~t[142] & ~t[143]) | (t[137] & ~t[138] & t[139] & t[140] & ~t[143]) | (t[137] & ~t[138] & t[141] & t[142] & ~t[143]) | (t[138] & ~t[140] & ~t[142] & t[143]) | (~t[138] & t[140] & t[142] & t[143]);
  assign t[113] = (t[137] & t[138] & t[139] & ~t[140] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[140] & ~t[141] & t[142] & t[143]) | (~t[138] & ~t[139] & t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[139] & t[140] & ~t[142] & ~t[143]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[143]) | (~t[138] & t[139] & t[140] & t[141] & ~t[142]) | (~t[139] & t[140] & t[141] & ~t[143]);
  assign t[114] = (t[137] & t[138] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[137] & ~t[138] & ~t[139] & t[142] & ~t[143]) | (~t[138] & t[139] & ~t[140] & t[141] & t[142]) | (t[139] & ~t[141] & t[142] & ~t[143]);
  assign t[115] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[116] = (t[145] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (~t[144] & t[145] & ~t[147] & ~t[148] & ~t[150]) | (~t[144] & t[145] & ~t[146] & ~t[149] & ~t[150]) | (t[144] & ~t[145] & t[146] & t[147] & ~t[150]) | (t[144] & ~t[145] & t[148] & t[149] & ~t[150]) | (t[145] & ~t[147] & ~t[149] & t[150]) | (~t[145] & t[147] & t[149] & t[150]);
  assign t[117] = (t[144] & t[145] & t[146] & ~t[147] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[147] & ~t[148] & t[149] & t[150]) | (~t[145] & ~t[146] & t[147] & ~t[148] & ~t[149]) | (~t[144] & ~t[146] & t[147] & ~t[149] & ~t[150]) | (~t[144] & ~t[145] & t[147] & ~t[148] & ~t[150]) | (~t[145] & t[146] & t[147] & t[148] & ~t[149]) | (~t[146] & t[147] & t[148] & ~t[150]);
  assign t[118] = (t[144] & t[145] & ~t[147] & t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & ~t[147] & ~t[148] & t[149]) | (~t[144] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[144] & ~t[145] & ~t[146] & t[149] & ~t[150]) | (~t[145] & t[146] & ~t[147] & t[148] & t[149]) | (t[146] & ~t[148] & t[149] & ~t[150]);
  assign t[119] = (t[124] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (~t[123] & t[124] & ~t[126] & ~t[127] & ~t[129]) | (~t[123] & t[124] & ~t[125] & ~t[128] & ~t[129]) | (t[123] & ~t[124] & t[125] & t[126] & ~t[129]) | (t[123] & ~t[124] & t[127] & t[128] & ~t[129]) | (t[124] & ~t[126] & ~t[128] & t[129]) | (~t[124] & t[126] & t[128] & t[129]);
  assign t[11] = t[20] ^ t[21];
  assign t[120] = (t[123] & t[124] & t[125] & ~t[126] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & ~t[126] & ~t[127] & t[128] & t[129]) | (~t[124] & ~t[125] & t[126] & ~t[127] & ~t[128]) | (~t[123] & ~t[125] & t[126] & ~t[128] & ~t[129]) | (~t[123] & ~t[124] & t[126] & ~t[127] & ~t[129]) | (~t[124] & t[125] & t[126] & t[127] & ~t[128]) | (~t[125] & t[126] & t[127] & ~t[129]);
  assign t[121] = (t[123] & t[124] & ~t[125] & ~t[127] & t[128] & ~t[129]) | (t[123] & t[125] & ~t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & t[127] & ~t[128] & ~t[129]) | (~t[123] & ~t[125] & ~t[126] & t[127] & ~t[128]) | (~t[123] & ~t[124] & ~t[126] & t[127] & ~t[129]) | (~t[123] & ~t[125] & t[126] & t[127] & t[128]) | (t[126] & t[127] & ~t[128] & ~t[129]);
  assign t[122] = (t[123] & t[124] & ~t[126] & t[127] & ~t[128] & ~t[129]) | (t[124] & ~t[125] & t[126] & ~t[127] & ~t[128] & t[129]) | (~t[124] & ~t[125] & ~t[126] & ~t[127] & t[128]) | (~t[123] & ~t[126] & ~t[127] & t[128] & ~t[129]) | (~t[123] & ~t[124] & ~t[125] & t[128] & ~t[129]) | (~t[124] & t[125] & ~t[126] & t[127] & t[128]) | (t[125] & ~t[127] & t[128] & ~t[129]);
  assign t[123] = t[151] ^ x[7];
  assign t[124] = t[152] ^ x[43];
  assign t[125] = t[153] ^ x[8];
  assign t[126] = t[154] ^ x[44];
  assign t[127] = t[155] ^ x[45];
  assign t[128] = t[156] ^ x[46];
  assign t[129] = t[157] ^ x[6];
  assign t[12] = t[22] ^ t[23];
  assign t[130] = t[158] ^ x[14];
  assign t[131] = t[159] ^ x[31];
  assign t[132] = t[160] ^ x[15];
  assign t[133] = t[161] ^ x[32];
  assign t[134] = t[162] ^ x[30];
  assign t[135] = t[163] ^ x[33];
  assign t[136] = t[164] ^ x[13];
  assign t[137] = t[165] ^ x[21];
  assign t[138] = t[166] ^ x[35];
  assign t[139] = t[167] ^ x[22];
  assign t[13] = t[24] ^ t[25];
  assign t[140] = t[168] ^ x[36];
  assign t[141] = t[169] ^ x[34];
  assign t[142] = t[170] ^ x[37];
  assign t[143] = t[171] ^ x[20];
  assign t[144] = t[172] ^ x[28];
  assign t[145] = t[173] ^ x[39];
  assign t[146] = t[174] ^ x[29];
  assign t[147] = t[175] ^ x[40];
  assign t[148] = t[176] ^ x[38];
  assign t[149] = t[177] ^ x[41];
  assign t[14] = t[26] ^ t[27];
  assign t[150] = t[178] ^ x[27];
  assign t[151] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[152] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[153] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[154] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[155] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[156] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[157] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[158] = (x[9] & ~x[10] & ~x[11]) | (~x[9] & x[10] & ~x[11]) | (~x[9] & ~x[10] & x[11]) | (x[9] & x[10] & x[11]);
  assign t[159] = (x[9] & ~x[10] & ~x[12]) | (~x[9] & x[10] & ~x[12]) | (~x[9] & ~x[10] & x[12]) | (x[9] & x[10] & x[12]);
  assign t[15] = t[28] & t[29];
  assign t[160] = (x[9] & ~x[11]) | (~x[9] & x[11]);
  assign t[161] = (x[9] & ~x[12]) | (~x[9] & x[12]);
  assign t[162] = (x[10] & ~x[11]) | (~x[10] & x[11]);
  assign t[163] = (x[10] & ~x[12]) | (~x[10] & x[12]);
  assign t[164] = (x[11] & ~x[12]) | (~x[11] & x[12]);
  assign t[165] = (x[16] & ~x[17] & ~x[18]) | (~x[16] & x[17] & ~x[18]) | (~x[16] & ~x[17] & x[18]) | (x[16] & x[17] & x[18]);
  assign t[166] = (x[16] & ~x[17] & ~x[19]) | (~x[16] & x[17] & ~x[19]) | (~x[16] & ~x[17] & x[19]) | (x[16] & x[17] & x[19]);
  assign t[167] = (x[16] & ~x[18]) | (~x[16] & x[18]);
  assign t[168] = (x[16] & ~x[19]) | (~x[16] & x[19]);
  assign t[169] = (x[17] & ~x[18]) | (~x[17] & x[18]);
  assign t[16] = t[30] ^ t[15];
  assign t[170] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[171] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[172] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[173] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[174] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[175] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[176] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[177] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[178] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[17] = t[62] ^ t[28];
  assign t[18] = t[31] ^ t[32];
  assign t[19] = t[33] & t[34];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[35] ^ t[19];
  assign t[21] = t[63] ^ t[33];
  assign t[22] = t[36] ^ t[37];
  assign t[23] = t[38] & t[39];
  assign t[24] = t[40] ^ t[23];
  assign t[25] = t[64] ^ t[38];
  assign t[26] = t[65] ^ t[66];
  assign t[27] = t[28] & t[41];
  assign t[28] = ~(t[66]);
  assign t[29] = ~(t[62] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[61]);
  assign t[30] = t[62] & t[42];
  assign t[31] = t[67] ^ t[68];
  assign t[32] = t[33] & t[43];
  assign t[33] = ~(t[68]);
  assign t[34] = ~(t[63] ^ t[33]);
  assign t[35] = t[63] & t[44];
  assign t[36] = t[69] ^ t[70];
  assign t[37] = t[38] & t[45];
  assign t[38] = ~(t[70]);
  assign t[39] = ~(t[64] ^ t[38]);
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[64] & t[46];
  assign t[41] = t[62] ^ t[47];
  assign t[42] = t[48] ^ t[27];
  assign t[43] = t[63] ^ t[49];
  assign t[44] = t[50] ^ t[32];
  assign t[45] = t[64] ^ t[51];
  assign t[46] = t[52] ^ t[37];
  assign t[47] = t[66] ^ t[71];
  assign t[48] = t[62] ^ t[26];
  assign t[49] = t[68] ^ t[72];
  assign t[4] = ~t[7];
  assign t[50] = t[63] ^ t[31];
  assign t[51] = t[70] ^ t[73];
  assign t[52] = t[64] ^ t[36];
  assign t[53] = x[0] ? x[42] : t[54];
  assign t[54] = ~(t[55] ^ t[56]);
  assign t[55] = ~(t[57] ^ t[74]);
  assign t[56] = ~(t[58] ^ t[59]);
  assign t[57] = ~t[60];
  assign t[58] = ~(t[8]);
  assign t[59] = ~(t[10]);
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = ~(t[12]);
  assign t[61] = (t[75] & ~t[76]) | (~t[75] & t[76]);
  assign t[62] = (t[77] & ~t[78]) | (~t[77] & t[78]);
  assign t[63] = (t[79] & ~t[80]) | (~t[79] & t[80]);
  assign t[64] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[65] = (t[77] & ~t[83]) | (~t[77] & t[83]);
  assign t[66] = (t[77] & ~t[85] & ~t[86]) | (~t[84] & t[85] & ~t[83]) | (~t[77] & ~t[85] & t[86]) | (t[84] & t[85] & t[83]);
  assign t[67] = (t[79] & ~t[87]) | (~t[79] & t[87]);
  assign t[68] = (t[79] & ~t[89] & ~t[90]) | (~t[88] & t[89] & ~t[87]) | (~t[79] & ~t[89] & t[90]) | (t[88] & t[89] & t[87]);
  assign t[69] = (t[81] & ~t[91]) | (~t[81] & t[91]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (t[81] & ~t[93] & ~t[94]) | (~t[92] & t[93] & ~t[91]) | (~t[81] & ~t[93] & t[94]) | (t[92] & t[93] & t[91]);
  assign t[71] = (t[77] & ~t[85] & ~t[83]) | (~t[84] & t[85] & ~t[86]) | (~t[77] & ~t[85] & t[83]) | (t[84] & t[85] & t[86]);
  assign t[72] = (t[79] & ~t[89] & ~t[87]) | (~t[88] & t[89] & ~t[90]) | (~t[79] & ~t[89] & t[87]) | (t[88] & t[89] & t[90]);
  assign t[73] = (t[81] & ~t[93] & ~t[91]) | (~t[92] & t[93] & ~t[94]) | (~t[81] & ~t[93] & t[91]) | (t[92] & t[93] & t[94]);
  assign t[74] = (t[75] & ~t[96] & ~t[97]) | (~t[95] & t[96] & ~t[98]) | (~t[75] & ~t[96] & t[97]) | (t[95] & t[96] & t[98]);
  assign t[75] = t[99] ^ x[7];
  assign t[76] = t[100] ^ x[8];
  assign t[77] = t[101] ^ x[14];
  assign t[78] = t[102] ^ x[15];
  assign t[79] = t[103] ^ x[21];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[104] ^ x[22];
  assign t[81] = t[105] ^ x[28];
  assign t[82] = t[106] ^ x[29];
  assign t[83] = t[107] ^ x[30];
  assign t[84] = t[108] ^ x[31];
  assign t[85] = t[109] ^ x[32];
  assign t[86] = t[110] ^ x[33];
  assign t[87] = t[111] ^ x[34];
  assign t[88] = t[112] ^ x[35];
  assign t[89] = t[113] ^ x[36];
  assign t[8] = t[14] ^ t[15];
  assign t[90] = t[114] ^ x[37];
  assign t[91] = t[115] ^ x[38];
  assign t[92] = t[116] ^ x[39];
  assign t[93] = t[117] ^ x[40];
  assign t[94] = t[118] ^ x[41];
  assign t[95] = t[119] ^ x[43];
  assign t[96] = t[120] ^ x[44];
  assign t[97] = t[121] ^ x[45];
  assign t[98] = t[122] ^ x[46];
  assign t[99] = (t[123] & ~t[125] & ~t[126] & ~t[127] & ~t[128]) | (t[123] & ~t[124] & ~t[126] & ~t[127] & ~t[129]) | (t[123] & ~t[124] & ~t[125] & ~t[128] & ~t[129]) | (~t[123] & t[124] & t[125] & t[126] & ~t[129]) | (~t[123] & t[124] & t[127] & t[128] & ~t[129]) | (t[123] & ~t[125] & ~t[127] & t[129]) | (~t[123] & t[125] & t[127] & t[129]);
  assign t[9] = t[16] ^ t[17];
  assign y = (t[0] & ~t[53]) | (~t[0] & t[53]);
endmodule

module R2ind160(x, y);
 input [46:0] x;
 output y;

 wire [161:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[127] & t[128] & t[129] & ~t[130] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & ~t[130] & ~t[131] & t[132] & t[133]) | (~t[128] & ~t[129] & t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[129] & t[130] & ~t[132] & ~t[133]) | (~t[127] & ~t[128] & t[130] & ~t[131] & ~t[133]) | (~t[128] & t[129] & t[130] & t[131] & ~t[132]) | (~t[129] & t[130] & t[131] & ~t[133]);
  assign t[101] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[102] = (t[127] & t[128] & ~t[130] & t[131] & ~t[132] & ~t[133]) | (t[128] & ~t[129] & t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & ~t[130] & ~t[131] & t[132]) | (~t[127] & ~t[130] & ~t[131] & t[132] & ~t[133]) | (~t[127] & ~t[128] & ~t[129] & t[132] & ~t[133]) | (~t[128] & t[129] & ~t[130] & t[131] & t[132]) | (t[129] & ~t[131] & t[132] & ~t[133]);
  assign t[103] = (t[113] & t[114] & ~t[115] & t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[115] & ~t[116] & t[117] & ~t[118] & t[119]) | (~t[114] & t[115] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[114] & t[115] & ~t[118] & ~t[119]) | (~t[113] & t[115] & t[116] & ~t[117] & t[118]) | (t[115] & ~t[116] & t[118] & ~t[119]);
  assign t[104] = (t[120] & t[121] & ~t[122] & t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[122] & ~t[123] & t[124] & ~t[125] & t[126]) | (~t[121] & t[122] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[121] & t[122] & ~t[125] & ~t[126]) | (~t[120] & t[122] & t[123] & ~t[124] & t[125]) | (t[122] & ~t[123] & t[125] & ~t[126]);
  assign t[105] = (t[127] & t[128] & ~t[129] & t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[129] & ~t[130] & t[131] & ~t[132] & t[133]) | (~t[128] & t[129] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & ~t[128] & t[129] & ~t[132] & ~t[133]) | (~t[127] & t[129] & t[130] & ~t[131] & t[132]) | (t[129] & ~t[130] & t[132] & ~t[133]);
  assign t[106] = t[134] ^ x[8];
  assign t[107] = t[135] ^ x[9];
  assign t[108] = t[136] ^ x[6];
  assign t[109] = t[137] ^ x[10];
  assign t[10] = t[15] ^ t[16];
  assign t[110] = t[138] ^ x[11];
  assign t[111] = t[139] ^ x[12];
  assign t[112] = t[140] ^ x[7];
  assign t[113] = t[141] ^ x[18];
  assign t[114] = t[142] ^ x[19];
  assign t[115] = t[143] ^ x[43];
  assign t[116] = t[144] ^ x[20];
  assign t[117] = t[145] ^ x[21];
  assign t[118] = t[146] ^ x[22];
  assign t[119] = t[147] ^ x[17];
  assign t[11] = t[47] ^ t[48];
  assign t[120] = t[148] ^ x[28];
  assign t[121] = t[149] ^ x[29];
  assign t[122] = t[150] ^ x[44];
  assign t[123] = t[151] ^ x[30];
  assign t[124] = t[152] ^ x[31];
  assign t[125] = t[153] ^ x[32];
  assign t[126] = t[154] ^ x[27];
  assign t[127] = t[155] ^ x[38];
  assign t[128] = t[156] ^ x[39];
  assign t[129] = t[157] ^ x[45];
  assign t[12] = t[17] & t[18];
  assign t[130] = t[158] ^ x[40];
  assign t[131] = t[159] ^ x[41];
  assign t[132] = t[160] ^ x[42];
  assign t[133] = t[161] ^ x[37];
  assign t[134] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[135] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[136] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[137] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[138] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[139] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[13] = t[49] ^ t[50];
  assign t[140] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[141] = (x[13] & ~x[14] & ~x[15]) | (~x[13] & x[14] & ~x[15]) | (~x[13] & ~x[14] & x[15]) | (x[13] & x[14] & x[15]);
  assign t[142] = (x[13] & ~x[14] & ~x[16]) | (~x[13] & x[14] & ~x[16]) | (~x[13] & ~x[14] & x[16]) | (x[13] & x[14] & x[16]);
  assign t[143] = (x[13] & ~x[15]) | (~x[13] & x[15]);
  assign t[144] = (x[13] & ~x[16]) | (~x[13] & x[16]);
  assign t[145] = (x[14] & ~x[15]) | (~x[14] & x[15]);
  assign t[146] = (x[14] & ~x[16]) | (~x[14] & x[16]);
  assign t[147] = (x[15] & ~x[16]) | (~x[15] & x[16]);
  assign t[148] = (x[23] & ~x[24] & ~x[25]) | (~x[23] & x[24] & ~x[25]) | (~x[23] & ~x[24] & x[25]) | (x[23] & x[24] & x[25]);
  assign t[149] = (x[23] & ~x[24] & ~x[26]) | (~x[23] & x[24] & ~x[26]) | (~x[23] & ~x[24] & x[26]) | (x[23] & x[24] & x[26]);
  assign t[14] = t[19] & t[20];
  assign t[150] = (x[23] & ~x[25]) | (~x[23] & x[25]);
  assign t[151] = (x[23] & ~x[26]) | (~x[23] & x[26]);
  assign t[152] = (x[24] & ~x[25]) | (~x[24] & x[25]);
  assign t[153] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[154] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[155] = (x[33] & ~x[34] & ~x[35]) | (~x[33] & x[34] & ~x[35]) | (~x[33] & ~x[34] & x[35]) | (x[33] & x[34] & x[35]);
  assign t[156] = (x[33] & ~x[34] & ~x[36]) | (~x[33] & x[34] & ~x[36]) | (~x[33] & ~x[34] & x[36]) | (x[33] & x[34] & x[36]);
  assign t[157] = (x[33] & ~x[35]) | (~x[33] & x[35]);
  assign t[158] = (x[33] & ~x[36]) | (~x[33] & x[36]);
  assign t[159] = (x[34] & ~x[35]) | (~x[34] & x[35]);
  assign t[15] = t[51] ^ t[52];
  assign t[160] = (x[34] & ~x[36]) | (~x[34] & x[36]);
  assign t[161] = (x[35] & ~x[36]) | (~x[35] & x[36]);
  assign t[16] = t[21] & t[22];
  assign t[17] = ~(t[47]);
  assign t[18] = ~(t[53] ^ t[17]);
  assign t[19] = ~(t[49]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[54] ^ t[19]);
  assign t[21] = ~(t[51]);
  assign t[22] = ~(t[55] ^ t[21]);
  assign t[23] = x[0] ? x[46] : t[24];
  assign t[24] = ~(t[25] ^ t[26]);
  assign t[25] = ~(t[27] ^ t[56]);
  assign t[26] = ~(t[28] ^ t[29]);
  assign t[27] = ~t[30];
  assign t[28] = ~(t[31]);
  assign t[29] = ~(t[32]);
  assign t[2] = ~(t[4] ^ t[46]);
  assign t[30] = ~(t[33]);
  assign t[31] = t[34] ^ t[12];
  assign t[32] = t[35] ^ t[14];
  assign t[33] = t[36] ^ t[16];
  assign t[34] = t[37] ^ t[38];
  assign t[35] = t[39] ^ t[40];
  assign t[36] = t[41] ^ t[42];
  assign t[37] = t[57] ^ t[47];
  assign t[38] = t[17] & t[43];
  assign t[39] = t[58] ^ t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[19] & t[44];
  assign t[41] = t[59] ^ t[51];
  assign t[42] = t[21] & t[45];
  assign t[43] = t[53] ^ t[11];
  assign t[44] = t[54] ^ t[13];
  assign t[45] = t[55] ^ t[15];
  assign t[46] = (t[60] & ~t[62] & ~t[64]) | (~t[61] & t[62] & ~t[63]) | (~t[60] & ~t[62] & t[64]) | (t[61] & t[62] & t[63]);
  assign t[47] = (t[65] & ~t[67] & ~t[69]) | (~t[66] & t[67] & ~t[68]) | (~t[65] & ~t[67] & t[69]) | (t[66] & t[67] & t[68]);
  assign t[48] = (t[65] & ~t[67] & ~t[68]) | (~t[66] & t[67] & ~t[69]) | (~t[65] & ~t[67] & t[68]) | (t[66] & t[67] & t[69]);
  assign t[49] = (t[70] & ~t[72] & ~t[74]) | (~t[71] & t[72] & ~t[73]) | (~t[70] & ~t[72] & t[74]) | (t[71] & t[72] & t[73]);
  assign t[4] = ~t[7];
  assign t[50] = (t[70] & ~t[72] & ~t[73]) | (~t[71] & t[72] & ~t[74]) | (~t[70] & ~t[72] & t[73]) | (t[71] & t[72] & t[74]);
  assign t[51] = (t[75] & ~t[77] & ~t[79]) | (~t[76] & t[77] & ~t[78]) | (~t[75] & ~t[77] & t[79]) | (t[76] & t[77] & t[78]);
  assign t[52] = (t[75] & ~t[77] & ~t[78]) | (~t[76] & t[77] & ~t[79]) | (~t[75] & ~t[77] & t[78]) | (t[76] & t[77] & t[79]);
  assign t[53] = (t[65] & ~t[80]) | (~t[65] & t[80]);
  assign t[54] = (t[70] & ~t[81]) | (~t[70] & t[81]);
  assign t[55] = (t[75] & ~t[82]) | (~t[75] & t[82]);
  assign t[56] = (t[60] & ~t[62] & ~t[63]) | (~t[61] & t[62] & ~t[64]) | (~t[60] & ~t[62] & t[63]) | (t[61] & t[62] & t[64]);
  assign t[57] = (t[65] & ~t[68]) | (~t[65] & t[68]);
  assign t[58] = (t[70] & ~t[73]) | (~t[70] & t[73]);
  assign t[59] = (t[75] & ~t[78]) | (~t[75] & t[78]);
  assign t[5] = ~(t[8]);
  assign t[60] = t[83] ^ x[8];
  assign t[61] = t[84] ^ x[9];
  assign t[62] = t[85] ^ x[10];
  assign t[63] = t[86] ^ x[11];
  assign t[64] = t[87] ^ x[12];
  assign t[65] = t[88] ^ x[18];
  assign t[66] = t[89] ^ x[19];
  assign t[67] = t[90] ^ x[20];
  assign t[68] = t[91] ^ x[21];
  assign t[69] = t[92] ^ x[22];
  assign t[6] = ~(t[9]);
  assign t[70] = t[93] ^ x[28];
  assign t[71] = t[94] ^ x[29];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[31];
  assign t[74] = t[97] ^ x[32];
  assign t[75] = t[98] ^ x[38];
  assign t[76] = t[99] ^ x[39];
  assign t[77] = t[100] ^ x[40];
  assign t[78] = t[101] ^ x[41];
  assign t[79] = t[102] ^ x[42];
  assign t[7] = ~(t[10]);
  assign t[80] = t[103] ^ x[43];
  assign t[81] = t[104] ^ x[44];
  assign t[82] = t[105] ^ x[45];
  assign t[83] = (t[106] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (t[106] & ~t[107] & ~t[109] & ~t[110] & ~t[112]) | (t[106] & ~t[107] & ~t[108] & ~t[111] & ~t[112]) | (~t[106] & t[107] & t[108] & t[109] & ~t[112]) | (~t[106] & t[107] & t[110] & t[111] & ~t[112]) | (t[106] & ~t[108] & ~t[110] & t[112]) | (~t[106] & t[108] & t[110] & t[112]);
  assign t[84] = (t[107] & ~t[108] & ~t[109] & ~t[110] & ~t[111]) | (~t[106] & t[107] & ~t[109] & ~t[110] & ~t[112]) | (~t[106] & t[107] & ~t[108] & ~t[111] & ~t[112]) | (t[106] & ~t[107] & t[108] & t[109] & ~t[112]) | (t[106] & ~t[107] & t[110] & t[111] & ~t[112]) | (t[107] & ~t[109] & ~t[111] & t[112]) | (~t[107] & t[109] & t[111] & t[112]);
  assign t[85] = (t[106] & t[107] & t[108] & ~t[109] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & ~t[109] & ~t[110] & t[111] & t[112]) | (~t[107] & ~t[108] & t[109] & ~t[110] & ~t[111]) | (~t[106] & ~t[108] & t[109] & ~t[111] & ~t[112]) | (~t[106] & ~t[107] & t[109] & ~t[110] & ~t[112]) | (~t[107] & t[108] & t[109] & t[110] & ~t[111]) | (~t[108] & t[109] & t[110] & ~t[112]);
  assign t[86] = (t[106] & t[107] & ~t[108] & ~t[110] & t[111] & ~t[112]) | (t[106] & t[108] & ~t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & t[110] & ~t[111] & ~t[112]) | (~t[106] & ~t[108] & ~t[109] & t[110] & ~t[111]) | (~t[106] & ~t[107] & ~t[109] & t[110] & ~t[112]) | (~t[106] & ~t[108] & t[109] & t[110] & t[111]) | (t[109] & t[110] & ~t[111] & ~t[112]);
  assign t[87] = (t[106] & t[107] & ~t[109] & t[110] & ~t[111] & ~t[112]) | (t[107] & ~t[108] & t[109] & ~t[110] & ~t[111] & t[112]) | (~t[107] & ~t[108] & ~t[109] & ~t[110] & t[111]) | (~t[106] & ~t[109] & ~t[110] & t[111] & ~t[112]) | (~t[106] & ~t[107] & ~t[108] & t[111] & ~t[112]) | (~t[107] & t[108] & ~t[109] & t[110] & t[111]) | (t[108] & ~t[110] & t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (t[113] & ~t[114] & ~t[116] & ~t[117] & ~t[119]) | (t[113] & ~t[114] & ~t[115] & ~t[118] & ~t[119]) | (~t[113] & t[114] & t[115] & t[116] & ~t[119]) | (~t[113] & t[114] & t[117] & t[118] & ~t[119]) | (t[113] & ~t[115] & ~t[117] & t[119]) | (~t[113] & t[115] & t[117] & t[119]);
  assign t[89] = (t[114] & ~t[115] & ~t[116] & ~t[117] & ~t[118]) | (~t[113] & t[114] & ~t[116] & ~t[117] & ~t[119]) | (~t[113] & t[114] & ~t[115] & ~t[118] & ~t[119]) | (t[113] & ~t[114] & t[115] & t[116] & ~t[119]) | (t[113] & ~t[114] & t[117] & t[118] & ~t[119]) | (t[114] & ~t[116] & ~t[118] & t[119]) | (~t[114] & t[116] & t[118] & t[119]);
  assign t[8] = t[11] ^ t[12];
  assign t[90] = (t[113] & t[114] & t[115] & ~t[116] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & ~t[116] & ~t[117] & t[118] & t[119]) | (~t[114] & ~t[115] & t[116] & ~t[117] & ~t[118]) | (~t[113] & ~t[115] & t[116] & ~t[118] & ~t[119]) | (~t[113] & ~t[114] & t[116] & ~t[117] & ~t[119]) | (~t[114] & t[115] & t[116] & t[117] & ~t[118]) | (~t[115] & t[116] & t[117] & ~t[119]);
  assign t[91] = (t[113] & t[114] & ~t[115] & ~t[117] & t[118] & ~t[119]) | (t[113] & t[115] & ~t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & t[117] & ~t[118] & ~t[119]) | (~t[113] & ~t[115] & ~t[116] & t[117] & ~t[118]) | (~t[113] & ~t[114] & ~t[116] & t[117] & ~t[119]) | (~t[113] & ~t[115] & t[116] & t[117] & t[118]) | (t[116] & t[117] & ~t[118] & ~t[119]);
  assign t[92] = (t[113] & t[114] & ~t[116] & t[117] & ~t[118] & ~t[119]) | (t[114] & ~t[115] & t[116] & ~t[117] & ~t[118] & t[119]) | (~t[114] & ~t[115] & ~t[116] & ~t[117] & t[118]) | (~t[113] & ~t[116] & ~t[117] & t[118] & ~t[119]) | (~t[113] & ~t[114] & ~t[115] & t[118] & ~t[119]) | (~t[114] & t[115] & ~t[116] & t[117] & t[118]) | (t[115] & ~t[117] & t[118] & ~t[119]);
  assign t[93] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[94] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[95] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[97] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[98] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[99] = (t[128] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (~t[127] & t[128] & ~t[130] & ~t[131] & ~t[133]) | (~t[127] & t[128] & ~t[129] & ~t[132] & ~t[133]) | (t[127] & ~t[128] & t[129] & t[130] & ~t[133]) | (t[127] & ~t[128] & t[131] & t[132] & ~t[133]) | (t[128] & ~t[130] & ~t[132] & t[133]) | (~t[128] & t[130] & t[132] & t[133]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0] & ~t[23]) | (~t[0] & t[23]);
endmodule

module R2ind161(x, y);
 input [71:0] x;
 output y;

 wire [265:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[114] & ~t[121] & ~t[122]) | (~t[120] & t[121] & ~t[123]) | (~t[114] & ~t[121] & t[122]) | (t[120] & t[121] & t[123]);
  assign t[101] = (t[124] & ~t[127] & ~t[129]) | (~t[126] & t[127] & ~t[128]) | (~t[124] & ~t[127] & t[129]) | (t[126] & t[127] & t[128]);
  assign t[102] = (t[124] & ~t[128]) | (~t[124] & t[128]);
  assign t[103] = (t[124] & ~t[127] & ~t[128]) | (~t[126] & t[127] & ~t[129]) | (~t[124] & ~t[127] & t[128]) | (t[126] & t[127] & t[129]);
  assign t[104] = (t[108] & ~t[130]) | (~t[108] & t[130]);
  assign t[105] = (t[131] & ~t[132]) | (~t[131] & t[132]);
  assign t[106] = (t[108] & ~t[134] & ~t[135]) | (~t[133] & t[134] & ~t[109]) | (~t[108] & ~t[134] & t[135]) | (t[133] & t[134] & t[109]);
  assign t[107] = (t[136] & ~t[137]) | (~t[136] & t[137]);
  assign t[108] = t[138] ^ x[7];
  assign t[109] = t[139] ^ x[8];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[140] ^ x[15];
  assign t[111] = t[141] ^ x[16];
  assign t[112] = t[142] ^ x[22];
  assign t[113] = t[143] ^ x[23];
  assign t[114] = t[144] ^ x[29];
  assign t[115] = t[145] ^ x[30];
  assign t[116] = t[146] ^ x[31];
  assign t[117] = t[147] ^ x[32];
  assign t[118] = t[148] ^ x[33];
  assign t[119] = t[149] ^ x[34];
  assign t[11] = t[19] & t[20];
  assign t[120] = t[150] ^ x[35];
  assign t[121] = t[151] ^ x[36];
  assign t[122] = t[152] ^ x[37];
  assign t[123] = t[153] ^ x[38];
  assign t[124] = t[154] ^ x[44];
  assign t[125] = t[155] ^ x[45];
  assign t[126] = t[156] ^ x[46];
  assign t[127] = t[157] ^ x[47];
  assign t[128] = t[158] ^ x[48];
  assign t[129] = t[159] ^ x[49];
  assign t[12] = ~t[21];
  assign t[130] = t[160] ^ x[51];
  assign t[131] = t[161] ^ x[58];
  assign t[132] = t[162] ^ x[59];
  assign t[133] = t[163] ^ x[61];
  assign t[134] = t[164] ^ x[62];
  assign t[135] = t[165] ^ x[63];
  assign t[136] = t[166] ^ x[70];
  assign t[137] = t[167] ^ x[71];
  assign t[138] = (t[168] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (t[168] & ~t[169] & ~t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[169] & ~t[170] & ~t[173] & ~t[174]) | (~t[168] & t[169] & t[170] & t[171] & ~t[174]) | (~t[168] & t[169] & t[172] & t[173] & ~t[174]) | (t[168] & ~t[170] & ~t[172] & t[174]) | (~t[168] & t[170] & t[172] & t[174]);
  assign t[139] = (t[168] & t[169] & ~t[170] & ~t[172] & t[173] & ~t[174]) | (t[168] & t[170] & ~t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & t[172] & ~t[173] & ~t[174]) | (~t[168] & ~t[170] & ~t[171] & t[172] & ~t[173]) | (~t[168] & ~t[169] & ~t[171] & t[172] & ~t[174]) | (~t[168] & ~t[170] & t[171] & t[172] & t[173]) | (t[171] & t[172] & ~t[173] & ~t[174]);
  assign t[13] = t[92] & t[22];
  assign t[140] = (t[175] & ~t[177] & ~t[178] & ~t[179] & ~t[180]) | (t[175] & ~t[176] & ~t[178] & ~t[179] & ~t[181]) | (t[175] & ~t[176] & ~t[177] & ~t[180] & ~t[181]) | (~t[175] & t[176] & t[177] & t[178] & ~t[181]) | (~t[175] & t[176] & t[179] & t[180] & ~t[181]) | (t[175] & ~t[177] & ~t[179] & t[181]) | (~t[175] & t[177] & t[179] & t[181]);
  assign t[141] = (t[175] & t[176] & ~t[177] & ~t[179] & t[180] & ~t[181]) | (t[175] & t[177] & ~t[178] & ~t[179] & ~t[180] & t[181]) | (~t[176] & ~t[177] & t[179] & ~t[180] & ~t[181]) | (~t[175] & ~t[177] & ~t[178] & t[179] & ~t[180]) | (~t[175] & ~t[176] & ~t[178] & t[179] & ~t[181]) | (~t[175] & ~t[177] & t[178] & t[179] & t[180]) | (t[178] & t[179] & ~t[180] & ~t[181]);
  assign t[142] = (t[182] & ~t[184] & ~t[185] & ~t[186] & ~t[187]) | (t[182] & ~t[183] & ~t[185] & ~t[186] & ~t[188]) | (t[182] & ~t[183] & ~t[184] & ~t[187] & ~t[188]) | (~t[182] & t[183] & t[184] & t[185] & ~t[188]) | (~t[182] & t[183] & t[186] & t[187] & ~t[188]) | (t[182] & ~t[184] & ~t[186] & t[188]) | (~t[182] & t[184] & t[186] & t[188]);
  assign t[143] = (t[182] & t[183] & ~t[184] & t[185] & ~t[186] & ~t[188]) | (t[182] & ~t[184] & ~t[185] & t[186] & ~t[187] & t[188]) | (~t[183] & t[184] & ~t[185] & ~t[186] & ~t[188]) | (~t[182] & t[184] & ~t[185] & ~t[186] & ~t[187]) | (~t[182] & ~t[183] & t[184] & ~t[187] & ~t[188]) | (~t[182] & t[184] & t[185] & ~t[186] & t[187]) | (t[184] & ~t[185] & t[187] & ~t[188]);
  assign t[144] = (t[189] & ~t[191] & ~t[192] & ~t[193] & ~t[194]) | (t[189] & ~t[190] & ~t[192] & ~t[193] & ~t[195]) | (t[189] & ~t[190] & ~t[191] & ~t[194] & ~t[195]) | (~t[189] & t[190] & t[191] & t[192] & ~t[195]) | (~t[189] & t[190] & t[193] & t[194] & ~t[195]) | (t[189] & ~t[191] & ~t[193] & t[195]) | (~t[189] & t[191] & t[193] & t[195]);
  assign t[145] = (t[189] & t[190] & ~t[191] & t[192] & ~t[193] & ~t[195]) | (t[189] & ~t[191] & ~t[192] & t[193] & ~t[194] & t[195]) | (~t[190] & t[191] & ~t[192] & ~t[193] & ~t[195]) | (~t[189] & t[191] & ~t[192] & ~t[193] & ~t[194]) | (~t[189] & ~t[190] & t[191] & ~t[194] & ~t[195]) | (~t[189] & t[191] & t[192] & ~t[193] & t[194]) | (t[191] & ~t[192] & t[194] & ~t[195]);
  assign t[146] = (t[183] & ~t[184] & ~t[185] & ~t[186] & ~t[187]) | (~t[182] & t[183] & ~t[185] & ~t[186] & ~t[188]) | (~t[182] & t[183] & ~t[184] & ~t[187] & ~t[188]) | (t[182] & ~t[183] & t[184] & t[185] & ~t[188]) | (t[182] & ~t[183] & t[186] & t[187] & ~t[188]) | (t[183] & ~t[185] & ~t[187] & t[188]) | (~t[183] & t[185] & t[187] & t[188]);
  assign t[147] = (t[182] & t[183] & t[184] & ~t[185] & ~t[187] & ~t[188]) | (t[183] & ~t[184] & ~t[185] & ~t[186] & t[187] & t[188]) | (~t[183] & ~t[184] & t[185] & ~t[186] & ~t[187]) | (~t[182] & ~t[184] & t[185] & ~t[187] & ~t[188]) | (~t[182] & ~t[183] & t[185] & ~t[186] & ~t[188]) | (~t[183] & t[184] & t[185] & t[186] & ~t[187]) | (~t[184] & t[185] & t[186] & ~t[188]);
  assign t[148] = (t[182] & t[183] & ~t[184] & ~t[186] & t[187] & ~t[188]) | (t[182] & t[184] & ~t[185] & ~t[186] & ~t[187] & t[188]) | (~t[183] & ~t[184] & t[186] & ~t[187] & ~t[188]) | (~t[182] & ~t[184] & ~t[185] & t[186] & ~t[187]) | (~t[182] & ~t[183] & ~t[185] & t[186] & ~t[188]) | (~t[182] & ~t[184] & t[185] & t[186] & t[187]) | (t[185] & t[186] & ~t[187] & ~t[188]);
  assign t[149] = (t[182] & t[183] & ~t[185] & t[186] & ~t[187] & ~t[188]) | (t[183] & ~t[184] & t[185] & ~t[186] & ~t[187] & t[188]) | (~t[183] & ~t[184] & ~t[185] & ~t[186] & t[187]) | (~t[182] & ~t[185] & ~t[186] & t[187] & ~t[188]) | (~t[182] & ~t[183] & ~t[184] & t[187] & ~t[188]) | (~t[183] & t[184] & ~t[185] & t[186] & t[187]) | (t[184] & ~t[186] & t[187] & ~t[188]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (t[190] & ~t[191] & ~t[192] & ~t[193] & ~t[194]) | (~t[189] & t[190] & ~t[192] & ~t[193] & ~t[195]) | (~t[189] & t[190] & ~t[191] & ~t[194] & ~t[195]) | (t[189] & ~t[190] & t[191] & t[192] & ~t[195]) | (t[189] & ~t[190] & t[193] & t[194] & ~t[195]) | (t[190] & ~t[192] & ~t[194] & t[195]) | (~t[190] & t[192] & t[194] & t[195]);
  assign t[151] = (t[189] & t[190] & t[191] & ~t[192] & ~t[194] & ~t[195]) | (t[190] & ~t[191] & ~t[192] & ~t[193] & t[194] & t[195]) | (~t[190] & ~t[191] & t[192] & ~t[193] & ~t[194]) | (~t[189] & ~t[191] & t[192] & ~t[194] & ~t[195]) | (~t[189] & ~t[190] & t[192] & ~t[193] & ~t[195]) | (~t[190] & t[191] & t[192] & t[193] & ~t[194]) | (~t[191] & t[192] & t[193] & ~t[195]);
  assign t[152] = (t[189] & t[190] & ~t[191] & ~t[193] & t[194] & ~t[195]) | (t[189] & t[191] & ~t[192] & ~t[193] & ~t[194] & t[195]) | (~t[190] & ~t[191] & t[193] & ~t[194] & ~t[195]) | (~t[189] & ~t[191] & ~t[192] & t[193] & ~t[194]) | (~t[189] & ~t[190] & ~t[192] & t[193] & ~t[195]) | (~t[189] & ~t[191] & t[192] & t[193] & t[194]) | (t[192] & t[193] & ~t[194] & ~t[195]);
  assign t[153] = (t[189] & t[190] & ~t[192] & t[193] & ~t[194] & ~t[195]) | (t[190] & ~t[191] & t[192] & ~t[193] & ~t[194] & t[195]) | (~t[190] & ~t[191] & ~t[192] & ~t[193] & t[194]) | (~t[189] & ~t[192] & ~t[193] & t[194] & ~t[195]) | (~t[189] & ~t[190] & ~t[191] & t[194] & ~t[195]) | (~t[190] & t[191] & ~t[192] & t[193] & t[194]) | (t[191] & ~t[193] & t[194] & ~t[195]);
  assign t[154] = (t[196] & ~t[198] & ~t[199] & ~t[200] & ~t[201]) | (t[196] & ~t[197] & ~t[199] & ~t[200] & ~t[202]) | (t[196] & ~t[197] & ~t[198] & ~t[201] & ~t[202]) | (~t[196] & t[197] & t[198] & t[199] & ~t[202]) | (~t[196] & t[197] & t[200] & t[201] & ~t[202]) | (t[196] & ~t[198] & ~t[200] & t[202]) | (~t[196] & t[198] & t[200] & t[202]);
  assign t[155] = (t[196] & t[197] & ~t[198] & t[199] & ~t[200] & ~t[202]) | (t[196] & ~t[198] & ~t[199] & t[200] & ~t[201] & t[202]) | (~t[197] & t[198] & ~t[199] & ~t[200] & ~t[202]) | (~t[196] & t[198] & ~t[199] & ~t[200] & ~t[201]) | (~t[196] & ~t[197] & t[198] & ~t[201] & ~t[202]) | (~t[196] & t[198] & t[199] & ~t[200] & t[201]) | (t[198] & ~t[199] & t[201] & ~t[202]);
  assign t[156] = (t[197] & ~t[198] & ~t[199] & ~t[200] & ~t[201]) | (~t[196] & t[197] & ~t[199] & ~t[200] & ~t[202]) | (~t[196] & t[197] & ~t[198] & ~t[201] & ~t[202]) | (t[196] & ~t[197] & t[198] & t[199] & ~t[202]) | (t[196] & ~t[197] & t[200] & t[201] & ~t[202]) | (t[197] & ~t[199] & ~t[201] & t[202]) | (~t[197] & t[199] & t[201] & t[202]);
  assign t[157] = (t[196] & t[197] & t[198] & ~t[199] & ~t[201] & ~t[202]) | (t[197] & ~t[198] & ~t[199] & ~t[200] & t[201] & t[202]) | (~t[197] & ~t[198] & t[199] & ~t[200] & ~t[201]) | (~t[196] & ~t[198] & t[199] & ~t[201] & ~t[202]) | (~t[196] & ~t[197] & t[199] & ~t[200] & ~t[202]) | (~t[197] & t[198] & t[199] & t[200] & ~t[201]) | (~t[198] & t[199] & t[200] & ~t[202]);
  assign t[158] = (t[196] & t[197] & ~t[198] & ~t[200] & t[201] & ~t[202]) | (t[196] & t[198] & ~t[199] & ~t[200] & ~t[201] & t[202]) | (~t[197] & ~t[198] & t[200] & ~t[201] & ~t[202]) | (~t[196] & ~t[198] & ~t[199] & t[200] & ~t[201]) | (~t[196] & ~t[197] & ~t[199] & t[200] & ~t[202]) | (~t[196] & ~t[198] & t[199] & t[200] & t[201]) | (t[199] & t[200] & ~t[201] & ~t[202]);
  assign t[159] = (t[196] & t[197] & ~t[199] & t[200] & ~t[201] & ~t[202]) | (t[197] & ~t[198] & t[199] & ~t[200] & ~t[201] & t[202]) | (~t[197] & ~t[198] & ~t[199] & ~t[200] & t[201]) | (~t[196] & ~t[199] & ~t[200] & t[201] & ~t[202]) | (~t[196] & ~t[197] & ~t[198] & t[201] & ~t[202]) | (~t[197] & t[198] & ~t[199] & t[200] & t[201]) | (t[198] & ~t[200] & t[201] & ~t[202]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = (t[168] & t[169] & ~t[170] & t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[170] & ~t[171] & t[172] & ~t[173] & t[174]) | (~t[169] & t[170] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[169] & t[170] & ~t[173] & ~t[174]) | (~t[168] & t[170] & t[171] & ~t[172] & t[173]) | (t[170] & ~t[171] & t[173] & ~t[174]);
  assign t[161] = (t[203] & ~t[205] & ~t[206] & ~t[207] & ~t[208]) | (t[203] & ~t[204] & ~t[206] & ~t[207] & ~t[209]) | (t[203] & ~t[204] & ~t[205] & ~t[208] & ~t[209]) | (~t[203] & t[204] & t[205] & t[206] & ~t[209]) | (~t[203] & t[204] & t[207] & t[208] & ~t[209]) | (t[203] & ~t[205] & ~t[207] & t[209]) | (~t[203] & t[205] & t[207] & t[209]);
  assign t[162] = (t[203] & t[204] & ~t[205] & ~t[207] & t[208] & ~t[209]) | (t[203] & t[205] & ~t[206] & ~t[207] & ~t[208] & t[209]) | (~t[204] & ~t[205] & t[207] & ~t[208] & ~t[209]) | (~t[203] & ~t[205] & ~t[206] & t[207] & ~t[208]) | (~t[203] & ~t[204] & ~t[206] & t[207] & ~t[209]) | (~t[203] & ~t[205] & t[206] & t[207] & t[208]) | (t[206] & t[207] & ~t[208] & ~t[209]);
  assign t[163] = (t[169] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & t[169] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[169] & ~t[170] & ~t[173] & ~t[174]) | (t[168] & ~t[169] & t[170] & t[171] & ~t[174]) | (t[168] & ~t[169] & t[172] & t[173] & ~t[174]) | (t[169] & ~t[171] & ~t[173] & t[174]) | (~t[169] & t[171] & t[173] & t[174]);
  assign t[164] = (t[168] & t[169] & t[170] & ~t[171] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & ~t[171] & ~t[172] & t[173] & t[174]) | (~t[169] & ~t[170] & t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[170] & t[171] & ~t[173] & ~t[174]) | (~t[168] & ~t[169] & t[171] & ~t[172] & ~t[174]) | (~t[169] & t[170] & t[171] & t[172] & ~t[173]) | (~t[170] & t[171] & t[172] & ~t[174]);
  assign t[165] = (t[168] & t[169] & ~t[171] & t[172] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & ~t[171] & ~t[172] & t[173]) | (~t[168] & ~t[171] & ~t[172] & t[173] & ~t[174]) | (~t[168] & ~t[169] & ~t[170] & t[173] & ~t[174]) | (~t[169] & t[170] & ~t[171] & t[172] & t[173]) | (t[170] & ~t[172] & t[173] & ~t[174]);
  assign t[166] = (t[210] & ~t[212] & ~t[213] & ~t[214] & ~t[215]) | (t[210] & ~t[211] & ~t[213] & ~t[214] & ~t[216]) | (t[210] & ~t[211] & ~t[212] & ~t[215] & ~t[216]) | (~t[210] & t[211] & t[212] & t[213] & ~t[216]) | (~t[210] & t[211] & t[214] & t[215] & ~t[216]) | (t[210] & ~t[212] & ~t[214] & t[216]) | (~t[210] & t[212] & t[214] & t[216]);
  assign t[167] = (t[210] & t[211] & ~t[212] & ~t[214] & t[215] & ~t[216]) | (t[210] & t[212] & ~t[213] & ~t[214] & ~t[215] & t[216]) | (~t[211] & ~t[212] & t[214] & ~t[215] & ~t[216]) | (~t[210] & ~t[212] & ~t[213] & t[214] & ~t[215]) | (~t[210] & ~t[211] & ~t[213] & t[214] & ~t[216]) | (~t[210] & ~t[212] & t[213] & t[214] & t[215]) | (t[213] & t[214] & ~t[215] & ~t[216]);
  assign t[168] = t[217] ^ x[7];
  assign t[169] = t[218] ^ x[61];
  assign t[16] = t[26] ^ t[14];
  assign t[170] = t[219] ^ x[51];
  assign t[171] = t[220] ^ x[62];
  assign t[172] = t[221] ^ x[8];
  assign t[173] = t[222] ^ x[63];
  assign t[174] = t[223] ^ x[6];
  assign t[175] = t[224] ^ x[15];
  assign t[176] = t[225] ^ x[10];
  assign t[177] = t[226] ^ x[11];
  assign t[178] = t[227] ^ x[12];
  assign t[179] = t[228] ^ x[16];
  assign t[17] = t[93] & t[27];
  assign t[180] = t[229] ^ x[13];
  assign t[181] = t[230] ^ x[14];
  assign t[182] = t[231] ^ x[22];
  assign t[183] = t[232] ^ x[31];
  assign t[184] = t[233] ^ x[23];
  assign t[185] = t[234] ^ x[32];
  assign t[186] = t[235] ^ x[33];
  assign t[187] = t[236] ^ x[34];
  assign t[188] = t[237] ^ x[21];
  assign t[189] = t[238] ^ x[29];
  assign t[18] = t[28] & t[29];
  assign t[190] = t[239] ^ x[35];
  assign t[191] = t[240] ^ x[30];
  assign t[192] = t[241] ^ x[36];
  assign t[193] = t[242] ^ x[37];
  assign t[194] = t[243] ^ x[38];
  assign t[195] = t[244] ^ x[28];
  assign t[196] = t[245] ^ x[44];
  assign t[197] = t[246] ^ x[46];
  assign t[198] = t[247] ^ x[45];
  assign t[199] = t[248] ^ x[47];
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = t[249] ^ x[48];
  assign t[201] = t[250] ^ x[49];
  assign t[202] = t[251] ^ x[43];
  assign t[203] = t[252] ^ x[58];
  assign t[204] = t[253] ^ x[53];
  assign t[205] = t[254] ^ x[54];
  assign t[206] = t[255] ^ x[55];
  assign t[207] = t[256] ^ x[59];
  assign t[208] = t[257] ^ x[56];
  assign t[209] = t[258] ^ x[57];
  assign t[20] = t[31] ^ t[18];
  assign t[210] = t[259] ^ x[70];
  assign t[211] = t[260] ^ x[65];
  assign t[212] = t[261] ^ x[66];
  assign t[213] = t[262] ^ x[67];
  assign t[214] = t[263] ^ x[71];
  assign t[215] = t[264] ^ x[68];
  assign t[216] = t[265] ^ x[69];
  assign t[217] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[218] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[219] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[21] = t[32] ^ t[33];
  assign t[220] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[221] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[222] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[223] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[224] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[225] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[226] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[227] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[228] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[229] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[22] = t[34] ^ t[35];
  assign t[230] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[231] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[232] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[233] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[234] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[235] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[236] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[237] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[238] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[239] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[23] = ~(t[94]);
  assign t[240] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[241] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[242] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[243] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[244] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[245] = (x[39] & ~x[40] & ~x[41]) | (~x[39] & x[40] & ~x[41]) | (~x[39] & ~x[40] & x[41]) | (x[39] & x[40] & x[41]);
  assign t[246] = (x[39] & ~x[40] & ~x[42]) | (~x[39] & x[40] & ~x[42]) | (~x[39] & ~x[40] & x[42]) | (x[39] & x[40] & x[42]);
  assign t[247] = (x[39] & ~x[41]) | (~x[39] & x[41]);
  assign t[248] = (x[39] & ~x[42]) | (~x[39] & x[42]);
  assign t[249] = (x[40] & ~x[41]) | (~x[40] & x[41]);
  assign t[24] = ~(t[92] ^ t[23]);
  assign t[250] = (x[40] & ~x[42]) | (~x[40] & x[42]);
  assign t[251] = (x[41] & ~x[42]) | (~x[41] & x[42]);
  assign t[252] = (x[52] & ~1'b0 & ~1'b0) | (~x[52] & 1'b0 & ~1'b0) | (~x[52] & ~1'b0 & 1'b0) | (x[52] & 1'b0 & 1'b0);
  assign t[253] = (x[52] & ~1'b0 & ~1'b0) | (~x[52] & 1'b0 & ~1'b0) | (~x[52] & ~1'b0 & 1'b0) | (x[52] & 1'b0 & 1'b0);
  assign t[254] = (x[52] & ~1'b0) | (~x[52] & 1'b0);
  assign t[255] = (x[52] & ~1'b0) | (~x[52] & 1'b0);
  assign t[256] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[257] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[258] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[259] = (x[64] & ~1'b0 & ~1'b0) | (~x[64] & 1'b0 & ~1'b0) | (~x[64] & ~1'b0 & 1'b0) | (x[64] & 1'b0 & 1'b0);
  assign t[25] = t[95] ^ t[94];
  assign t[260] = (x[64] & ~1'b0 & ~1'b0) | (~x[64] & 1'b0 & ~1'b0) | (~x[64] & ~1'b0 & 1'b0) | (x[64] & 1'b0 & 1'b0);
  assign t[261] = (x[64] & ~1'b0) | (~x[64] & 1'b0);
  assign t[262] = (x[64] & ~1'b0) | (~x[64] & 1'b0);
  assign t[263] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[264] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[265] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[96]);
  assign t[29] = ~(t[93] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[90]);
  assign t[30] = t[97] ^ t[96];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[92] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[92] ^ t[44];
  assign t[37] = t[93] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[93] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[98] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[94] ^ t[99];
  assign t[45] = t[96] ^ t[100];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[101]);
  assign t[48] = ~(t[98] ^ t[47]);
  assign t[49] = t[102] ^ t[101];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[98] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[98] ^ t[54];
  assign t[54] = t[101] ^ t[103];
  assign t[55] = x[0] ? x[50] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[104]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63] ^ t[64]);
  assign t[61] = ~(t[65] ^ t[66]);
  assign t[62] = ~(t[67] ^ t[105]);
  assign t[63] = t[68] ^ t[14];
  assign t[64] = t[8] ^ t[69];
  assign t[65] = t[70] ^ t[18];
  assign t[66] = t[10] ^ t[71];
  assign t[67] = ~t[72];
  assign t[68] = t[25] ^ t[35];
  assign t[69] = t[92] ^ t[23];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[30] ^ t[38];
  assign t[71] = t[93] ^ t[28];
  assign t[72] = ~(t[73] ^ t[74]);
  assign t[73] = t[75] ^ t[41];
  assign t[74] = t[32] ^ t[76];
  assign t[75] = t[49] ^ t[52];
  assign t[76] = t[98] ^ t[47];
  assign t[77] = x[0] ? x[60] : t[78];
  assign t[78] = ~(t[79] ^ t[80]);
  assign t[79] = ~(t[81] ^ t[106]);
  assign t[7] = ~(t[12] ^ t[91]);
  assign t[80] = ~(t[82] ^ t[83]);
  assign t[81] = ~t[84];
  assign t[82] = ~(t[85]);
  assign t[83] = ~(t[86]);
  assign t[84] = ~(t[87] ^ t[107]);
  assign t[85] = t[44] ^ t[14];
  assign t[86] = t[45] ^ t[18];
  assign t[87] = ~t[88];
  assign t[88] = ~(t[89]);
  assign t[89] = t[54] ^ t[41];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[108] & ~t[109]) | (~t[108] & t[109]);
  assign t[91] = (t[110] & ~t[111]) | (~t[110] & t[111]);
  assign t[92] = (t[112] & ~t[113]) | (~t[112] & t[113]);
  assign t[93] = (t[114] & ~t[115]) | (~t[114] & t[115]);
  assign t[94] = (t[112] & ~t[117] & ~t[119]) | (~t[116] & t[117] & ~t[118]) | (~t[112] & ~t[117] & t[119]) | (t[116] & t[117] & t[118]);
  assign t[95] = (t[112] & ~t[118]) | (~t[112] & t[118]);
  assign t[96] = (t[114] & ~t[121] & ~t[123]) | (~t[120] & t[121] & ~t[122]) | (~t[114] & ~t[121] & t[123]) | (t[120] & t[121] & t[122]);
  assign t[97] = (t[114] & ~t[122]) | (~t[114] & t[122]);
  assign t[98] = (t[124] & ~t[125]) | (~t[124] & t[125]);
  assign t[99] = (t[112] & ~t[117] & ~t[118]) | (~t[116] & t[117] & ~t[119]) | (~t[112] & ~t[117] & t[118]) | (t[116] & t[117] & t[119]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[55] & ~t[77]) | (~t[0] & t[55] & ~t[77]) | (~t[0] & ~t[55] & t[77]) | (t[0] & t[55] & t[77]);
endmodule

module R2ind162(x, y);
 input [71:0] x;
 output y;

 wire [262:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[121] & ~t[124] & ~t[125]) | (~t[123] & t[124] & ~t[126]) | (~t[121] & ~t[124] & t[125]) | (t[123] & t[124] & t[126]);
  assign t[101] = (t[105] & ~t[127]) | (~t[105] & t[127]);
  assign t[102] = (t[128] & ~t[129]) | (~t[128] & t[129]);
  assign t[103] = (t[105] & ~t[131] & ~t[106]) | (~t[130] & t[131] & ~t[132]) | (~t[105] & ~t[131] & t[106]) | (t[130] & t[131] & t[132]);
  assign t[104] = (t[133] & ~t[134]) | (~t[133] & t[134]);
  assign t[105] = t[135] ^ x[7];
  assign t[106] = t[136] ^ x[8];
  assign t[107] = t[137] ^ x[15];
  assign t[108] = t[138] ^ x[16];
  assign t[109] = t[139] ^ x[22];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[140] ^ x[23];
  assign t[111] = t[141] ^ x[29];
  assign t[112] = t[142] ^ x[30];
  assign t[113] = t[143] ^ x[31];
  assign t[114] = t[144] ^ x[32];
  assign t[115] = t[145] ^ x[33];
  assign t[116] = t[146] ^ x[34];
  assign t[117] = t[147] ^ x[35];
  assign t[118] = t[148] ^ x[36];
  assign t[119] = t[149] ^ x[37];
  assign t[11] = t[19] & t[20];
  assign t[120] = t[150] ^ x[38];
  assign t[121] = t[151] ^ x[44];
  assign t[122] = t[152] ^ x[45];
  assign t[123] = t[153] ^ x[46];
  assign t[124] = t[154] ^ x[47];
  assign t[125] = t[155] ^ x[48];
  assign t[126] = t[156] ^ x[49];
  assign t[127] = t[157] ^ x[51];
  assign t[128] = t[158] ^ x[58];
  assign t[129] = t[159] ^ x[59];
  assign t[12] = ~t[21];
  assign t[130] = t[160] ^ x[61];
  assign t[131] = t[161] ^ x[62];
  assign t[132] = t[162] ^ x[63];
  assign t[133] = t[163] ^ x[70];
  assign t[134] = t[164] ^ x[71];
  assign t[135] = (t[165] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (t[165] & ~t[166] & ~t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[166] & ~t[167] & ~t[170] & ~t[171]) | (~t[165] & t[166] & t[167] & t[168] & ~t[171]) | (~t[165] & t[166] & t[169] & t[170] & ~t[171]) | (t[165] & ~t[167] & ~t[169] & t[171]) | (~t[165] & t[167] & t[169] & t[171]);
  assign t[136] = (t[165] & t[166] & ~t[167] & ~t[169] & t[170] & ~t[171]) | (t[165] & t[167] & ~t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & t[169] & ~t[170] & ~t[171]) | (~t[165] & ~t[167] & ~t[168] & t[169] & ~t[170]) | (~t[165] & ~t[166] & ~t[168] & t[169] & ~t[171]) | (~t[165] & ~t[167] & t[168] & t[169] & t[170]) | (t[168] & t[169] & ~t[170] & ~t[171]);
  assign t[137] = (t[172] & ~t[174] & ~t[175] & ~t[176] & ~t[177]) | (t[172] & ~t[173] & ~t[175] & ~t[176] & ~t[178]) | (t[172] & ~t[173] & ~t[174] & ~t[177] & ~t[178]) | (~t[172] & t[173] & t[174] & t[175] & ~t[178]) | (~t[172] & t[173] & t[176] & t[177] & ~t[178]) | (t[172] & ~t[174] & ~t[176] & t[178]) | (~t[172] & t[174] & t[176] & t[178]);
  assign t[138] = (t[172] & t[173] & ~t[174] & ~t[176] & t[177] & ~t[178]) | (t[172] & t[174] & ~t[175] & ~t[176] & ~t[177] & t[178]) | (~t[173] & ~t[174] & t[176] & ~t[177] & ~t[178]) | (~t[172] & ~t[174] & ~t[175] & t[176] & ~t[177]) | (~t[172] & ~t[173] & ~t[175] & t[176] & ~t[178]) | (~t[172] & ~t[174] & t[175] & t[176] & t[177]) | (t[175] & t[176] & ~t[177] & ~t[178]);
  assign t[139] = (t[179] & ~t[181] & ~t[182] & ~t[183] & ~t[184]) | (t[179] & ~t[180] & ~t[182] & ~t[183] & ~t[185]) | (t[179] & ~t[180] & ~t[181] & ~t[184] & ~t[185]) | (~t[179] & t[180] & t[181] & t[182] & ~t[185]) | (~t[179] & t[180] & t[183] & t[184] & ~t[185]) | (t[179] & ~t[181] & ~t[183] & t[185]) | (~t[179] & t[181] & t[183] & t[185]);
  assign t[13] = t[89] & t[22];
  assign t[140] = (t[179] & t[180] & ~t[181] & t[182] & ~t[183] & ~t[185]) | (t[179] & ~t[181] & ~t[182] & t[183] & ~t[184] & t[185]) | (~t[180] & t[181] & ~t[182] & ~t[183] & ~t[185]) | (~t[179] & t[181] & ~t[182] & ~t[183] & ~t[184]) | (~t[179] & ~t[180] & t[181] & ~t[184] & ~t[185]) | (~t[179] & t[181] & t[182] & ~t[183] & t[184]) | (t[181] & ~t[182] & t[184] & ~t[185]);
  assign t[141] = (t[186] & ~t[188] & ~t[189] & ~t[190] & ~t[191]) | (t[186] & ~t[187] & ~t[189] & ~t[190] & ~t[192]) | (t[186] & ~t[187] & ~t[188] & ~t[191] & ~t[192]) | (~t[186] & t[187] & t[188] & t[189] & ~t[192]) | (~t[186] & t[187] & t[190] & t[191] & ~t[192]) | (t[186] & ~t[188] & ~t[190] & t[192]) | (~t[186] & t[188] & t[190] & t[192]);
  assign t[142] = (t[186] & t[187] & ~t[188] & t[189] & ~t[190] & ~t[192]) | (t[186] & ~t[188] & ~t[189] & t[190] & ~t[191] & t[192]) | (~t[187] & t[188] & ~t[189] & ~t[190] & ~t[192]) | (~t[186] & t[188] & ~t[189] & ~t[190] & ~t[191]) | (~t[186] & ~t[187] & t[188] & ~t[191] & ~t[192]) | (~t[186] & t[188] & t[189] & ~t[190] & t[191]) | (t[188] & ~t[189] & t[191] & ~t[192]);
  assign t[143] = (t[180] & ~t[181] & ~t[182] & ~t[183] & ~t[184]) | (~t[179] & t[180] & ~t[182] & ~t[183] & ~t[185]) | (~t[179] & t[180] & ~t[181] & ~t[184] & ~t[185]) | (t[179] & ~t[180] & t[181] & t[182] & ~t[185]) | (t[179] & ~t[180] & t[183] & t[184] & ~t[185]) | (t[180] & ~t[182] & ~t[184] & t[185]) | (~t[180] & t[182] & t[184] & t[185]);
  assign t[144] = (t[179] & t[180] & t[181] & ~t[182] & ~t[184] & ~t[185]) | (t[180] & ~t[181] & ~t[182] & ~t[183] & t[184] & t[185]) | (~t[180] & ~t[181] & t[182] & ~t[183] & ~t[184]) | (~t[179] & ~t[181] & t[182] & ~t[184] & ~t[185]) | (~t[179] & ~t[180] & t[182] & ~t[183] & ~t[185]) | (~t[180] & t[181] & t[182] & t[183] & ~t[184]) | (~t[181] & t[182] & t[183] & ~t[185]);
  assign t[145] = (t[179] & t[180] & ~t[181] & ~t[183] & t[184] & ~t[185]) | (t[179] & t[181] & ~t[182] & ~t[183] & ~t[184] & t[185]) | (~t[180] & ~t[181] & t[183] & ~t[184] & ~t[185]) | (~t[179] & ~t[181] & ~t[182] & t[183] & ~t[184]) | (~t[179] & ~t[180] & ~t[182] & t[183] & ~t[185]) | (~t[179] & ~t[181] & t[182] & t[183] & t[184]) | (t[182] & t[183] & ~t[184] & ~t[185]);
  assign t[146] = (t[179] & t[180] & ~t[182] & t[183] & ~t[184] & ~t[185]) | (t[180] & ~t[181] & t[182] & ~t[183] & ~t[184] & t[185]) | (~t[180] & ~t[181] & ~t[182] & ~t[183] & t[184]) | (~t[179] & ~t[182] & ~t[183] & t[184] & ~t[185]) | (~t[179] & ~t[180] & ~t[181] & t[184] & ~t[185]) | (~t[180] & t[181] & ~t[182] & t[183] & t[184]) | (t[181] & ~t[183] & t[184] & ~t[185]);
  assign t[147] = (t[187] & ~t[188] & ~t[189] & ~t[190] & ~t[191]) | (~t[186] & t[187] & ~t[189] & ~t[190] & ~t[192]) | (~t[186] & t[187] & ~t[188] & ~t[191] & ~t[192]) | (t[186] & ~t[187] & t[188] & t[189] & ~t[192]) | (t[186] & ~t[187] & t[190] & t[191] & ~t[192]) | (t[187] & ~t[189] & ~t[191] & t[192]) | (~t[187] & t[189] & t[191] & t[192]);
  assign t[148] = (t[186] & t[187] & t[188] & ~t[189] & ~t[191] & ~t[192]) | (t[187] & ~t[188] & ~t[189] & ~t[190] & t[191] & t[192]) | (~t[187] & ~t[188] & t[189] & ~t[190] & ~t[191]) | (~t[186] & ~t[188] & t[189] & ~t[191] & ~t[192]) | (~t[186] & ~t[187] & t[189] & ~t[190] & ~t[192]) | (~t[187] & t[188] & t[189] & t[190] & ~t[191]) | (~t[188] & t[189] & t[190] & ~t[192]);
  assign t[149] = (t[186] & t[187] & ~t[188] & ~t[190] & t[191] & ~t[192]) | (t[186] & t[188] & ~t[189] & ~t[190] & ~t[191] & t[192]) | (~t[187] & ~t[188] & t[190] & ~t[191] & ~t[192]) | (~t[186] & ~t[188] & ~t[189] & t[190] & ~t[191]) | (~t[186] & ~t[187] & ~t[189] & t[190] & ~t[192]) | (~t[186] & ~t[188] & t[189] & t[190] & t[191]) | (t[189] & t[190] & ~t[191] & ~t[192]);
  assign t[14] = t[23] & t[24];
  assign t[150] = (t[186] & t[187] & ~t[189] & t[190] & ~t[191] & ~t[192]) | (t[187] & ~t[188] & t[189] & ~t[190] & ~t[191] & t[192]) | (~t[187] & ~t[188] & ~t[189] & ~t[190] & t[191]) | (~t[186] & ~t[189] & ~t[190] & t[191] & ~t[192]) | (~t[186] & ~t[187] & ~t[188] & t[191] & ~t[192]) | (~t[187] & t[188] & ~t[189] & t[190] & t[191]) | (t[188] & ~t[190] & t[191] & ~t[192]);
  assign t[151] = (t[193] & ~t[195] & ~t[196] & ~t[197] & ~t[198]) | (t[193] & ~t[194] & ~t[196] & ~t[197] & ~t[199]) | (t[193] & ~t[194] & ~t[195] & ~t[198] & ~t[199]) | (~t[193] & t[194] & t[195] & t[196] & ~t[199]) | (~t[193] & t[194] & t[197] & t[198] & ~t[199]) | (t[193] & ~t[195] & ~t[197] & t[199]) | (~t[193] & t[195] & t[197] & t[199]);
  assign t[152] = (t[193] & t[194] & ~t[195] & t[196] & ~t[197] & ~t[199]) | (t[193] & ~t[195] & ~t[196] & t[197] & ~t[198] & t[199]) | (~t[194] & t[195] & ~t[196] & ~t[197] & ~t[199]) | (~t[193] & t[195] & ~t[196] & ~t[197] & ~t[198]) | (~t[193] & ~t[194] & t[195] & ~t[198] & ~t[199]) | (~t[193] & t[195] & t[196] & ~t[197] & t[198]) | (t[195] & ~t[196] & t[198] & ~t[199]);
  assign t[153] = (t[194] & ~t[195] & ~t[196] & ~t[197] & ~t[198]) | (~t[193] & t[194] & ~t[196] & ~t[197] & ~t[199]) | (~t[193] & t[194] & ~t[195] & ~t[198] & ~t[199]) | (t[193] & ~t[194] & t[195] & t[196] & ~t[199]) | (t[193] & ~t[194] & t[197] & t[198] & ~t[199]) | (t[194] & ~t[196] & ~t[198] & t[199]) | (~t[194] & t[196] & t[198] & t[199]);
  assign t[154] = (t[193] & t[194] & t[195] & ~t[196] & ~t[198] & ~t[199]) | (t[194] & ~t[195] & ~t[196] & ~t[197] & t[198] & t[199]) | (~t[194] & ~t[195] & t[196] & ~t[197] & ~t[198]) | (~t[193] & ~t[195] & t[196] & ~t[198] & ~t[199]) | (~t[193] & ~t[194] & t[196] & ~t[197] & ~t[199]) | (~t[194] & t[195] & t[196] & t[197] & ~t[198]) | (~t[195] & t[196] & t[197] & ~t[199]);
  assign t[155] = (t[193] & t[194] & ~t[195] & ~t[197] & t[198] & ~t[199]) | (t[193] & t[195] & ~t[196] & ~t[197] & ~t[198] & t[199]) | (~t[194] & ~t[195] & t[197] & ~t[198] & ~t[199]) | (~t[193] & ~t[195] & ~t[196] & t[197] & ~t[198]) | (~t[193] & ~t[194] & ~t[196] & t[197] & ~t[199]) | (~t[193] & ~t[195] & t[196] & t[197] & t[198]) | (t[196] & t[197] & ~t[198] & ~t[199]);
  assign t[156] = (t[193] & t[194] & ~t[196] & t[197] & ~t[198] & ~t[199]) | (t[194] & ~t[195] & t[196] & ~t[197] & ~t[198] & t[199]) | (~t[194] & ~t[195] & ~t[196] & ~t[197] & t[198]) | (~t[193] & ~t[196] & ~t[197] & t[198] & ~t[199]) | (~t[193] & ~t[194] & ~t[195] & t[198] & ~t[199]) | (~t[194] & t[195] & ~t[196] & t[197] & t[198]) | (t[195] & ~t[197] & t[198] & ~t[199]);
  assign t[157] = (t[165] & t[166] & ~t[167] & t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[167] & ~t[168] & t[169] & ~t[170] & t[171]) | (~t[166] & t[167] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[166] & t[167] & ~t[170] & ~t[171]) | (~t[165] & t[167] & t[168] & ~t[169] & t[170]) | (t[167] & ~t[168] & t[170] & ~t[171]);
  assign t[158] = (t[200] & ~t[202] & ~t[203] & ~t[204] & ~t[205]) | (t[200] & ~t[201] & ~t[203] & ~t[204] & ~t[206]) | (t[200] & ~t[201] & ~t[202] & ~t[205] & ~t[206]) | (~t[200] & t[201] & t[202] & t[203] & ~t[206]) | (~t[200] & t[201] & t[204] & t[205] & ~t[206]) | (t[200] & ~t[202] & ~t[204] & t[206]) | (~t[200] & t[202] & t[204] & t[206]);
  assign t[159] = (t[200] & t[201] & ~t[202] & ~t[204] & t[205] & ~t[206]) | (t[200] & t[202] & ~t[203] & ~t[204] & ~t[205] & t[206]) | (~t[201] & ~t[202] & t[204] & ~t[205] & ~t[206]) | (~t[200] & ~t[202] & ~t[203] & t[204] & ~t[205]) | (~t[200] & ~t[201] & ~t[203] & t[204] & ~t[206]) | (~t[200] & ~t[202] & t[203] & t[204] & t[205]) | (t[203] & t[204] & ~t[205] & ~t[206]);
  assign t[15] = t[25] ^ t[23];
  assign t[160] = (t[166] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & t[166] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[166] & ~t[167] & ~t[170] & ~t[171]) | (t[165] & ~t[166] & t[167] & t[168] & ~t[171]) | (t[165] & ~t[166] & t[169] & t[170] & ~t[171]) | (t[166] & ~t[168] & ~t[170] & t[171]) | (~t[166] & t[168] & t[170] & t[171]);
  assign t[161] = (t[165] & t[166] & t[167] & ~t[168] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & ~t[168] & ~t[169] & t[170] & t[171]) | (~t[166] & ~t[167] & t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[167] & t[168] & ~t[170] & ~t[171]) | (~t[165] & ~t[166] & t[168] & ~t[169] & ~t[171]) | (~t[166] & t[167] & t[168] & t[169] & ~t[170]) | (~t[167] & t[168] & t[169] & ~t[171]);
  assign t[162] = (t[165] & t[166] & ~t[168] & t[169] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & ~t[168] & ~t[169] & t[170]) | (~t[165] & ~t[168] & ~t[169] & t[170] & ~t[171]) | (~t[165] & ~t[166] & ~t[167] & t[170] & ~t[171]) | (~t[166] & t[167] & ~t[168] & t[169] & t[170]) | (t[167] & ~t[169] & t[170] & ~t[171]);
  assign t[163] = (t[207] & ~t[209] & ~t[210] & ~t[211] & ~t[212]) | (t[207] & ~t[208] & ~t[210] & ~t[211] & ~t[213]) | (t[207] & ~t[208] & ~t[209] & ~t[212] & ~t[213]) | (~t[207] & t[208] & t[209] & t[210] & ~t[213]) | (~t[207] & t[208] & t[211] & t[212] & ~t[213]) | (t[207] & ~t[209] & ~t[211] & t[213]) | (~t[207] & t[209] & t[211] & t[213]);
  assign t[164] = (t[207] & t[208] & ~t[209] & ~t[211] & t[212] & ~t[213]) | (t[207] & t[209] & ~t[210] & ~t[211] & ~t[212] & t[213]) | (~t[208] & ~t[209] & t[211] & ~t[212] & ~t[213]) | (~t[207] & ~t[209] & ~t[210] & t[211] & ~t[212]) | (~t[207] & ~t[208] & ~t[210] & t[211] & ~t[213]) | (~t[207] & ~t[209] & t[210] & t[211] & t[212]) | (t[210] & t[211] & ~t[212] & ~t[213]);
  assign t[165] = t[214] ^ x[7];
  assign t[166] = t[215] ^ x[61];
  assign t[167] = t[216] ^ x[51];
  assign t[168] = t[217] ^ x[62];
  assign t[169] = t[218] ^ x[8];
  assign t[16] = t[26] ^ t[14];
  assign t[170] = t[219] ^ x[63];
  assign t[171] = t[220] ^ x[6];
  assign t[172] = t[221] ^ x[15];
  assign t[173] = t[222] ^ x[10];
  assign t[174] = t[223] ^ x[11];
  assign t[175] = t[224] ^ x[12];
  assign t[176] = t[225] ^ x[16];
  assign t[177] = t[226] ^ x[13];
  assign t[178] = t[227] ^ x[14];
  assign t[179] = t[228] ^ x[22];
  assign t[17] = t[90] & t[27];
  assign t[180] = t[229] ^ x[31];
  assign t[181] = t[230] ^ x[23];
  assign t[182] = t[231] ^ x[32];
  assign t[183] = t[232] ^ x[33];
  assign t[184] = t[233] ^ x[34];
  assign t[185] = t[234] ^ x[21];
  assign t[186] = t[235] ^ x[29];
  assign t[187] = t[236] ^ x[35];
  assign t[188] = t[237] ^ x[30];
  assign t[189] = t[238] ^ x[36];
  assign t[18] = t[28] & t[29];
  assign t[190] = t[239] ^ x[37];
  assign t[191] = t[240] ^ x[38];
  assign t[192] = t[241] ^ x[28];
  assign t[193] = t[242] ^ x[44];
  assign t[194] = t[243] ^ x[46];
  assign t[195] = t[244] ^ x[45];
  assign t[196] = t[245] ^ x[47];
  assign t[197] = t[246] ^ x[48];
  assign t[198] = t[247] ^ x[49];
  assign t[199] = t[248] ^ x[43];
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = t[249] ^ x[58];
  assign t[201] = t[250] ^ x[53];
  assign t[202] = t[251] ^ x[54];
  assign t[203] = t[252] ^ x[55];
  assign t[204] = t[253] ^ x[59];
  assign t[205] = t[254] ^ x[56];
  assign t[206] = t[255] ^ x[57];
  assign t[207] = t[256] ^ x[70];
  assign t[208] = t[257] ^ x[65];
  assign t[209] = t[258] ^ x[66];
  assign t[20] = t[31] ^ t[18];
  assign t[210] = t[259] ^ x[67];
  assign t[211] = t[260] ^ x[71];
  assign t[212] = t[261] ^ x[68];
  assign t[213] = t[262] ^ x[69];
  assign t[214] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[215] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[216] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[217] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[218] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[219] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[21] = t[32] ^ t[33];
  assign t[220] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[221] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[222] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[223] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[224] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[225] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[226] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[227] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[228] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[229] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[22] = t[34] ^ t[35];
  assign t[230] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[231] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[232] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[233] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[234] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[235] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[236] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[237] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[238] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[239] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[23] = ~(t[91]);
  assign t[240] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[241] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[242] = (x[39] & ~x[40] & ~x[41]) | (~x[39] & x[40] & ~x[41]) | (~x[39] & ~x[40] & x[41]) | (x[39] & x[40] & x[41]);
  assign t[243] = (x[39] & ~x[40] & ~x[42]) | (~x[39] & x[40] & ~x[42]) | (~x[39] & ~x[40] & x[42]) | (x[39] & x[40] & x[42]);
  assign t[244] = (x[39] & ~x[41]) | (~x[39] & x[41]);
  assign t[245] = (x[39] & ~x[42]) | (~x[39] & x[42]);
  assign t[246] = (x[40] & ~x[41]) | (~x[40] & x[41]);
  assign t[247] = (x[40] & ~x[42]) | (~x[40] & x[42]);
  assign t[248] = (x[41] & ~x[42]) | (~x[41] & x[42]);
  assign t[249] = (x[52] & ~1'b0 & ~1'b0) | (~x[52] & 1'b0 & ~1'b0) | (~x[52] & ~1'b0 & 1'b0) | (x[52] & 1'b0 & 1'b0);
  assign t[24] = ~(t[89] ^ t[23]);
  assign t[250] = (x[52] & ~1'b0 & ~1'b0) | (~x[52] & 1'b0 & ~1'b0) | (~x[52] & ~1'b0 & 1'b0) | (x[52] & 1'b0 & 1'b0);
  assign t[251] = (x[52] & ~1'b0) | (~x[52] & 1'b0);
  assign t[252] = (x[52] & ~1'b0) | (~x[52] & 1'b0);
  assign t[253] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[254] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[255] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[256] = (x[64] & ~1'b0 & ~1'b0) | (~x[64] & 1'b0 & ~1'b0) | (~x[64] & ~1'b0 & 1'b0) | (x[64] & 1'b0 & 1'b0);
  assign t[257] = (x[64] & ~1'b0 & ~1'b0) | (~x[64] & 1'b0 & ~1'b0) | (~x[64] & ~1'b0 & 1'b0) | (x[64] & 1'b0 & 1'b0);
  assign t[258] = (x[64] & ~1'b0) | (~x[64] & 1'b0);
  assign t[259] = (x[64] & ~1'b0) | (~x[64] & 1'b0);
  assign t[25] = t[92] ^ t[91];
  assign t[260] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[261] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[262] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[93]);
  assign t[29] = ~(t[90] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[87]);
  assign t[30] = t[94] ^ t[93];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[89] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[89] ^ t[44];
  assign t[37] = t[90] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[90] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[95] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[91] ^ t[96];
  assign t[45] = t[93] ^ t[97];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[98]);
  assign t[48] = ~(t[95] ^ t[47]);
  assign t[49] = t[99] ^ t[98];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[95] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[95] ^ t[54];
  assign t[54] = t[98] ^ t[100];
  assign t[55] = x[0] ? x[50] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[101]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63] ^ t[64]);
  assign t[61] = ~(t[65] ^ t[66]);
  assign t[62] = ~(t[67] ^ t[102]);
  assign t[63] = t[68] ^ t[14];
  assign t[64] = t[8] ^ t[69];
  assign t[65] = t[70] ^ t[18];
  assign t[66] = t[10] ^ t[71];
  assign t[67] = ~t[72];
  assign t[68] = t[25] ^ t[35];
  assign t[69] = t[89] ^ t[23];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[30] ^ t[38];
  assign t[71] = t[90] ^ t[28];
  assign t[72] = ~(t[73] ^ t[74]);
  assign t[73] = t[75] ^ t[41];
  assign t[74] = t[32] ^ t[76];
  assign t[75] = t[49] ^ t[52];
  assign t[76] = t[95] ^ t[47];
  assign t[77] = x[0] ? x[60] : t[78];
  assign t[78] = ~(t[79] ^ t[80]);
  assign t[79] = ~(t[81] ^ t[103]);
  assign t[7] = ~(t[12] ^ t[88]);
  assign t[80] = ~(t[82] ^ t[83]);
  assign t[81] = ~t[84];
  assign t[82] = ~(t[63]);
  assign t[83] = ~(t[65]);
  assign t[84] = ~(t[85] ^ t[104]);
  assign t[85] = ~t[86];
  assign t[86] = ~(t[73]);
  assign t[87] = (t[105] & ~t[106]) | (~t[105] & t[106]);
  assign t[88] = (t[107] & ~t[108]) | (~t[107] & t[108]);
  assign t[89] = (t[109] & ~t[110]) | (~t[109] & t[110]);
  assign t[8] = t[13] ^ t[14];
  assign t[90] = (t[111] & ~t[112]) | (~t[111] & t[112]);
  assign t[91] = (t[109] & ~t[114] & ~t[116]) | (~t[113] & t[114] & ~t[115]) | (~t[109] & ~t[114] & t[116]) | (t[113] & t[114] & t[115]);
  assign t[92] = (t[109] & ~t[115]) | (~t[109] & t[115]);
  assign t[93] = (t[111] & ~t[118] & ~t[120]) | (~t[117] & t[118] & ~t[119]) | (~t[111] & ~t[118] & t[120]) | (t[117] & t[118] & t[119]);
  assign t[94] = (t[111] & ~t[119]) | (~t[111] & t[119]);
  assign t[95] = (t[121] & ~t[122]) | (~t[121] & t[122]);
  assign t[96] = (t[109] & ~t[114] & ~t[115]) | (~t[113] & t[114] & ~t[116]) | (~t[109] & ~t[114] & t[115]) | (t[113] & t[114] & t[116]);
  assign t[97] = (t[111] & ~t[118] & ~t[119]) | (~t[117] & t[118] & ~t[120]) | (~t[111] & ~t[118] & t[119]) | (t[117] & t[118] & t[120]);
  assign t[98] = (t[121] & ~t[124] & ~t[126]) | (~t[123] & t[124] & ~t[125]) | (~t[121] & ~t[124] & t[126]) | (t[123] & t[124] & t[125]);
  assign t[99] = (t[121] & ~t[125]) | (~t[121] & t[125]);
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[55] & ~t[77]) | (~t[0] & t[55] & ~t[77]) | (~t[0] & ~t[55] & t[77]) | (t[0] & t[55] & t[77]);
endmodule

module R2ind163(x, y);
 input [62:0] x;
 output y;

 wire [221:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[127] ^ x[45];
  assign t[101] = t[128] ^ x[46];
  assign t[102] = t[129] ^ x[47];
  assign t[103] = t[130] ^ x[48];
  assign t[104] = t[131] ^ x[49];
  assign t[105] = t[132] ^ x[50];
  assign t[106] = t[133] ^ x[52];
  assign t[107] = t[134] ^ x[53];
  assign t[108] = t[135] ^ x[54];
  assign t[109] = t[136] ^ x[61];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[137] ^ x[62];
  assign t[111] = (t[138] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[141] & ~t[142] & ~t[144]) | (t[138] & ~t[139] & ~t[140] & ~t[143] & ~t[144]) | (~t[138] & t[139] & t[140] & t[141] & ~t[144]) | (~t[138] & t[139] & t[142] & t[143] & ~t[144]) | (t[138] & ~t[140] & ~t[142] & t[144]) | (~t[138] & t[140] & t[142] & t[144]);
  assign t[112] = (t[138] & t[139] & ~t[140] & ~t[142] & t[143] & ~t[144]) | (t[138] & t[140] & ~t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & t[142] & ~t[143] & ~t[144]) | (~t[138] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[138] & ~t[139] & ~t[141] & t[142] & ~t[144]) | (~t[138] & ~t[140] & t[141] & t[142] & t[143]) | (t[141] & t[142] & ~t[143] & ~t[144]);
  assign t[113] = (t[145] & ~t[147] & ~t[148] & ~t[149] & ~t[150]) | (t[145] & ~t[146] & ~t[148] & ~t[149] & ~t[151]) | (t[145] & ~t[146] & ~t[147] & ~t[150] & ~t[151]) | (~t[145] & t[146] & t[147] & t[148] & ~t[151]) | (~t[145] & t[146] & t[149] & t[150] & ~t[151]) | (t[145] & ~t[147] & ~t[149] & t[151]) | (~t[145] & t[147] & t[149] & t[151]);
  assign t[114] = (t[145] & t[146] & ~t[147] & ~t[149] & t[150] & ~t[151]) | (t[145] & t[147] & ~t[148] & ~t[149] & ~t[150] & t[151]) | (~t[146] & ~t[147] & t[149] & ~t[150] & ~t[151]) | (~t[145] & ~t[147] & ~t[148] & t[149] & ~t[150]) | (~t[145] & ~t[146] & ~t[148] & t[149] & ~t[151]) | (~t[145] & ~t[147] & t[148] & t[149] & t[150]) | (t[148] & t[149] & ~t[150] & ~t[151]);
  assign t[115] = (t[152] & ~t[154] & ~t[155] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & ~t[155] & ~t[156] & ~t[158]) | (t[152] & ~t[153] & ~t[154] & ~t[157] & ~t[158]) | (~t[152] & t[153] & t[154] & t[155] & ~t[158]) | (~t[152] & t[153] & t[156] & t[157] & ~t[158]) | (t[152] & ~t[154] & ~t[156] & t[158]) | (~t[152] & t[154] & t[156] & t[158]);
  assign t[116] = (t[152] & t[153] & ~t[154] & t[155] & ~t[156] & ~t[158]) | (t[152] & ~t[154] & ~t[155] & t[156] & ~t[157] & t[158]) | (~t[153] & t[154] & ~t[155] & ~t[156] & ~t[158]) | (~t[152] & t[154] & ~t[155] & ~t[156] & ~t[157]) | (~t[152] & ~t[153] & t[154] & ~t[157] & ~t[158]) | (~t[152] & t[154] & t[155] & ~t[156] & t[157]) | (t[154] & ~t[155] & t[157] & ~t[158]);
  assign t[117] = (t[159] & ~t[161] & ~t[162] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & ~t[162] & ~t[163] & ~t[165]) | (t[159] & ~t[160] & ~t[161] & ~t[164] & ~t[165]) | (~t[159] & t[160] & t[161] & t[162] & ~t[165]) | (~t[159] & t[160] & t[163] & t[164] & ~t[165]) | (t[159] & ~t[161] & ~t[163] & t[165]) | (~t[159] & t[161] & t[163] & t[165]);
  assign t[118] = (t[159] & t[160] & ~t[161] & t[162] & ~t[163] & ~t[165]) | (t[159] & ~t[161] & ~t[162] & t[163] & ~t[164] & t[165]) | (~t[160] & t[161] & ~t[162] & ~t[163] & ~t[165]) | (~t[159] & t[161] & ~t[162] & ~t[163] & ~t[164]) | (~t[159] & ~t[160] & t[161] & ~t[164] & ~t[165]) | (~t[159] & t[161] & t[162] & ~t[163] & t[164]) | (t[161] & ~t[162] & t[164] & ~t[165]);
  assign t[119] = (t[153] & ~t[154] & ~t[155] & ~t[156] & ~t[157]) | (~t[152] & t[153] & ~t[155] & ~t[156] & ~t[158]) | (~t[152] & t[153] & ~t[154] & ~t[157] & ~t[158]) | (t[152] & ~t[153] & t[154] & t[155] & ~t[158]) | (t[152] & ~t[153] & t[156] & t[157] & ~t[158]) | (t[153] & ~t[155] & ~t[157] & t[158]) | (~t[153] & t[155] & t[157] & t[158]);
  assign t[11] = t[19] & t[20];
  assign t[120] = (t[152] & t[153] & t[154] & ~t[155] & ~t[157] & ~t[158]) | (t[153] & ~t[154] & ~t[155] & ~t[156] & t[157] & t[158]) | (~t[153] & ~t[154] & t[155] & ~t[156] & ~t[157]) | (~t[152] & ~t[154] & t[155] & ~t[157] & ~t[158]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[158]) | (~t[153] & t[154] & t[155] & t[156] & ~t[157]) | (~t[154] & t[155] & t[156] & ~t[158]);
  assign t[121] = (t[152] & t[153] & ~t[154] & ~t[156] & t[157] & ~t[158]) | (t[152] & t[154] & ~t[155] & ~t[156] & ~t[157] & t[158]) | (~t[153] & ~t[154] & t[156] & ~t[157] & ~t[158]) | (~t[152] & ~t[154] & ~t[155] & t[156] & ~t[157]) | (~t[152] & ~t[153] & ~t[155] & t[156] & ~t[158]) | (~t[152] & ~t[154] & t[155] & t[156] & t[157]) | (t[155] & t[156] & ~t[157] & ~t[158]);
  assign t[122] = (t[152] & t[153] & ~t[155] & t[156] & ~t[157] & ~t[158]) | (t[153] & ~t[154] & t[155] & ~t[156] & ~t[157] & t[158]) | (~t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[155] & ~t[156] & t[157] & ~t[158]) | (~t[152] & ~t[153] & ~t[154] & t[157] & ~t[158]) | (~t[153] & t[154] & ~t[155] & t[156] & t[157]) | (t[154] & ~t[156] & t[157] & ~t[158]);
  assign t[123] = (t[160] & ~t[161] & ~t[162] & ~t[163] & ~t[164]) | (~t[159] & t[160] & ~t[162] & ~t[163] & ~t[165]) | (~t[159] & t[160] & ~t[161] & ~t[164] & ~t[165]) | (t[159] & ~t[160] & t[161] & t[162] & ~t[165]) | (t[159] & ~t[160] & t[163] & t[164] & ~t[165]) | (t[160] & ~t[162] & ~t[164] & t[165]) | (~t[160] & t[162] & t[164] & t[165]);
  assign t[124] = (t[159] & t[160] & t[161] & ~t[162] & ~t[164] & ~t[165]) | (t[160] & ~t[161] & ~t[162] & ~t[163] & t[164] & t[165]) | (~t[160] & ~t[161] & t[162] & ~t[163] & ~t[164]) | (~t[159] & ~t[161] & t[162] & ~t[164] & ~t[165]) | (~t[159] & ~t[160] & t[162] & ~t[163] & ~t[165]) | (~t[160] & t[161] & t[162] & t[163] & ~t[164]) | (~t[161] & t[162] & t[163] & ~t[165]);
  assign t[125] = (t[159] & t[160] & ~t[161] & ~t[163] & t[164] & ~t[165]) | (t[159] & t[161] & ~t[162] & ~t[163] & ~t[164] & t[165]) | (~t[160] & ~t[161] & t[163] & ~t[164] & ~t[165]) | (~t[159] & ~t[161] & ~t[162] & t[163] & ~t[164]) | (~t[159] & ~t[160] & ~t[162] & t[163] & ~t[165]) | (~t[159] & ~t[161] & t[162] & t[163] & t[164]) | (t[162] & t[163] & ~t[164] & ~t[165]);
  assign t[126] = (t[159] & t[160] & ~t[162] & t[163] & ~t[164] & ~t[165]) | (t[160] & ~t[161] & t[162] & ~t[163] & ~t[164] & t[165]) | (~t[160] & ~t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[162] & ~t[163] & t[164] & ~t[165]) | (~t[159] & ~t[160] & ~t[161] & t[164] & ~t[165]) | (~t[160] & t[161] & ~t[162] & t[163] & t[164]) | (t[161] & ~t[163] & t[164] & ~t[165]);
  assign t[127] = (t[166] & ~t[168] & ~t[169] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & ~t[169] & ~t[170] & ~t[172]) | (t[166] & ~t[167] & ~t[168] & ~t[171] & ~t[172]) | (~t[166] & t[167] & t[168] & t[169] & ~t[172]) | (~t[166] & t[167] & t[170] & t[171] & ~t[172]) | (t[166] & ~t[168] & ~t[170] & t[172]) | (~t[166] & t[168] & t[170] & t[172]);
  assign t[128] = (t[166] & t[167] & ~t[168] & t[169] & ~t[170] & ~t[172]) | (t[166] & ~t[168] & ~t[169] & t[170] & ~t[171] & t[172]) | (~t[167] & t[168] & ~t[169] & ~t[170] & ~t[172]) | (~t[166] & t[168] & ~t[169] & ~t[170] & ~t[171]) | (~t[166] & ~t[167] & t[168] & ~t[171] & ~t[172]) | (~t[166] & t[168] & t[169] & ~t[170] & t[171]) | (t[168] & ~t[169] & t[171] & ~t[172]);
  assign t[129] = (t[167] & ~t[168] & ~t[169] & ~t[170] & ~t[171]) | (~t[166] & t[167] & ~t[169] & ~t[170] & ~t[172]) | (~t[166] & t[167] & ~t[168] & ~t[171] & ~t[172]) | (t[166] & ~t[167] & t[168] & t[169] & ~t[172]) | (t[166] & ~t[167] & t[170] & t[171] & ~t[172]) | (t[167] & ~t[169] & ~t[171] & t[172]) | (~t[167] & t[169] & t[171] & t[172]);
  assign t[12] = ~t[21];
  assign t[130] = (t[166] & t[167] & t[168] & ~t[169] & ~t[171] & ~t[172]) | (t[167] & ~t[168] & ~t[169] & ~t[170] & t[171] & t[172]) | (~t[167] & ~t[168] & t[169] & ~t[170] & ~t[171]) | (~t[166] & ~t[168] & t[169] & ~t[171] & ~t[172]) | (~t[166] & ~t[167] & t[169] & ~t[170] & ~t[172]) | (~t[167] & t[168] & t[169] & t[170] & ~t[171]) | (~t[168] & t[169] & t[170] & ~t[172]);
  assign t[131] = (t[166] & t[167] & ~t[168] & ~t[170] & t[171] & ~t[172]) | (t[166] & t[168] & ~t[169] & ~t[170] & ~t[171] & t[172]) | (~t[167] & ~t[168] & t[170] & ~t[171] & ~t[172]) | (~t[166] & ~t[168] & ~t[169] & t[170] & ~t[171]) | (~t[166] & ~t[167] & ~t[169] & t[170] & ~t[172]) | (~t[166] & ~t[168] & t[169] & t[170] & t[171]) | (t[169] & t[170] & ~t[171] & ~t[172]);
  assign t[132] = (t[166] & t[167] & ~t[169] & t[170] & ~t[171] & ~t[172]) | (t[167] & ~t[168] & t[169] & ~t[170] & ~t[171] & t[172]) | (~t[167] & ~t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[169] & ~t[170] & t[171] & ~t[172]) | (~t[166] & ~t[167] & ~t[168] & t[171] & ~t[172]) | (~t[167] & t[168] & ~t[169] & t[170] & t[171]) | (t[168] & ~t[170] & t[171] & ~t[172]);
  assign t[133] = (t[139] & ~t[140] & ~t[141] & ~t[142] & ~t[143]) | (~t[138] & t[139] & ~t[141] & ~t[142] & ~t[144]) | (~t[138] & t[139] & ~t[140] & ~t[143] & ~t[144]) | (t[138] & ~t[139] & t[140] & t[141] & ~t[144]) | (t[138] & ~t[139] & t[142] & t[143] & ~t[144]) | (t[139] & ~t[141] & ~t[143] & t[144]) | (~t[139] & t[141] & t[143] & t[144]);
  assign t[134] = (t[138] & t[139] & t[140] & ~t[141] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & ~t[141] & ~t[142] & t[143] & t[144]) | (~t[139] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (~t[138] & ~t[140] & t[141] & ~t[143] & ~t[144]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[144]) | (~t[139] & t[140] & t[141] & t[142] & ~t[143]) | (~t[140] & t[141] & t[142] & ~t[144]);
  assign t[135] = (t[138] & t[139] & ~t[141] & t[142] & ~t[143] & ~t[144]) | (t[139] & ~t[140] & t[141] & ~t[142] & ~t[143] & t[144]) | (~t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[141] & ~t[142] & t[143] & ~t[144]) | (~t[138] & ~t[139] & ~t[140] & t[143] & ~t[144]) | (~t[139] & t[140] & ~t[141] & t[142] & t[143]) | (t[140] & ~t[142] & t[143] & ~t[144]);
  assign t[136] = (t[173] & ~t[175] & ~t[176] & ~t[177] & ~t[178]) | (t[173] & ~t[174] & ~t[176] & ~t[177] & ~t[179]) | (t[173] & ~t[174] & ~t[175] & ~t[178] & ~t[179]) | (~t[173] & t[174] & t[175] & t[176] & ~t[179]) | (~t[173] & t[174] & t[177] & t[178] & ~t[179]) | (t[173] & ~t[175] & ~t[177] & t[179]) | (~t[173] & t[175] & t[177] & t[179]);
  assign t[137] = (t[173] & t[174] & ~t[175] & ~t[177] & t[178] & ~t[179]) | (t[173] & t[175] & ~t[176] & ~t[177] & ~t[178] & t[179]) | (~t[174] & ~t[175] & t[177] & ~t[178] & ~t[179]) | (~t[173] & ~t[175] & ~t[176] & t[177] & ~t[178]) | (~t[173] & ~t[174] & ~t[176] & t[177] & ~t[179]) | (~t[173] & ~t[175] & t[176] & t[177] & t[178]) | (t[176] & t[177] & ~t[178] & ~t[179]);
  assign t[138] = t[180] ^ x[8];
  assign t[139] = t[181] ^ x[52];
  assign t[13] = t[70] & t[22];
  assign t[140] = t[182] ^ x[6];
  assign t[141] = t[183] ^ x[53];
  assign t[142] = t[184] ^ x[9];
  assign t[143] = t[185] ^ x[54];
  assign t[144] = t[186] ^ x[7];
  assign t[145] = t[187] ^ x[16];
  assign t[146] = t[188] ^ x[11];
  assign t[147] = t[189] ^ x[12];
  assign t[148] = t[190] ^ x[13];
  assign t[149] = t[191] ^ x[17];
  assign t[14] = t[23] & t[24];
  assign t[150] = t[192] ^ x[14];
  assign t[151] = t[193] ^ x[15];
  assign t[152] = t[194] ^ x[23];
  assign t[153] = t[195] ^ x[32];
  assign t[154] = t[196] ^ x[24];
  assign t[155] = t[197] ^ x[33];
  assign t[156] = t[198] ^ x[34];
  assign t[157] = t[199] ^ x[35];
  assign t[158] = t[200] ^ x[22];
  assign t[159] = t[201] ^ x[30];
  assign t[15] = t[25] ^ t[23];
  assign t[160] = t[202] ^ x[36];
  assign t[161] = t[203] ^ x[31];
  assign t[162] = t[204] ^ x[37];
  assign t[163] = t[205] ^ x[38];
  assign t[164] = t[206] ^ x[39];
  assign t[165] = t[207] ^ x[29];
  assign t[166] = t[208] ^ x[45];
  assign t[167] = t[209] ^ x[47];
  assign t[168] = t[210] ^ x[46];
  assign t[169] = t[211] ^ x[48];
  assign t[16] = t[26] ^ t[14];
  assign t[170] = t[212] ^ x[49];
  assign t[171] = t[213] ^ x[50];
  assign t[172] = t[214] ^ x[44];
  assign t[173] = t[215] ^ x[61];
  assign t[174] = t[216] ^ x[56];
  assign t[175] = t[217] ^ x[57];
  assign t[176] = t[218] ^ x[58];
  assign t[177] = t[219] ^ x[62];
  assign t[178] = t[220] ^ x[59];
  assign t[179] = t[221] ^ x[60];
  assign t[17] = t[71] & t[27];
  assign t[180] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[181] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[182] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[183] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[184] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[185] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[186] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[187] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[188] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[189] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[192] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[193] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[194] = (x[18] & ~x[19] & ~x[20]) | (~x[18] & x[19] & ~x[20]) | (~x[18] & ~x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[195] = (x[18] & ~x[19] & ~x[21]) | (~x[18] & x[19] & ~x[21]) | (~x[18] & ~x[19] & x[21]) | (x[18] & x[19] & x[21]);
  assign t[196] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[197] = (x[18] & ~x[21]) | (~x[18] & x[21]);
  assign t[198] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[199] = (x[19] & ~x[21]) | (~x[19] & x[21]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[20] & ~x[21]) | (~x[20] & x[21]);
  assign t[201] = (x[25] & ~x[26] & ~x[27]) | (~x[25] & x[26] & ~x[27]) | (~x[25] & ~x[26] & x[27]) | (x[25] & x[26] & x[27]);
  assign t[202] = (x[25] & ~x[26] & ~x[28]) | (~x[25] & x[26] & ~x[28]) | (~x[25] & ~x[26] & x[28]) | (x[25] & x[26] & x[28]);
  assign t[203] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[204] = (x[25] & ~x[28]) | (~x[25] & x[28]);
  assign t[205] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[206] = (x[26] & ~x[28]) | (~x[26] & x[28]);
  assign t[207] = (x[27] & ~x[28]) | (~x[27] & x[28]);
  assign t[208] = (x[40] & ~x[41] & ~x[42]) | (~x[40] & x[41] & ~x[42]) | (~x[40] & ~x[41] & x[42]) | (x[40] & x[41] & x[42]);
  assign t[209] = (x[40] & ~x[41] & ~x[43]) | (~x[40] & x[41] & ~x[43]) | (~x[40] & ~x[41] & x[43]) | (x[40] & x[41] & x[43]);
  assign t[20] = t[31] ^ t[18];
  assign t[210] = (x[40] & ~x[42]) | (~x[40] & x[42]);
  assign t[211] = (x[40] & ~x[43]) | (~x[40] & x[43]);
  assign t[212] = (x[41] & ~x[42]) | (~x[41] & x[42]);
  assign t[213] = (x[41] & ~x[43]) | (~x[41] & x[43]);
  assign t[214] = (x[42] & ~x[43]) | (~x[42] & x[43]);
  assign t[215] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[216] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[217] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[218] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[219] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[21] = t[32] ^ t[33];
  assign t[220] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[221] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[72]);
  assign t[24] = ~(t[70] ^ t[23]);
  assign t[25] = t[73] ^ t[72];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[74]);
  assign t[29] = ~(t[71] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[68]);
  assign t[30] = t[75] ^ t[74];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[70] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[70] ^ t[44];
  assign t[37] = t[71] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[71] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[76] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[72] ^ t[77];
  assign t[45] = t[74] ^ t[78];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[79]);
  assign t[48] = ~(t[76] ^ t[47]);
  assign t[49] = t[80] ^ t[79];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[76] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[76] ^ t[54];
  assign t[54] = t[79] ^ t[81];
  assign t[55] = x[0] ? x[51] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[82]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = ~(t[64]);
  assign t[62] = ~(t[65] ^ t[83]);
  assign t[63] = t[44] ^ t[14];
  assign t[64] = t[45] ^ t[18];
  assign t[65] = ~t[66];
  assign t[66] = ~(t[67]);
  assign t[67] = t[54] ^ t[41];
  assign t[68] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[69] = (t[86] & ~t[87]) | (~t[86] & t[87]);
  assign t[6] = t[10] ^ t[11];
  assign t[70] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[71] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[72] = (t[88] & ~t[93] & ~t[95]) | (~t[92] & t[93] & ~t[94]) | (~t[88] & ~t[93] & t[95]) | (t[92] & t[93] & t[94]);
  assign t[73] = (t[88] & ~t[94]) | (~t[88] & t[94]);
  assign t[74] = (t[90] & ~t[97] & ~t[99]) | (~t[96] & t[97] & ~t[98]) | (~t[90] & ~t[97] & t[99]) | (t[96] & t[97] & t[98]);
  assign t[75] = (t[90] & ~t[98]) | (~t[90] & t[98]);
  assign t[76] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[77] = (t[88] & ~t[93] & ~t[94]) | (~t[92] & t[93] & ~t[95]) | (~t[88] & ~t[93] & t[94]) | (t[92] & t[93] & t[95]);
  assign t[78] = (t[90] & ~t[97] & ~t[98]) | (~t[96] & t[97] & ~t[99]) | (~t[90] & ~t[97] & t[98]) | (t[96] & t[97] & t[99]);
  assign t[79] = (t[100] & ~t[103] & ~t[105]) | (~t[102] & t[103] & ~t[104]) | (~t[100] & ~t[103] & t[105]) | (t[102] & t[103] & t[104]);
  assign t[7] = ~(t[12] ^ t[69]);
  assign t[80] = (t[100] & ~t[104]) | (~t[100] & t[104]);
  assign t[81] = (t[100] & ~t[103] & ~t[104]) | (~t[102] & t[103] & ~t[105]) | (~t[100] & ~t[103] & t[104]) | (t[102] & t[103] & t[105]);
  assign t[82] = (t[84] & ~t[107] & ~t[108]) | (~t[106] & t[107] & ~t[85]) | (~t[84] & ~t[107] & t[108]) | (t[106] & t[107] & t[85]);
  assign t[83] = (t[109] & ~t[110]) | (~t[109] & t[110]);
  assign t[84] = t[111] ^ x[8];
  assign t[85] = t[112] ^ x[9];
  assign t[86] = t[113] ^ x[16];
  assign t[87] = t[114] ^ x[17];
  assign t[88] = t[115] ^ x[23];
  assign t[89] = t[116] ^ x[24];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[117] ^ x[30];
  assign t[91] = t[118] ^ x[31];
  assign t[92] = t[119] ^ x[32];
  assign t[93] = t[120] ^ x[33];
  assign t[94] = t[121] ^ x[34];
  assign t[95] = t[122] ^ x[35];
  assign t[96] = t[123] ^ x[36];
  assign t[97] = t[124] ^ x[37];
  assign t[98] = t[125] ^ x[38];
  assign t[99] = t[126] ^ x[39];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[55]) | (~t[0] & t[55]);
endmodule

module R2ind164(x, y);
 input [62:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[127] ^ x[37];
  assign t[101] = t[128] ^ x[38];
  assign t[102] = t[129] ^ x[39];
  assign t[103] = t[130] ^ x[45];
  assign t[104] = t[131] ^ x[46];
  assign t[105] = t[132] ^ x[47];
  assign t[106] = t[133] ^ x[48];
  assign t[107] = t[134] ^ x[49];
  assign t[108] = t[135] ^ x[50];
  assign t[109] = t[136] ^ x[52];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[137] ^ x[53];
  assign t[111] = t[138] ^ x[54];
  assign t[112] = t[139] ^ x[61];
  assign t[113] = t[140] ^ x[62];
  assign t[114] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[115] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[116] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[117] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[118] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[119] = (t[155] & t[156] & ~t[157] & t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[157] & ~t[158] & t[159] & ~t[160] & t[161]) | (~t[156] & t[157] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[156] & t[157] & ~t[160] & ~t[161]) | (~t[155] & t[157] & t[158] & ~t[159] & t[160]) | (t[157] & ~t[158] & t[160] & ~t[161]);
  assign t[11] = t[19] & t[20];
  assign t[120] = (t[162] & ~t[164] & ~t[165] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & ~t[165] & ~t[166] & ~t[168]) | (t[162] & ~t[163] & ~t[164] & ~t[167] & ~t[168]) | (~t[162] & t[163] & t[164] & t[165] & ~t[168]) | (~t[162] & t[163] & t[166] & t[167] & ~t[168]) | (t[162] & ~t[164] & ~t[166] & t[168]) | (~t[162] & t[164] & t[166] & t[168]);
  assign t[121] = (t[162] & t[163] & ~t[164] & t[165] & ~t[166] & ~t[168]) | (t[162] & ~t[164] & ~t[165] & t[166] & ~t[167] & t[168]) | (~t[163] & t[164] & ~t[165] & ~t[166] & ~t[168]) | (~t[162] & t[164] & ~t[165] & ~t[166] & ~t[167]) | (~t[162] & ~t[163] & t[164] & ~t[167] & ~t[168]) | (~t[162] & t[164] & t[165] & ~t[166] & t[167]) | (t[164] & ~t[165] & t[167] & ~t[168]);
  assign t[122] = (t[156] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (~t[155] & t[156] & ~t[158] & ~t[159] & ~t[161]) | (~t[155] & t[156] & ~t[157] & ~t[160] & ~t[161]) | (t[155] & ~t[156] & t[157] & t[158] & ~t[161]) | (t[155] & ~t[156] & t[159] & t[160] & ~t[161]) | (t[156] & ~t[158] & ~t[160] & t[161]) | (~t[156] & t[158] & t[160] & t[161]);
  assign t[123] = (t[155] & t[156] & t[157] & ~t[158] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & ~t[158] & ~t[159] & t[160] & t[161]) | (~t[156] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (~t[155] & ~t[157] & t[158] & ~t[160] & ~t[161]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[161]) | (~t[156] & t[157] & t[158] & t[159] & ~t[160]) | (~t[157] & t[158] & t[159] & ~t[161]);
  assign t[124] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[125] = (t[155] & t[156] & ~t[158] & t[159] & ~t[160] & ~t[161]) | (t[156] & ~t[157] & t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[158] & ~t[159] & t[160] & ~t[161]) | (~t[155] & ~t[156] & ~t[157] & t[160] & ~t[161]) | (~t[156] & t[157] & ~t[158] & t[159] & t[160]) | (t[157] & ~t[159] & t[160] & ~t[161]);
  assign t[126] = (t[163] & ~t[164] & ~t[165] & ~t[166] & ~t[167]) | (~t[162] & t[163] & ~t[165] & ~t[166] & ~t[168]) | (~t[162] & t[163] & ~t[164] & ~t[167] & ~t[168]) | (t[162] & ~t[163] & t[164] & t[165] & ~t[168]) | (t[162] & ~t[163] & t[166] & t[167] & ~t[168]) | (t[163] & ~t[165] & ~t[167] & t[168]) | (~t[163] & t[165] & t[167] & t[168]);
  assign t[127] = (t[162] & t[163] & t[164] & ~t[165] & ~t[167] & ~t[168]) | (t[163] & ~t[164] & ~t[165] & ~t[166] & t[167] & t[168]) | (~t[163] & ~t[164] & t[165] & ~t[166] & ~t[167]) | (~t[162] & ~t[164] & t[165] & ~t[167] & ~t[168]) | (~t[162] & ~t[163] & t[165] & ~t[166] & ~t[168]) | (~t[163] & t[164] & t[165] & t[166] & ~t[167]) | (~t[164] & t[165] & t[166] & ~t[168]);
  assign t[128] = (t[162] & t[163] & ~t[164] & ~t[166] & t[167] & ~t[168]) | (t[162] & t[164] & ~t[165] & ~t[166] & ~t[167] & t[168]) | (~t[163] & ~t[164] & t[166] & ~t[167] & ~t[168]) | (~t[162] & ~t[164] & ~t[165] & t[166] & ~t[167]) | (~t[162] & ~t[163] & ~t[165] & t[166] & ~t[168]) | (~t[162] & ~t[164] & t[165] & t[166] & t[167]) | (t[165] & t[166] & ~t[167] & ~t[168]);
  assign t[129] = (t[162] & t[163] & ~t[165] & t[166] & ~t[167] & ~t[168]) | (t[163] & ~t[164] & t[165] & ~t[166] & ~t[167] & t[168]) | (~t[163] & ~t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[165] & ~t[166] & t[167] & ~t[168]) | (~t[162] & ~t[163] & ~t[164] & t[167] & ~t[168]) | (~t[163] & t[164] & ~t[165] & t[166] & t[167]) | (t[164] & ~t[166] & t[167] & ~t[168]);
  assign t[12] = ~t[21];
  assign t[130] = (t[169] & ~t[171] & ~t[172] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & ~t[172] & ~t[173] & ~t[175]) | (t[169] & ~t[170] & ~t[171] & ~t[174] & ~t[175]) | (~t[169] & t[170] & t[171] & t[172] & ~t[175]) | (~t[169] & t[170] & t[173] & t[174] & ~t[175]) | (t[169] & ~t[171] & ~t[173] & t[175]) | (~t[169] & t[171] & t[173] & t[175]);
  assign t[131] = (t[169] & t[170] & ~t[171] & t[172] & ~t[173] & ~t[175]) | (t[169] & ~t[171] & ~t[172] & t[173] & ~t[174] & t[175]) | (~t[170] & t[171] & ~t[172] & ~t[173] & ~t[175]) | (~t[169] & t[171] & ~t[172] & ~t[173] & ~t[174]) | (~t[169] & ~t[170] & t[171] & ~t[174] & ~t[175]) | (~t[169] & t[171] & t[172] & ~t[173] & t[174]) | (t[171] & ~t[172] & t[174] & ~t[175]);
  assign t[132] = (t[170] & ~t[171] & ~t[172] & ~t[173] & ~t[174]) | (~t[169] & t[170] & ~t[172] & ~t[173] & ~t[175]) | (~t[169] & t[170] & ~t[171] & ~t[174] & ~t[175]) | (t[169] & ~t[170] & t[171] & t[172] & ~t[175]) | (t[169] & ~t[170] & t[173] & t[174] & ~t[175]) | (t[170] & ~t[172] & ~t[174] & t[175]) | (~t[170] & t[172] & t[174] & t[175]);
  assign t[133] = (t[169] & t[170] & t[171] & ~t[172] & ~t[174] & ~t[175]) | (t[170] & ~t[171] & ~t[172] & ~t[173] & t[174] & t[175]) | (~t[170] & ~t[171] & t[172] & ~t[173] & ~t[174]) | (~t[169] & ~t[171] & t[172] & ~t[174] & ~t[175]) | (~t[169] & ~t[170] & t[172] & ~t[173] & ~t[175]) | (~t[170] & t[171] & t[172] & t[173] & ~t[174]) | (~t[171] & t[172] & t[173] & ~t[175]);
  assign t[134] = (t[169] & t[170] & ~t[171] & ~t[173] & t[174] & ~t[175]) | (t[169] & t[171] & ~t[172] & ~t[173] & ~t[174] & t[175]) | (~t[170] & ~t[171] & t[173] & ~t[174] & ~t[175]) | (~t[169] & ~t[171] & ~t[172] & t[173] & ~t[174]) | (~t[169] & ~t[170] & ~t[172] & t[173] & ~t[175]) | (~t[169] & ~t[171] & t[172] & t[173] & t[174]) | (t[172] & t[173] & ~t[174] & ~t[175]);
  assign t[135] = (t[169] & t[170] & ~t[172] & t[173] & ~t[174] & ~t[175]) | (t[170] & ~t[171] & t[172] & ~t[173] & ~t[174] & t[175]) | (~t[170] & ~t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[172] & ~t[173] & t[174] & ~t[175]) | (~t[169] & ~t[170] & ~t[171] & t[174] & ~t[175]) | (~t[170] & t[171] & ~t[172] & t[173] & t[174]) | (t[171] & ~t[173] & t[174] & ~t[175]);
  assign t[136] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[137] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[138] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[139] = (t[176] & ~t[178] & ~t[179] & ~t[180] & ~t[181]) | (t[176] & ~t[177] & ~t[179] & ~t[180] & ~t[182]) | (t[176] & ~t[177] & ~t[178] & ~t[181] & ~t[182]) | (~t[176] & t[177] & t[178] & t[179] & ~t[182]) | (~t[176] & t[177] & t[180] & t[181] & ~t[182]) | (t[176] & ~t[178] & ~t[180] & t[182]) | (~t[176] & t[178] & t[180] & t[182]);
  assign t[13] = t[73] & t[22];
  assign t[140] = (t[176] & t[177] & ~t[178] & ~t[180] & t[181] & ~t[182]) | (t[176] & t[178] & ~t[179] & ~t[180] & ~t[181] & t[182]) | (~t[177] & ~t[178] & t[180] & ~t[181] & ~t[182]) | (~t[176] & ~t[178] & ~t[179] & t[180] & ~t[181]) | (~t[176] & ~t[177] & ~t[179] & t[180] & ~t[182]) | (~t[176] & ~t[178] & t[179] & t[180] & t[181]) | (t[179] & t[180] & ~t[181] & ~t[182]);
  assign t[141] = t[183] ^ x[8];
  assign t[142] = t[184] ^ x[52];
  assign t[143] = t[185] ^ x[6];
  assign t[144] = t[186] ^ x[53];
  assign t[145] = t[187] ^ x[9];
  assign t[146] = t[188] ^ x[54];
  assign t[147] = t[189] ^ x[7];
  assign t[148] = t[190] ^ x[16];
  assign t[149] = t[191] ^ x[11];
  assign t[14] = t[23] & t[24];
  assign t[150] = t[192] ^ x[12];
  assign t[151] = t[193] ^ x[13];
  assign t[152] = t[194] ^ x[17];
  assign t[153] = t[195] ^ x[14];
  assign t[154] = t[196] ^ x[15];
  assign t[155] = t[197] ^ x[23];
  assign t[156] = t[198] ^ x[32];
  assign t[157] = t[199] ^ x[24];
  assign t[158] = t[200] ^ x[33];
  assign t[159] = t[201] ^ x[34];
  assign t[15] = t[25] ^ t[23];
  assign t[160] = t[202] ^ x[35];
  assign t[161] = t[203] ^ x[22];
  assign t[162] = t[204] ^ x[30];
  assign t[163] = t[205] ^ x[36];
  assign t[164] = t[206] ^ x[31];
  assign t[165] = t[207] ^ x[37];
  assign t[166] = t[208] ^ x[38];
  assign t[167] = t[209] ^ x[39];
  assign t[168] = t[210] ^ x[29];
  assign t[169] = t[211] ^ x[45];
  assign t[16] = t[26] ^ t[14];
  assign t[170] = t[212] ^ x[47];
  assign t[171] = t[213] ^ x[46];
  assign t[172] = t[214] ^ x[48];
  assign t[173] = t[215] ^ x[49];
  assign t[174] = t[216] ^ x[50];
  assign t[175] = t[217] ^ x[44];
  assign t[176] = t[218] ^ x[61];
  assign t[177] = t[219] ^ x[56];
  assign t[178] = t[220] ^ x[57];
  assign t[179] = t[221] ^ x[58];
  assign t[17] = t[74] & t[27];
  assign t[180] = t[222] ^ x[62];
  assign t[181] = t[223] ^ x[59];
  assign t[182] = t[224] ^ x[60];
  assign t[183] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[184] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[185] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[186] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[187] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[188] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[189] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[18] = t[28] & t[29];
  assign t[190] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[191] = (x[10] & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0);
  assign t[192] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[193] = (x[10] & ~1'b0) | (~x[10] & 1'b0);
  assign t[194] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[195] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[196] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[197] = (x[18] & ~x[19] & ~x[20]) | (~x[18] & x[19] & ~x[20]) | (~x[18] & ~x[19] & x[20]) | (x[18] & x[19] & x[20]);
  assign t[198] = (x[18] & ~x[19] & ~x[21]) | (~x[18] & x[19] & ~x[21]) | (~x[18] & ~x[19] & x[21]) | (x[18] & x[19] & x[21]);
  assign t[199] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[19] = t[30] ^ t[28];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[18] & ~x[21]) | (~x[18] & x[21]);
  assign t[201] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[202] = (x[19] & ~x[21]) | (~x[19] & x[21]);
  assign t[203] = (x[20] & ~x[21]) | (~x[20] & x[21]);
  assign t[204] = (x[25] & ~x[26] & ~x[27]) | (~x[25] & x[26] & ~x[27]) | (~x[25] & ~x[26] & x[27]) | (x[25] & x[26] & x[27]);
  assign t[205] = (x[25] & ~x[26] & ~x[28]) | (~x[25] & x[26] & ~x[28]) | (~x[25] & ~x[26] & x[28]) | (x[25] & x[26] & x[28]);
  assign t[206] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[207] = (x[25] & ~x[28]) | (~x[25] & x[28]);
  assign t[208] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[209] = (x[26] & ~x[28]) | (~x[26] & x[28]);
  assign t[20] = t[31] ^ t[18];
  assign t[210] = (x[27] & ~x[28]) | (~x[27] & x[28]);
  assign t[211] = (x[40] & ~x[41] & ~x[42]) | (~x[40] & x[41] & ~x[42]) | (~x[40] & ~x[41] & x[42]) | (x[40] & x[41] & x[42]);
  assign t[212] = (x[40] & ~x[41] & ~x[43]) | (~x[40] & x[41] & ~x[43]) | (~x[40] & ~x[41] & x[43]) | (x[40] & x[41] & x[43]);
  assign t[213] = (x[40] & ~x[42]) | (~x[40] & x[42]);
  assign t[214] = (x[40] & ~x[43]) | (~x[40] & x[43]);
  assign t[215] = (x[41] & ~x[42]) | (~x[41] & x[42]);
  assign t[216] = (x[41] & ~x[43]) | (~x[41] & x[43]);
  assign t[217] = (x[42] & ~x[43]) | (~x[42] & x[43]);
  assign t[218] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[219] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[21] = t[32] ^ t[33];
  assign t[220] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[221] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[222] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[223] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[224] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[22] = t[34] ^ t[35];
  assign t[23] = ~(t[75]);
  assign t[24] = ~(t[73] ^ t[23]);
  assign t[25] = t[76] ^ t[75];
  assign t[26] = ~(t[36] ^ t[15]);
  assign t[27] = t[37] ^ t[38];
  assign t[28] = ~(t[77]);
  assign t[29] = ~(t[74] ^ t[28]);
  assign t[2] = ~(t[4] ^ t[71]);
  assign t[30] = t[78] ^ t[77];
  assign t[31] = ~(t[39] ^ t[19]);
  assign t[32] = t[40] ^ t[41];
  assign t[33] = t[42] & t[43];
  assign t[34] = t[73] ^ t[25];
  assign t[35] = t[23] & t[36];
  assign t[36] = t[73] ^ t[44];
  assign t[37] = t[74] ^ t[30];
  assign t[38] = t[28] & t[39];
  assign t[39] = t[74] ^ t[45];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[79] & t[46];
  assign t[41] = t[47] & t[48];
  assign t[42] = t[49] ^ t[47];
  assign t[43] = t[50] ^ t[41];
  assign t[44] = t[75] ^ t[80];
  assign t[45] = t[77] ^ t[81];
  assign t[46] = t[51] ^ t[52];
  assign t[47] = ~(t[82]);
  assign t[48] = ~(t[79] ^ t[47]);
  assign t[49] = t[83] ^ t[82];
  assign t[4] = ~t[7];
  assign t[50] = ~(t[53] ^ t[42]);
  assign t[51] = t[79] ^ t[49];
  assign t[52] = t[47] & t[53];
  assign t[53] = t[79] ^ t[54];
  assign t[54] = t[82] ^ t[84];
  assign t[55] = x[0] ? x[51] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[85]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = t[8] ^ t[9];
  assign t[60] = ~(t[63]);
  assign t[61] = ~(t[64]);
  assign t[62] = ~(t[65] ^ t[86]);
  assign t[63] = t[66] ^ t[14];
  assign t[64] = t[67] ^ t[18];
  assign t[65] = ~t[68];
  assign t[66] = t[25] ^ t[35];
  assign t[67] = t[30] ^ t[38];
  assign t[68] = ~(t[69]);
  assign t[69] = t[70] ^ t[41];
  assign t[6] = t[10] ^ t[11];
  assign t[70] = t[49] ^ t[52];
  assign t[71] = (t[87] & ~t[88]) | (~t[87] & t[88]);
  assign t[72] = (t[89] & ~t[90]) | (~t[89] & t[90]);
  assign t[73] = (t[91] & ~t[92]) | (~t[91] & t[92]);
  assign t[74] = (t[93] & ~t[94]) | (~t[93] & t[94]);
  assign t[75] = (t[91] & ~t[96] & ~t[98]) | (~t[95] & t[96] & ~t[97]) | (~t[91] & ~t[96] & t[98]) | (t[95] & t[96] & t[97]);
  assign t[76] = (t[91] & ~t[97]) | (~t[91] & t[97]);
  assign t[77] = (t[93] & ~t[100] & ~t[102]) | (~t[99] & t[100] & ~t[101]) | (~t[93] & ~t[100] & t[102]) | (t[99] & t[100] & t[101]);
  assign t[78] = (t[93] & ~t[101]) | (~t[93] & t[101]);
  assign t[79] = (t[103] & ~t[104]) | (~t[103] & t[104]);
  assign t[7] = ~(t[12] ^ t[72]);
  assign t[80] = (t[91] & ~t[96] & ~t[97]) | (~t[95] & t[96] & ~t[98]) | (~t[91] & ~t[96] & t[97]) | (t[95] & t[96] & t[98]);
  assign t[81] = (t[93] & ~t[100] & ~t[101]) | (~t[99] & t[100] & ~t[102]) | (~t[93] & ~t[100] & t[101]) | (t[99] & t[100] & t[102]);
  assign t[82] = (t[103] & ~t[106] & ~t[108]) | (~t[105] & t[106] & ~t[107]) | (~t[103] & ~t[106] & t[108]) | (t[105] & t[106] & t[107]);
  assign t[83] = (t[103] & ~t[107]) | (~t[103] & t[107]);
  assign t[84] = (t[103] & ~t[106] & ~t[107]) | (~t[105] & t[106] & ~t[108]) | (~t[103] & ~t[106] & t[107]) | (t[105] & t[106] & t[108]);
  assign t[85] = (t[87] & ~t[110] & ~t[88]) | (~t[109] & t[110] & ~t[111]) | (~t[87] & ~t[110] & t[88]) | (t[109] & t[110] & t[111]);
  assign t[86] = (t[112] & ~t[113]) | (~t[112] & t[113]);
  assign t[87] = t[114] ^ x[8];
  assign t[88] = t[115] ^ x[9];
  assign t[89] = t[116] ^ x[16];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[117] ^ x[17];
  assign t[91] = t[118] ^ x[23];
  assign t[92] = t[119] ^ x[24];
  assign t[93] = t[120] ^ x[30];
  assign t[94] = t[121] ^ x[31];
  assign t[95] = t[122] ^ x[32];
  assign t[96] = t[123] ^ x[33];
  assign t[97] = t[124] ^ x[34];
  assign t[98] = t[125] ^ x[35];
  assign t[99] = t[126] ^ x[36];
  assign t[9] = t[15] & t[16];
  assign y = (t[0] & ~t[55]) | (~t[0] & t[55]);
endmodule

module R2ind165(x, y);
 input [62:0] x;
 output y;

 wire [223:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] ^ x[44];
  assign t[101] = t[129] ^ x[45];
  assign t[102] = t[130] ^ x[46];
  assign t[103] = t[131] ^ x[47];
  assign t[104] = t[132] ^ x[48];
  assign t[105] = t[133] ^ x[49];
  assign t[106] = t[134] ^ x[51];
  assign t[107] = t[135] ^ x[52];
  assign t[108] = t[136] ^ x[53];
  assign t[109] = t[137] ^ x[54];
  assign t[10] = t[17] ^ t[18];
  assign t[110] = t[138] ^ x[61];
  assign t[111] = t[139] ^ x[62];
  assign t[112] = (t[140] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (t[140] & ~t[141] & ~t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[141] & ~t[142] & ~t[145] & ~t[146]) | (~t[140] & t[141] & t[142] & t[143] & ~t[146]) | (~t[140] & t[141] & t[144] & t[145] & ~t[146]) | (t[140] & ~t[142] & ~t[144] & t[146]) | (~t[140] & t[142] & t[144] & t[146]);
  assign t[113] = (t[140] & t[141] & ~t[142] & t[143] & ~t[144] & ~t[146]) | (t[140] & ~t[142] & ~t[143] & t[144] & ~t[145] & t[146]) | (~t[141] & t[142] & ~t[143] & ~t[144] & ~t[146]) | (~t[140] & t[142] & ~t[143] & ~t[144] & ~t[145]) | (~t[140] & ~t[141] & t[142] & ~t[145] & ~t[146]) | (~t[140] & t[142] & t[143] & ~t[144] & t[145]) | (t[142] & ~t[143] & t[145] & ~t[146]);
  assign t[114] = (t[147] & ~t[149] & ~t[150] & ~t[151] & ~t[152]) | (t[147] & ~t[148] & ~t[150] & ~t[151] & ~t[153]) | (t[147] & ~t[148] & ~t[149] & ~t[152] & ~t[153]) | (~t[147] & t[148] & t[149] & t[150] & ~t[153]) | (~t[147] & t[148] & t[151] & t[152] & ~t[153]) | (t[147] & ~t[149] & ~t[151] & t[153]) | (~t[147] & t[149] & t[151] & t[153]);
  assign t[115] = (t[147] & t[148] & ~t[149] & ~t[151] & t[152] & ~t[153]) | (t[147] & t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[153]) | (~t[147] & ~t[149] & ~t[150] & t[151] & ~t[152]) | (~t[147] & ~t[148] & ~t[150] & t[151] & ~t[153]) | (~t[147] & ~t[149] & t[150] & t[151] & t[152]) | (t[150] & t[151] & ~t[152] & ~t[153]);
  assign t[116] = (t[154] & ~t[156] & ~t[157] & ~t[158] & ~t[159]) | (t[154] & ~t[155] & ~t[157] & ~t[158] & ~t[160]) | (t[154] & ~t[155] & ~t[156] & ~t[159] & ~t[160]) | (~t[154] & t[155] & t[156] & t[157] & ~t[160]) | (~t[154] & t[155] & t[158] & t[159] & ~t[160]) | (t[154] & ~t[156] & ~t[158] & t[160]) | (~t[154] & t[156] & t[158] & t[160]);
  assign t[117] = (t[154] & t[155] & ~t[156] & t[157] & ~t[158] & ~t[160]) | (t[154] & ~t[156] & ~t[157] & t[158] & ~t[159] & t[160]) | (~t[155] & t[156] & ~t[157] & ~t[158] & ~t[160]) | (~t[154] & t[156] & ~t[157] & ~t[158] & ~t[159]) | (~t[154] & ~t[155] & t[156] & ~t[159] & ~t[160]) | (~t[154] & t[156] & t[157] & ~t[158] & t[159]) | (t[156] & ~t[157] & t[159] & ~t[160]);
  assign t[118] = (t[161] & ~t[163] & ~t[164] & ~t[165] & ~t[166]) | (t[161] & ~t[162] & ~t[164] & ~t[165] & ~t[167]) | (t[161] & ~t[162] & ~t[163] & ~t[166] & ~t[167]) | (~t[161] & t[162] & t[163] & t[164] & ~t[167]) | (~t[161] & t[162] & t[165] & t[166] & ~t[167]) | (t[161] & ~t[163] & ~t[165] & t[167]) | (~t[161] & t[163] & t[165] & t[167]);
  assign t[119] = (t[161] & t[162] & ~t[163] & t[164] & ~t[165] & ~t[167]) | (t[161] & ~t[163] & ~t[164] & t[165] & ~t[166] & t[167]) | (~t[162] & t[163] & ~t[164] & ~t[165] & ~t[167]) | (~t[161] & t[163] & ~t[164] & ~t[165] & ~t[166]) | (~t[161] & ~t[162] & t[163] & ~t[166] & ~t[167]) | (~t[161] & t[163] & t[164] & ~t[165] & t[166]) | (t[163] & ~t[164] & t[166] & ~t[167]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = (t[154] & t[155] & ~t[156] & ~t[158] & t[159] & ~t[160]) | (t[154] & t[156] & ~t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[156] & t[158] & ~t[159] & ~t[160]) | (~t[154] & ~t[156] & ~t[157] & t[158] & ~t[159]) | (~t[154] & ~t[155] & ~t[157] & t[158] & ~t[160]) | (~t[154] & ~t[156] & t[157] & t[158] & t[159]) | (t[157] & t[158] & ~t[159] & ~t[160]);
  assign t[121] = (t[155] & ~t[156] & ~t[157] & ~t[158] & ~t[159]) | (~t[154] & t[155] & ~t[157] & ~t[158] & ~t[160]) | (~t[154] & t[155] & ~t[156] & ~t[159] & ~t[160]) | (t[154] & ~t[155] & t[156] & t[157] & ~t[160]) | (t[154] & ~t[155] & t[158] & t[159] & ~t[160]) | (t[155] & ~t[157] & ~t[159] & t[160]) | (~t[155] & t[157] & t[159] & t[160]);
  assign t[122] = (t[154] & t[155] & t[156] & ~t[157] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[157] & ~t[158] & t[159] & t[160]) | (~t[155] & ~t[156] & t[157] & ~t[158] & ~t[159]) | (~t[154] & ~t[156] & t[157] & ~t[159] & ~t[160]) | (~t[154] & ~t[155] & t[157] & ~t[158] & ~t[160]) | (~t[155] & t[156] & t[157] & t[158] & ~t[159]) | (~t[156] & t[157] & t[158] & ~t[160]);
  assign t[123] = (t[154] & t[155] & ~t[157] & t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & t[157] & ~t[158] & ~t[159] & t[160]) | (~t[155] & ~t[156] & ~t[157] & ~t[158] & t[159]) | (~t[154] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[154] & ~t[155] & ~t[156] & t[159] & ~t[160]) | (~t[155] & t[156] & ~t[157] & t[158] & t[159]) | (t[156] & ~t[158] & t[159] & ~t[160]);
  assign t[124] = (t[161] & t[162] & ~t[163] & ~t[165] & t[166] & ~t[167]) | (t[161] & t[163] & ~t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[163] & t[165] & ~t[166] & ~t[167]) | (~t[161] & ~t[163] & ~t[164] & t[165] & ~t[166]) | (~t[161] & ~t[162] & ~t[164] & t[165] & ~t[167]) | (~t[161] & ~t[163] & t[164] & t[165] & t[166]) | (t[164] & t[165] & ~t[166] & ~t[167]);
  assign t[125] = (t[162] & ~t[163] & ~t[164] & ~t[165] & ~t[166]) | (~t[161] & t[162] & ~t[164] & ~t[165] & ~t[167]) | (~t[161] & t[162] & ~t[163] & ~t[166] & ~t[167]) | (t[161] & ~t[162] & t[163] & t[164] & ~t[167]) | (t[161] & ~t[162] & t[165] & t[166] & ~t[167]) | (t[162] & ~t[164] & ~t[166] & t[167]) | (~t[162] & t[164] & t[166] & t[167]);
  assign t[126] = (t[161] & t[162] & t[163] & ~t[164] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & ~t[164] & ~t[165] & t[166] & t[167]) | (~t[162] & ~t[163] & t[164] & ~t[165] & ~t[166]) | (~t[161] & ~t[163] & t[164] & ~t[166] & ~t[167]) | (~t[161] & ~t[162] & t[164] & ~t[165] & ~t[167]) | (~t[162] & t[163] & t[164] & t[165] & ~t[166]) | (~t[163] & t[164] & t[165] & ~t[167]);
  assign t[127] = (t[161] & t[162] & ~t[164] & t[165] & ~t[166] & ~t[167]) | (t[162] & ~t[163] & t[164] & ~t[165] & ~t[166] & t[167]) | (~t[162] & ~t[163] & ~t[164] & ~t[165] & t[166]) | (~t[161] & ~t[164] & ~t[165] & t[166] & ~t[167]) | (~t[161] & ~t[162] & ~t[163] & t[166] & ~t[167]) | (~t[162] & t[163] & ~t[164] & t[165] & t[166]) | (t[163] & ~t[165] & t[166] & ~t[167]);
  assign t[128] = (t[168] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (t[168] & ~t[169] & ~t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[169] & ~t[170] & ~t[173] & ~t[174]) | (~t[168] & t[169] & t[170] & t[171] & ~t[174]) | (~t[168] & t[169] & t[172] & t[173] & ~t[174]) | (t[168] & ~t[170] & ~t[172] & t[174]) | (~t[168] & t[170] & t[172] & t[174]);
  assign t[129] = (t[168] & t[169] & ~t[170] & t[171] & ~t[172] & ~t[174]) | (t[168] & ~t[170] & ~t[171] & t[172] & ~t[173] & t[174]) | (~t[169] & t[170] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[169] & t[170] & ~t[173] & ~t[174]) | (~t[168] & t[170] & t[171] & ~t[172] & t[173]) | (t[170] & ~t[171] & t[173] & ~t[174]);
  assign t[12] = ~t[21];
  assign t[130] = (t[168] & t[169] & ~t[170] & ~t[172] & t[173] & ~t[174]) | (t[168] & t[170] & ~t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & t[172] & ~t[173] & ~t[174]) | (~t[168] & ~t[170] & ~t[171] & t[172] & ~t[173]) | (~t[168] & ~t[169] & ~t[171] & t[172] & ~t[174]) | (~t[168] & ~t[170] & t[171] & t[172] & t[173]) | (t[171] & t[172] & ~t[173] & ~t[174]);
  assign t[131] = (t[169] & ~t[170] & ~t[171] & ~t[172] & ~t[173]) | (~t[168] & t[169] & ~t[171] & ~t[172] & ~t[174]) | (~t[168] & t[169] & ~t[170] & ~t[173] & ~t[174]) | (t[168] & ~t[169] & t[170] & t[171] & ~t[174]) | (t[168] & ~t[169] & t[172] & t[173] & ~t[174]) | (t[169] & ~t[171] & ~t[173] & t[174]) | (~t[169] & t[171] & t[173] & t[174]);
  assign t[132] = (t[168] & t[169] & t[170] & ~t[171] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & ~t[171] & ~t[172] & t[173] & t[174]) | (~t[169] & ~t[170] & t[171] & ~t[172] & ~t[173]) | (~t[168] & ~t[170] & t[171] & ~t[173] & ~t[174]) | (~t[168] & ~t[169] & t[171] & ~t[172] & ~t[174]) | (~t[169] & t[170] & t[171] & t[172] & ~t[173]) | (~t[170] & t[171] & t[172] & ~t[174]);
  assign t[133] = (t[168] & t[169] & ~t[171] & t[172] & ~t[173] & ~t[174]) | (t[169] & ~t[170] & t[171] & ~t[172] & ~t[173] & t[174]) | (~t[169] & ~t[170] & ~t[171] & ~t[172] & t[173]) | (~t[168] & ~t[171] & ~t[172] & t[173] & ~t[174]) | (~t[168] & ~t[169] & ~t[170] & t[173] & ~t[174]) | (~t[169] & t[170] & ~t[171] & t[172] & t[173]) | (t[170] & ~t[172] & t[173] & ~t[174]);
  assign t[134] = (t[141] & ~t[142] & ~t[143] & ~t[144] & ~t[145]) | (~t[140] & t[141] & ~t[143] & ~t[144] & ~t[146]) | (~t[140] & t[141] & ~t[142] & ~t[145] & ~t[146]) | (t[140] & ~t[141] & t[142] & t[143] & ~t[146]) | (t[140] & ~t[141] & t[144] & t[145] & ~t[146]) | (t[141] & ~t[143] & ~t[145] & t[146]) | (~t[141] & t[143] & t[145] & t[146]);
  assign t[135] = (t[140] & t[141] & t[142] & ~t[143] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[143] & ~t[144] & t[145] & t[146]) | (~t[141] & ~t[142] & t[143] & ~t[144] & ~t[145]) | (~t[140] & ~t[142] & t[143] & ~t[145] & ~t[146]) | (~t[140] & ~t[141] & t[143] & ~t[144] & ~t[146]) | (~t[141] & t[142] & t[143] & t[144] & ~t[145]) | (~t[142] & t[143] & t[144] & ~t[146]);
  assign t[136] = (t[140] & t[141] & ~t[142] & ~t[144] & t[145] & ~t[146]) | (t[140] & t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[146]) | (~t[140] & ~t[142] & ~t[143] & t[144] & ~t[145]) | (~t[140] & ~t[141] & ~t[143] & t[144] & ~t[146]) | (~t[140] & ~t[142] & t[143] & t[144] & t[145]) | (t[143] & t[144] & ~t[145] & ~t[146]);
  assign t[137] = (t[140] & t[141] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[142] & ~t[143] & ~t[144] & t[145]) | (~t[140] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[140] & ~t[141] & ~t[142] & t[145] & ~t[146]) | (~t[141] & t[142] & ~t[143] & t[144] & t[145]) | (t[142] & ~t[144] & t[145] & ~t[146]);
  assign t[138] = (t[175] & ~t[177] & ~t[178] & ~t[179] & ~t[180]) | (t[175] & ~t[176] & ~t[178] & ~t[179] & ~t[181]) | (t[175] & ~t[176] & ~t[177] & ~t[180] & ~t[181]) | (~t[175] & t[176] & t[177] & t[178] & ~t[181]) | (~t[175] & t[176] & t[179] & t[180] & ~t[181]) | (t[175] & ~t[177] & ~t[179] & t[181]) | (~t[175] & t[177] & t[179] & t[181]);
  assign t[139] = (t[175] & t[176] & ~t[177] & ~t[179] & t[180] & ~t[181]) | (t[175] & t[177] & ~t[178] & ~t[179] & ~t[180] & t[181]) | (~t[176] & ~t[177] & t[179] & ~t[180] & ~t[181]) | (~t[175] & ~t[177] & ~t[178] & t[179] & ~t[180]) | (~t[175] & ~t[176] & ~t[178] & t[179] & ~t[181]) | (~t[175] & ~t[177] & t[178] & t[179] & t[180]) | (t[178] & t[179] & ~t[180] & ~t[181]);
  assign t[13] = t[22] ^ t[23];
  assign t[140] = t[182] ^ x[7];
  assign t[141] = t[183] ^ x[51];
  assign t[142] = t[184] ^ x[8];
  assign t[143] = t[185] ^ x[52];
  assign t[144] = t[186] ^ x[53];
  assign t[145] = t[187] ^ x[54];
  assign t[146] = t[188] ^ x[6];
  assign t[147] = t[189] ^ x[15];
  assign t[148] = t[190] ^ x[10];
  assign t[149] = t[191] ^ x[11];
  assign t[14] = t[24] & t[25];
  assign t[150] = t[192] ^ x[12];
  assign t[151] = t[193] ^ x[16];
  assign t[152] = t[194] ^ x[13];
  assign t[153] = t[195] ^ x[14];
  assign t[154] = t[196] ^ x[22];
  assign t[155] = t[197] ^ x[32];
  assign t[156] = t[198] ^ x[23];
  assign t[157] = t[199] ^ x[33];
  assign t[158] = t[200] ^ x[31];
  assign t[159] = t[201] ^ x[34];
  assign t[15] = t[26] ^ t[14];
  assign t[160] = t[202] ^ x[21];
  assign t[161] = t[203] ^ x[29];
  assign t[162] = t[204] ^ x[36];
  assign t[163] = t[205] ^ x[30];
  assign t[164] = t[206] ^ x[37];
  assign t[165] = t[207] ^ x[35];
  assign t[166] = t[208] ^ x[38];
  assign t[167] = t[209] ^ x[28];
  assign t[168] = t[210] ^ x[44];
  assign t[169] = t[211] ^ x[47];
  assign t[16] = t[70] ^ t[24];
  assign t[170] = t[212] ^ x[45];
  assign t[171] = t[213] ^ x[48];
  assign t[172] = t[214] ^ x[46];
  assign t[173] = t[215] ^ x[49];
  assign t[174] = t[216] ^ x[43];
  assign t[175] = t[217] ^ x[61];
  assign t[176] = t[218] ^ x[56];
  assign t[177] = t[219] ^ x[57];
  assign t[178] = t[220] ^ x[58];
  assign t[179] = t[221] ^ x[62];
  assign t[17] = t[27] ^ t[28];
  assign t[180] = t[222] ^ x[59];
  assign t[181] = t[223] ^ x[60];
  assign t[182] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[183] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[184] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[185] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[186] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[187] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[188] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[189] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[18] = t[29] & t[30];
  assign t[190] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[191] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[192] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[193] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[194] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[195] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[196] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[197] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[198] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[199] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[201] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[202] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[203] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[204] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[205] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[206] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[207] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[208] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[209] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[20] = t[71] ^ t[29];
  assign t[210] = (x[39] & ~x[40] & ~x[41]) | (~x[39] & x[40] & ~x[41]) | (~x[39] & ~x[40] & x[41]) | (x[39] & x[40] & x[41]);
  assign t[211] = (x[39] & ~x[40] & ~x[42]) | (~x[39] & x[40] & ~x[42]) | (~x[39] & ~x[40] & x[42]) | (x[39] & x[40] & x[42]);
  assign t[212] = (x[39] & ~x[41]) | (~x[39] & x[41]);
  assign t[213] = (x[39] & ~x[42]) | (~x[39] & x[42]);
  assign t[214] = (x[40] & ~x[41]) | (~x[40] & x[41]);
  assign t[215] = (x[40] & ~x[42]) | (~x[40] & x[42]);
  assign t[216] = (x[41] & ~x[42]) | (~x[41] & x[42]);
  assign t[217] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[218] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[219] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[220] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[221] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[222] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[223] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[22] = t[72] ^ t[73];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[73]);
  assign t[25] = ~(t[70] ^ t[24]);
  assign t[26] = t[70] & t[35];
  assign t[27] = t[74] ^ t[75];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[75]);
  assign t[2] = ~(t[4] ^ t[68]);
  assign t[30] = ~(t[71] ^ t[29]);
  assign t[31] = t[71] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[70] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[71] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[76] ^ t[48];
  assign t[42] = t[73] ^ t[77];
  assign t[43] = t[70] ^ t[22];
  assign t[44] = t[75] ^ t[78];
  assign t[45] = t[71] ^ t[27];
  assign t[46] = t[79] ^ t[80];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[80]);
  assign t[49] = ~(t[76] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[76] & t[52];
  assign t[51] = t[76] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[80] ^ t[81];
  assign t[54] = t[76] ^ t[46];
  assign t[55] = x[0] ? x[50] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[82]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = ~(t[63]);
  assign t[61] = ~(t[64]);
  assign t[62] = ~(t[65] ^ t[83]);
  assign t[63] = t[42] ^ t[14];
  assign t[64] = t[44] ^ t[18];
  assign t[65] = ~t[66];
  assign t[66] = ~(t[67]);
  assign t[67] = t[53] ^ t[39];
  assign t[68] = (t[84] & ~t[85]) | (~t[84] & t[85]);
  assign t[69] = (t[86] & ~t[87]) | (~t[86] & t[87]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (t[88] & ~t[89]) | (~t[88] & t[89]);
  assign t[71] = (t[90] & ~t[91]) | (~t[90] & t[91]);
  assign t[72] = (t[88] & ~t[92]) | (~t[88] & t[92]);
  assign t[73] = (t[88] & ~t[94] & ~t[95]) | (~t[93] & t[94] & ~t[92]) | (~t[88] & ~t[94] & t[95]) | (t[93] & t[94] & t[92]);
  assign t[74] = (t[90] & ~t[96]) | (~t[90] & t[96]);
  assign t[75] = (t[90] & ~t[98] & ~t[99]) | (~t[97] & t[98] & ~t[96]) | (~t[90] & ~t[98] & t[99]) | (t[97] & t[98] & t[96]);
  assign t[76] = (t[100] & ~t[101]) | (~t[100] & t[101]);
  assign t[77] = (t[88] & ~t[94] & ~t[92]) | (~t[93] & t[94] & ~t[95]) | (~t[88] & ~t[94] & t[92]) | (t[93] & t[94] & t[95]);
  assign t[78] = (t[90] & ~t[98] & ~t[96]) | (~t[97] & t[98] & ~t[99]) | (~t[90] & ~t[98] & t[96]) | (t[97] & t[98] & t[99]);
  assign t[79] = (t[100] & ~t[102]) | (~t[100] & t[102]);
  assign t[7] = ~(t[12] ^ t[69]);
  assign t[80] = (t[100] & ~t[104] & ~t[105]) | (~t[103] & t[104] & ~t[102]) | (~t[100] & ~t[104] & t[105]) | (t[103] & t[104] & t[102]);
  assign t[81] = (t[100] & ~t[104] & ~t[102]) | (~t[103] & t[104] & ~t[105]) | (~t[100] & ~t[104] & t[102]) | (t[103] & t[104] & t[105]);
  assign t[82] = (t[84] & ~t[107] & ~t[109]) | (~t[106] & t[107] & ~t[108]) | (~t[84] & ~t[107] & t[109]) | (t[106] & t[107] & t[108]);
  assign t[83] = (t[110] & ~t[111]) | (~t[110] & t[111]);
  assign t[84] = t[112] ^ x[7];
  assign t[85] = t[113] ^ x[8];
  assign t[86] = t[114] ^ x[15];
  assign t[87] = t[115] ^ x[16];
  assign t[88] = t[116] ^ x[22];
  assign t[89] = t[117] ^ x[23];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[118] ^ x[29];
  assign t[91] = t[119] ^ x[30];
  assign t[92] = t[120] ^ x[31];
  assign t[93] = t[121] ^ x[32];
  assign t[94] = t[122] ^ x[33];
  assign t[95] = t[123] ^ x[34];
  assign t[96] = t[124] ^ x[35];
  assign t[97] = t[125] ^ x[36];
  assign t[98] = t[126] ^ x[37];
  assign t[99] = t[127] ^ x[38];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0] & ~t[55]) | (~t[0] & t[55]);
endmodule

module R2ind166(x, y);
 input [62:0] x;
 output y;

 wire [220:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = t[128] ^ x[47];
  assign t[101] = t[129] ^ x[48];
  assign t[102] = t[130] ^ x[49];
  assign t[103] = t[131] ^ x[51];
  assign t[104] = t[132] ^ x[52];
  assign t[105] = t[133] ^ x[53];
  assign t[106] = t[134] ^ x[54];
  assign t[107] = t[135] ^ x[61];
  assign t[108] = t[136] ^ x[62];
  assign t[109] = (t[137] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (t[137] & ~t[138] & ~t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[138] & ~t[139] & ~t[142] & ~t[143]) | (~t[137] & t[138] & t[139] & t[140] & ~t[143]) | (~t[137] & t[138] & t[141] & t[142] & ~t[143]) | (t[137] & ~t[139] & ~t[141] & t[143]) | (~t[137] & t[139] & t[141] & t[143]);
  assign t[10] = t[17] ^ t[18];
  assign t[110] = (t[137] & t[138] & ~t[139] & t[140] & ~t[141] & ~t[143]) | (t[137] & ~t[139] & ~t[140] & t[141] & ~t[142] & t[143]) | (~t[138] & t[139] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[138] & t[139] & ~t[142] & ~t[143]) | (~t[137] & t[139] & t[140] & ~t[141] & t[142]) | (t[139] & ~t[140] & t[142] & ~t[143]);
  assign t[111] = (t[144] & ~t[146] & ~t[147] & ~t[148] & ~t[149]) | (t[144] & ~t[145] & ~t[147] & ~t[148] & ~t[150]) | (t[144] & ~t[145] & ~t[146] & ~t[149] & ~t[150]) | (~t[144] & t[145] & t[146] & t[147] & ~t[150]) | (~t[144] & t[145] & t[148] & t[149] & ~t[150]) | (t[144] & ~t[146] & ~t[148] & t[150]) | (~t[144] & t[146] & t[148] & t[150]);
  assign t[112] = (t[144] & t[145] & ~t[146] & ~t[148] & t[149] & ~t[150]) | (t[144] & t[146] & ~t[147] & ~t[148] & ~t[149] & t[150]) | (~t[145] & ~t[146] & t[148] & ~t[149] & ~t[150]) | (~t[144] & ~t[146] & ~t[147] & t[148] & ~t[149]) | (~t[144] & ~t[145] & ~t[147] & t[148] & ~t[150]) | (~t[144] & ~t[146] & t[147] & t[148] & t[149]) | (t[147] & t[148] & ~t[149] & ~t[150]);
  assign t[113] = (t[151] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (t[151] & ~t[152] & ~t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[152] & ~t[153] & ~t[156] & ~t[157]) | (~t[151] & t[152] & t[153] & t[154] & ~t[157]) | (~t[151] & t[152] & t[155] & t[156] & ~t[157]) | (t[151] & ~t[153] & ~t[155] & t[157]) | (~t[151] & t[153] & t[155] & t[157]);
  assign t[114] = (t[151] & t[152] & ~t[153] & t[154] & ~t[155] & ~t[157]) | (t[151] & ~t[153] & ~t[154] & t[155] & ~t[156] & t[157]) | (~t[152] & t[153] & ~t[154] & ~t[155] & ~t[157]) | (~t[151] & t[153] & ~t[154] & ~t[155] & ~t[156]) | (~t[151] & ~t[152] & t[153] & ~t[156] & ~t[157]) | (~t[151] & t[153] & t[154] & ~t[155] & t[156]) | (t[153] & ~t[154] & t[156] & ~t[157]);
  assign t[115] = (t[158] & ~t[160] & ~t[161] & ~t[162] & ~t[163]) | (t[158] & ~t[159] & ~t[161] & ~t[162] & ~t[164]) | (t[158] & ~t[159] & ~t[160] & ~t[163] & ~t[164]) | (~t[158] & t[159] & t[160] & t[161] & ~t[164]) | (~t[158] & t[159] & t[162] & t[163] & ~t[164]) | (t[158] & ~t[160] & ~t[162] & t[164]) | (~t[158] & t[160] & t[162] & t[164]);
  assign t[116] = (t[158] & t[159] & ~t[160] & t[161] & ~t[162] & ~t[164]) | (t[158] & ~t[160] & ~t[161] & t[162] & ~t[163] & t[164]) | (~t[159] & t[160] & ~t[161] & ~t[162] & ~t[164]) | (~t[158] & t[160] & ~t[161] & ~t[162] & ~t[163]) | (~t[158] & ~t[159] & t[160] & ~t[163] & ~t[164]) | (~t[158] & t[160] & t[161] & ~t[162] & t[163]) | (t[160] & ~t[161] & t[163] & ~t[164]);
  assign t[117] = (t[151] & t[152] & ~t[153] & ~t[155] & t[156] & ~t[157]) | (t[151] & t[153] & ~t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & t[155] & ~t[156] & ~t[157]) | (~t[151] & ~t[153] & ~t[154] & t[155] & ~t[156]) | (~t[151] & ~t[152] & ~t[154] & t[155] & ~t[157]) | (~t[151] & ~t[153] & t[154] & t[155] & t[156]) | (t[154] & t[155] & ~t[156] & ~t[157]);
  assign t[118] = (t[152] & ~t[153] & ~t[154] & ~t[155] & ~t[156]) | (~t[151] & t[152] & ~t[154] & ~t[155] & ~t[157]) | (~t[151] & t[152] & ~t[153] & ~t[156] & ~t[157]) | (t[151] & ~t[152] & t[153] & t[154] & ~t[157]) | (t[151] & ~t[152] & t[155] & t[156] & ~t[157]) | (t[152] & ~t[154] & ~t[156] & t[157]) | (~t[152] & t[154] & t[156] & t[157]);
  assign t[119] = (t[151] & t[152] & t[153] & ~t[154] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & ~t[154] & ~t[155] & t[156] & t[157]) | (~t[152] & ~t[153] & t[154] & ~t[155] & ~t[156]) | (~t[151] & ~t[153] & t[154] & ~t[156] & ~t[157]) | (~t[151] & ~t[152] & t[154] & ~t[155] & ~t[157]) | (~t[152] & t[153] & t[154] & t[155] & ~t[156]) | (~t[153] & t[154] & t[155] & ~t[157]);
  assign t[11] = t[19] ^ t[20];
  assign t[120] = (t[151] & t[152] & ~t[154] & t[155] & ~t[156] & ~t[157]) | (t[152] & ~t[153] & t[154] & ~t[155] & ~t[156] & t[157]) | (~t[152] & ~t[153] & ~t[154] & ~t[155] & t[156]) | (~t[151] & ~t[154] & ~t[155] & t[156] & ~t[157]) | (~t[151] & ~t[152] & ~t[153] & t[156] & ~t[157]) | (~t[152] & t[153] & ~t[154] & t[155] & t[156]) | (t[153] & ~t[155] & t[156] & ~t[157]);
  assign t[121] = (t[158] & t[159] & ~t[160] & ~t[162] & t[163] & ~t[164]) | (t[158] & t[160] & ~t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[160] & t[162] & ~t[163] & ~t[164]) | (~t[158] & ~t[160] & ~t[161] & t[162] & ~t[163]) | (~t[158] & ~t[159] & ~t[161] & t[162] & ~t[164]) | (~t[158] & ~t[160] & t[161] & t[162] & t[163]) | (t[161] & t[162] & ~t[163] & ~t[164]);
  assign t[122] = (t[159] & ~t[160] & ~t[161] & ~t[162] & ~t[163]) | (~t[158] & t[159] & ~t[161] & ~t[162] & ~t[164]) | (~t[158] & t[159] & ~t[160] & ~t[163] & ~t[164]) | (t[158] & ~t[159] & t[160] & t[161] & ~t[164]) | (t[158] & ~t[159] & t[162] & t[163] & ~t[164]) | (t[159] & ~t[161] & ~t[163] & t[164]) | (~t[159] & t[161] & t[163] & t[164]);
  assign t[123] = (t[158] & t[159] & t[160] & ~t[161] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & ~t[161] & ~t[162] & t[163] & t[164]) | (~t[159] & ~t[160] & t[161] & ~t[162] & ~t[163]) | (~t[158] & ~t[160] & t[161] & ~t[163] & ~t[164]) | (~t[158] & ~t[159] & t[161] & ~t[162] & ~t[164]) | (~t[159] & t[160] & t[161] & t[162] & ~t[163]) | (~t[160] & t[161] & t[162] & ~t[164]);
  assign t[124] = (t[158] & t[159] & ~t[161] & t[162] & ~t[163] & ~t[164]) | (t[159] & ~t[160] & t[161] & ~t[162] & ~t[163] & t[164]) | (~t[159] & ~t[160] & ~t[161] & ~t[162] & t[163]) | (~t[158] & ~t[161] & ~t[162] & t[163] & ~t[164]) | (~t[158] & ~t[159] & ~t[160] & t[163] & ~t[164]) | (~t[159] & t[160] & ~t[161] & t[162] & t[163]) | (t[160] & ~t[162] & t[163] & ~t[164]);
  assign t[125] = (t[165] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (t[165] & ~t[166] & ~t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[166] & ~t[167] & ~t[170] & ~t[171]) | (~t[165] & t[166] & t[167] & t[168] & ~t[171]) | (~t[165] & t[166] & t[169] & t[170] & ~t[171]) | (t[165] & ~t[167] & ~t[169] & t[171]) | (~t[165] & t[167] & t[169] & t[171]);
  assign t[126] = (t[165] & t[166] & ~t[167] & t[168] & ~t[169] & ~t[171]) | (t[165] & ~t[167] & ~t[168] & t[169] & ~t[170] & t[171]) | (~t[166] & t[167] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[166] & t[167] & ~t[170] & ~t[171]) | (~t[165] & t[167] & t[168] & ~t[169] & t[170]) | (t[167] & ~t[168] & t[170] & ~t[171]);
  assign t[127] = (t[165] & t[166] & ~t[167] & ~t[169] & t[170] & ~t[171]) | (t[165] & t[167] & ~t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & t[169] & ~t[170] & ~t[171]) | (~t[165] & ~t[167] & ~t[168] & t[169] & ~t[170]) | (~t[165] & ~t[166] & ~t[168] & t[169] & ~t[171]) | (~t[165] & ~t[167] & t[168] & t[169] & t[170]) | (t[168] & t[169] & ~t[170] & ~t[171]);
  assign t[128] = (t[166] & ~t[167] & ~t[168] & ~t[169] & ~t[170]) | (~t[165] & t[166] & ~t[168] & ~t[169] & ~t[171]) | (~t[165] & t[166] & ~t[167] & ~t[170] & ~t[171]) | (t[165] & ~t[166] & t[167] & t[168] & ~t[171]) | (t[165] & ~t[166] & t[169] & t[170] & ~t[171]) | (t[166] & ~t[168] & ~t[170] & t[171]) | (~t[166] & t[168] & t[170] & t[171]);
  assign t[129] = (t[165] & t[166] & t[167] & ~t[168] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & ~t[168] & ~t[169] & t[170] & t[171]) | (~t[166] & ~t[167] & t[168] & ~t[169] & ~t[170]) | (~t[165] & ~t[167] & t[168] & ~t[170] & ~t[171]) | (~t[165] & ~t[166] & t[168] & ~t[169] & ~t[171]) | (~t[166] & t[167] & t[168] & t[169] & ~t[170]) | (~t[167] & t[168] & t[169] & ~t[171]);
  assign t[12] = ~t[21];
  assign t[130] = (t[165] & t[166] & ~t[168] & t[169] & ~t[170] & ~t[171]) | (t[166] & ~t[167] & t[168] & ~t[169] & ~t[170] & t[171]) | (~t[166] & ~t[167] & ~t[168] & ~t[169] & t[170]) | (~t[165] & ~t[168] & ~t[169] & t[170] & ~t[171]) | (~t[165] & ~t[166] & ~t[167] & t[170] & ~t[171]) | (~t[166] & t[167] & ~t[168] & t[169] & t[170]) | (t[167] & ~t[169] & t[170] & ~t[171]);
  assign t[131] = (t[138] & ~t[139] & ~t[140] & ~t[141] & ~t[142]) | (~t[137] & t[138] & ~t[140] & ~t[141] & ~t[143]) | (~t[137] & t[138] & ~t[139] & ~t[142] & ~t[143]) | (t[137] & ~t[138] & t[139] & t[140] & ~t[143]) | (t[137] & ~t[138] & t[141] & t[142] & ~t[143]) | (t[138] & ~t[140] & ~t[142] & t[143]) | (~t[138] & t[140] & t[142] & t[143]);
  assign t[132] = (t[137] & t[138] & t[139] & ~t[140] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & ~t[140] & ~t[141] & t[142] & t[143]) | (~t[138] & ~t[139] & t[140] & ~t[141] & ~t[142]) | (~t[137] & ~t[139] & t[140] & ~t[142] & ~t[143]) | (~t[137] & ~t[138] & t[140] & ~t[141] & ~t[143]) | (~t[138] & t[139] & t[140] & t[141] & ~t[142]) | (~t[139] & t[140] & t[141] & ~t[143]);
  assign t[133] = (t[137] & t[138] & ~t[139] & ~t[141] & t[142] & ~t[143]) | (t[137] & t[139] & ~t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & t[141] & ~t[142] & ~t[143]) | (~t[137] & ~t[139] & ~t[140] & t[141] & ~t[142]) | (~t[137] & ~t[138] & ~t[140] & t[141] & ~t[143]) | (~t[137] & ~t[139] & t[140] & t[141] & t[142]) | (t[140] & t[141] & ~t[142] & ~t[143]);
  assign t[134] = (t[137] & t[138] & ~t[140] & t[141] & ~t[142] & ~t[143]) | (t[138] & ~t[139] & t[140] & ~t[141] & ~t[142] & t[143]) | (~t[138] & ~t[139] & ~t[140] & ~t[141] & t[142]) | (~t[137] & ~t[140] & ~t[141] & t[142] & ~t[143]) | (~t[137] & ~t[138] & ~t[139] & t[142] & ~t[143]) | (~t[138] & t[139] & ~t[140] & t[141] & t[142]) | (t[139] & ~t[141] & t[142] & ~t[143]);
  assign t[135] = (t[172] & ~t[174] & ~t[175] & ~t[176] & ~t[177]) | (t[172] & ~t[173] & ~t[175] & ~t[176] & ~t[178]) | (t[172] & ~t[173] & ~t[174] & ~t[177] & ~t[178]) | (~t[172] & t[173] & t[174] & t[175] & ~t[178]) | (~t[172] & t[173] & t[176] & t[177] & ~t[178]) | (t[172] & ~t[174] & ~t[176] & t[178]) | (~t[172] & t[174] & t[176] & t[178]);
  assign t[136] = (t[172] & t[173] & ~t[174] & ~t[176] & t[177] & ~t[178]) | (t[172] & t[174] & ~t[175] & ~t[176] & ~t[177] & t[178]) | (~t[173] & ~t[174] & t[176] & ~t[177] & ~t[178]) | (~t[172] & ~t[174] & ~t[175] & t[176] & ~t[177]) | (~t[172] & ~t[173] & ~t[175] & t[176] & ~t[178]) | (~t[172] & ~t[174] & t[175] & t[176] & t[177]) | (t[175] & t[176] & ~t[177] & ~t[178]);
  assign t[137] = t[179] ^ x[7];
  assign t[138] = t[180] ^ x[51];
  assign t[139] = t[181] ^ x[8];
  assign t[13] = t[22] ^ t[23];
  assign t[140] = t[182] ^ x[52];
  assign t[141] = t[183] ^ x[53];
  assign t[142] = t[184] ^ x[54];
  assign t[143] = t[185] ^ x[6];
  assign t[144] = t[186] ^ x[15];
  assign t[145] = t[187] ^ x[10];
  assign t[146] = t[188] ^ x[11];
  assign t[147] = t[189] ^ x[12];
  assign t[148] = t[190] ^ x[16];
  assign t[149] = t[191] ^ x[13];
  assign t[14] = t[24] & t[25];
  assign t[150] = t[192] ^ x[14];
  assign t[151] = t[193] ^ x[22];
  assign t[152] = t[194] ^ x[32];
  assign t[153] = t[195] ^ x[23];
  assign t[154] = t[196] ^ x[33];
  assign t[155] = t[197] ^ x[31];
  assign t[156] = t[198] ^ x[34];
  assign t[157] = t[199] ^ x[21];
  assign t[158] = t[200] ^ x[29];
  assign t[159] = t[201] ^ x[36];
  assign t[15] = t[26] ^ t[14];
  assign t[160] = t[202] ^ x[30];
  assign t[161] = t[203] ^ x[37];
  assign t[162] = t[204] ^ x[35];
  assign t[163] = t[205] ^ x[38];
  assign t[164] = t[206] ^ x[28];
  assign t[165] = t[207] ^ x[44];
  assign t[166] = t[208] ^ x[47];
  assign t[167] = t[209] ^ x[45];
  assign t[168] = t[210] ^ x[48];
  assign t[169] = t[211] ^ x[46];
  assign t[16] = t[67] ^ t[24];
  assign t[170] = t[212] ^ x[49];
  assign t[171] = t[213] ^ x[43];
  assign t[172] = t[214] ^ x[61];
  assign t[173] = t[215] ^ x[56];
  assign t[174] = t[216] ^ x[57];
  assign t[175] = t[217] ^ x[58];
  assign t[176] = t[218] ^ x[62];
  assign t[177] = t[219] ^ x[59];
  assign t[178] = t[220] ^ x[60];
  assign t[179] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[17] = t[27] ^ t[28];
  assign t[180] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[181] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[182] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[183] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[184] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[185] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[186] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[187] = (x[9] & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0);
  assign t[188] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[189] = (x[9] & ~1'b0) | (~x[9] & 1'b0);
  assign t[18] = t[29] & t[30];
  assign t[190] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[191] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[192] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[193] = (x[17] & ~x[18] & ~x[19]) | (~x[17] & x[18] & ~x[19]) | (~x[17] & ~x[18] & x[19]) | (x[17] & x[18] & x[19]);
  assign t[194] = (x[17] & ~x[18] & ~x[20]) | (~x[17] & x[18] & ~x[20]) | (~x[17] & ~x[18] & x[20]) | (x[17] & x[18] & x[20]);
  assign t[195] = (x[17] & ~x[19]) | (~x[17] & x[19]);
  assign t[196] = (x[17] & ~x[20]) | (~x[17] & x[20]);
  assign t[197] = (x[18] & ~x[19]) | (~x[18] & x[19]);
  assign t[198] = (x[18] & ~x[20]) | (~x[18] & x[20]);
  assign t[199] = (x[19] & ~x[20]) | (~x[19] & x[20]);
  assign t[19] = t[31] ^ t[18];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[24] & ~x[25] & ~x[26]) | (~x[24] & x[25] & ~x[26]) | (~x[24] & ~x[25] & x[26]) | (x[24] & x[25] & x[26]);
  assign t[201] = (x[24] & ~x[25] & ~x[27]) | (~x[24] & x[25] & ~x[27]) | (~x[24] & ~x[25] & x[27]) | (x[24] & x[25] & x[27]);
  assign t[202] = (x[24] & ~x[26]) | (~x[24] & x[26]);
  assign t[203] = (x[24] & ~x[27]) | (~x[24] & x[27]);
  assign t[204] = (x[25] & ~x[26]) | (~x[25] & x[26]);
  assign t[205] = (x[25] & ~x[27]) | (~x[25] & x[27]);
  assign t[206] = (x[26] & ~x[27]) | (~x[26] & x[27]);
  assign t[207] = (x[39] & ~x[40] & ~x[41]) | (~x[39] & x[40] & ~x[41]) | (~x[39] & ~x[40] & x[41]) | (x[39] & x[40] & x[41]);
  assign t[208] = (x[39] & ~x[40] & ~x[42]) | (~x[39] & x[40] & ~x[42]) | (~x[39] & ~x[40] & x[42]) | (x[39] & x[40] & x[42]);
  assign t[209] = (x[39] & ~x[41]) | (~x[39] & x[41]);
  assign t[20] = t[68] ^ t[29];
  assign t[210] = (x[39] & ~x[42]) | (~x[39] & x[42]);
  assign t[211] = (x[40] & ~x[41]) | (~x[40] & x[41]);
  assign t[212] = (x[40] & ~x[42]) | (~x[40] & x[42]);
  assign t[213] = (x[41] & ~x[42]) | (~x[41] & x[42]);
  assign t[214] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[215] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[216] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[217] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[218] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[219] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[21] = ~(t[32] ^ t[33]);
  assign t[220] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[22] = t[69] ^ t[70];
  assign t[23] = t[24] & t[34];
  assign t[24] = ~(t[70]);
  assign t[25] = ~(t[67] ^ t[24]);
  assign t[26] = t[67] & t[35];
  assign t[27] = t[71] ^ t[72];
  assign t[28] = t[29] & t[36];
  assign t[29] = ~(t[72]);
  assign t[2] = ~(t[4] ^ t[65]);
  assign t[30] = ~(t[68] ^ t[29]);
  assign t[31] = t[68] & t[37];
  assign t[32] = t[38] ^ t[39];
  assign t[33] = t[40] ^ t[41];
  assign t[34] = t[67] ^ t[42];
  assign t[35] = t[43] ^ t[23];
  assign t[36] = t[68] ^ t[44];
  assign t[37] = t[45] ^ t[28];
  assign t[38] = t[46] ^ t[47];
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[50] ^ t[39];
  assign t[41] = t[73] ^ t[48];
  assign t[42] = t[70] ^ t[74];
  assign t[43] = t[67] ^ t[22];
  assign t[44] = t[72] ^ t[75];
  assign t[45] = t[68] ^ t[27];
  assign t[46] = t[76] ^ t[77];
  assign t[47] = t[48] & t[51];
  assign t[48] = ~(t[77]);
  assign t[49] = ~(t[73] ^ t[48]);
  assign t[4] = ~t[7];
  assign t[50] = t[73] & t[52];
  assign t[51] = t[73] ^ t[53];
  assign t[52] = t[54] ^ t[47];
  assign t[53] = t[77] ^ t[78];
  assign t[54] = t[73] ^ t[46];
  assign t[55] = x[0] ? x[50] : t[56];
  assign t[56] = ~(t[57] ^ t[58]);
  assign t[57] = ~(t[59] ^ t[79]);
  assign t[58] = ~(t[60] ^ t[61]);
  assign t[59] = ~t[62];
  assign t[5] = ~(t[8] ^ t[9]);
  assign t[60] = ~(t[8]);
  assign t[61] = ~(t[10]);
  assign t[62] = ~(t[63] ^ t[80]);
  assign t[63] = ~t[64];
  assign t[64] = ~(t[32]);
  assign t[65] = (t[81] & ~t[82]) | (~t[81] & t[82]);
  assign t[66] = (t[83] & ~t[84]) | (~t[83] & t[84]);
  assign t[67] = (t[85] & ~t[86]) | (~t[85] & t[86]);
  assign t[68] = (t[87] & ~t[88]) | (~t[87] & t[88]);
  assign t[69] = (t[85] & ~t[89]) | (~t[85] & t[89]);
  assign t[6] = ~(t[10] ^ t[11]);
  assign t[70] = (t[85] & ~t[91] & ~t[92]) | (~t[90] & t[91] & ~t[89]) | (~t[85] & ~t[91] & t[92]) | (t[90] & t[91] & t[89]);
  assign t[71] = (t[87] & ~t[93]) | (~t[87] & t[93]);
  assign t[72] = (t[87] & ~t[95] & ~t[96]) | (~t[94] & t[95] & ~t[93]) | (~t[87] & ~t[95] & t[96]) | (t[94] & t[95] & t[93]);
  assign t[73] = (t[97] & ~t[98]) | (~t[97] & t[98]);
  assign t[74] = (t[85] & ~t[91] & ~t[89]) | (~t[90] & t[91] & ~t[92]) | (~t[85] & ~t[91] & t[89]) | (t[90] & t[91] & t[92]);
  assign t[75] = (t[87] & ~t[95] & ~t[93]) | (~t[94] & t[95] & ~t[96]) | (~t[87] & ~t[95] & t[93]) | (t[94] & t[95] & t[96]);
  assign t[76] = (t[97] & ~t[99]) | (~t[97] & t[99]);
  assign t[77] = (t[97] & ~t[101] & ~t[102]) | (~t[100] & t[101] & ~t[99]) | (~t[97] & ~t[101] & t[102]) | (t[100] & t[101] & t[99]);
  assign t[78] = (t[97] & ~t[101] & ~t[99]) | (~t[100] & t[101] & ~t[102]) | (~t[97] & ~t[101] & t[99]) | (t[100] & t[101] & t[102]);
  assign t[79] = (t[81] & ~t[104] & ~t[105]) | (~t[103] & t[104] & ~t[106]) | (~t[81] & ~t[104] & t[105]) | (t[103] & t[104] & t[106]);
  assign t[7] = ~(t[12] ^ t[66]);
  assign t[80] = (t[107] & ~t[108]) | (~t[107] & t[108]);
  assign t[81] = t[109] ^ x[7];
  assign t[82] = t[110] ^ x[8];
  assign t[83] = t[111] ^ x[15];
  assign t[84] = t[112] ^ x[16];
  assign t[85] = t[113] ^ x[22];
  assign t[86] = t[114] ^ x[23];
  assign t[87] = t[115] ^ x[29];
  assign t[88] = t[116] ^ x[30];
  assign t[89] = t[117] ^ x[31];
  assign t[8] = t[13] ^ t[14];
  assign t[90] = t[118] ^ x[32];
  assign t[91] = t[119] ^ x[33];
  assign t[92] = t[120] ^ x[34];
  assign t[93] = t[121] ^ x[35];
  assign t[94] = t[122] ^ x[36];
  assign t[95] = t[123] ^ x[37];
  assign t[96] = t[124] ^ x[38];
  assign t[97] = t[125] ^ x[44];
  assign t[98] = t[126] ^ x[45];
  assign t[99] = t[127] ^ x[46];
  assign t[9] = t[15] ^ t[16];
  assign y = (t[0] & ~t[55]) | (~t[0] & t[55]);
endmodule

module R2ind167(x, y);
 input [62:0] x;
 output y;

 wire [203:0] t;
  assign t[0] = x[0] ? x[1] : t[1];
  assign t[100] = (t[134] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (t[134] & ~t[135] & ~t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[135] & ~t[136] & ~t[139] & ~t[140]) | (~t[134] & t[135] & t[136] & t[137] & ~t[140]) | (~t[134] & t[135] & t[138] & t[139] & ~t[140]) | (t[134] & ~t[136] & ~t[138] & t[140]) | (~t[134] & t[136] & t[138] & t[140]);
  assign t[101] = (t[135] & ~t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & t[135] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[135] & ~t[136] & ~t[139] & ~t[140]) | (t[134] & ~t[135] & t[136] & t[137] & ~t[140]) | (t[134] & ~t[135] & t[138] & t[139] & ~t[140]) | (t[135] & ~t[137] & ~t[139] & t[140]) | (~t[135] & t[137] & t[139] & t[140]);
  assign t[102] = (t[134] & t[135] & t[136] & ~t[137] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & ~t[137] & ~t[138] & t[139] & t[140]) | (~t[135] & ~t[136] & t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[136] & t[137] & ~t[139] & ~t[140]) | (~t[134] & ~t[135] & t[137] & ~t[138] & ~t[140]) | (~t[135] & t[136] & t[137] & t[138] & ~t[139]) | (~t[136] & t[137] & t[138] & ~t[140]);
  assign t[103] = (t[134] & t[135] & ~t[136] & ~t[138] & t[139] & ~t[140]) | (t[134] & t[136] & ~t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & t[138] & ~t[139] & ~t[140]) | (~t[134] & ~t[136] & ~t[137] & t[138] & ~t[139]) | (~t[134] & ~t[135] & ~t[137] & t[138] & ~t[140]) | (~t[134] & ~t[136] & t[137] & t[138] & t[139]) | (t[137] & t[138] & ~t[139] & ~t[140]);
  assign t[104] = (t[134] & t[135] & ~t[137] & t[138] & ~t[139] & ~t[140]) | (t[135] & ~t[136] & t[137] & ~t[138] & ~t[139] & t[140]) | (~t[135] & ~t[136] & ~t[137] & ~t[138] & t[139]) | (~t[134] & ~t[137] & ~t[138] & t[139] & ~t[140]) | (~t[134] & ~t[135] & ~t[136] & t[139] & ~t[140]) | (~t[135] & t[136] & ~t[137] & t[138] & t[139]) | (t[136] & ~t[138] & t[139] & ~t[140]);
  assign t[105] = (t[141] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (t[141] & ~t[142] & ~t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[142] & ~t[143] & ~t[146] & ~t[147]) | (~t[141] & t[142] & t[143] & t[144] & ~t[147]) | (~t[141] & t[142] & t[145] & t[146] & ~t[147]) | (t[141] & ~t[143] & ~t[145] & t[147]) | (~t[141] & t[143] & t[145] & t[147]);
  assign t[106] = (t[142] & ~t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & t[142] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[142] & ~t[143] & ~t[146] & ~t[147]) | (t[141] & ~t[142] & t[143] & t[144] & ~t[147]) | (t[141] & ~t[142] & t[145] & t[146] & ~t[147]) | (t[142] & ~t[144] & ~t[146] & t[147]) | (~t[142] & t[144] & t[146] & t[147]);
  assign t[107] = (t[141] & t[142] & t[143] & ~t[144] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & ~t[144] & ~t[145] & t[146] & t[147]) | (~t[142] & ~t[143] & t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[143] & t[144] & ~t[146] & ~t[147]) | (~t[141] & ~t[142] & t[144] & ~t[145] & ~t[147]) | (~t[142] & t[143] & t[144] & t[145] & ~t[146]) | (~t[143] & t[144] & t[145] & ~t[147]);
  assign t[108] = (t[141] & t[142] & ~t[143] & ~t[145] & t[146] & ~t[147]) | (t[141] & t[143] & ~t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & t[145] & ~t[146] & ~t[147]) | (~t[141] & ~t[143] & ~t[144] & t[145] & ~t[146]) | (~t[141] & ~t[142] & ~t[144] & t[145] & ~t[147]) | (~t[141] & ~t[143] & t[144] & t[145] & t[146]) | (t[144] & t[145] & ~t[146] & ~t[147]);
  assign t[109] = (t[141] & t[142] & ~t[144] & t[145] & ~t[146] & ~t[147]) | (t[142] & ~t[143] & t[144] & ~t[145] & ~t[146] & t[147]) | (~t[142] & ~t[143] & ~t[144] & ~t[145] & t[146]) | (~t[141] & ~t[144] & ~t[145] & t[146] & ~t[147]) | (~t[141] & ~t[142] & ~t[143] & t[146] & ~t[147]) | (~t[142] & t[143] & ~t[144] & t[145] & t[146]) | (t[143] & ~t[145] & t[146] & ~t[147]);
  assign t[10] = ~t[15];
  assign t[110] = (t[134] & t[135] & ~t[136] & t[137] & ~t[138] & ~t[140]) | (t[134] & ~t[136] & ~t[137] & t[138] & ~t[139] & t[140]) | (~t[135] & t[136] & ~t[137] & ~t[138] & ~t[140]) | (~t[134] & t[136] & ~t[137] & ~t[138] & ~t[139]) | (~t[134] & ~t[135] & t[136] & ~t[139] & ~t[140]) | (~t[134] & t[136] & t[137] & ~t[138] & t[139]) | (t[136] & ~t[137] & t[139] & ~t[140]);
  assign t[111] = (t[141] & t[142] & ~t[143] & t[144] & ~t[145] & ~t[147]) | (t[141] & ~t[143] & ~t[144] & t[145] & ~t[146] & t[147]) | (~t[142] & t[143] & ~t[144] & ~t[145] & ~t[147]) | (~t[141] & t[143] & ~t[144] & ~t[145] & ~t[146]) | (~t[141] & ~t[142] & t[143] & ~t[146] & ~t[147]) | (~t[141] & t[143] & t[144] & ~t[145] & t[146]) | (t[143] & ~t[144] & t[146] & ~t[147]);
  assign t[112] = (t[148] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (t[148] & ~t[149] & ~t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[149] & ~t[150] & ~t[153] & ~t[154]) | (~t[148] & t[149] & t[150] & t[151] & ~t[154]) | (~t[148] & t[149] & t[152] & t[153] & ~t[154]) | (t[148] & ~t[150] & ~t[152] & t[154]) | (~t[148] & t[150] & t[152] & t[154]);
  assign t[113] = (t[149] & ~t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & t[149] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[149] & ~t[150] & ~t[153] & ~t[154]) | (t[148] & ~t[149] & t[150] & t[151] & ~t[154]) | (t[148] & ~t[149] & t[152] & t[153] & ~t[154]) | (t[149] & ~t[151] & ~t[153] & t[154]) | (~t[149] & t[151] & t[153] & t[154]);
  assign t[114] = (t[148] & t[149] & t[150] & ~t[151] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & ~t[151] & ~t[152] & t[153] & t[154]) | (~t[149] & ~t[150] & t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[150] & t[151] & ~t[153] & ~t[154]) | (~t[148] & ~t[149] & t[151] & ~t[152] & ~t[154]) | (~t[149] & t[150] & t[151] & t[152] & ~t[153]) | (~t[150] & t[151] & t[152] & ~t[154]);
  assign t[115] = (t[148] & t[149] & ~t[150] & ~t[152] & t[153] & ~t[154]) | (t[148] & t[150] & ~t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & t[152] & ~t[153] & ~t[154]) | (~t[148] & ~t[150] & ~t[151] & t[152] & ~t[153]) | (~t[148] & ~t[149] & ~t[151] & t[152] & ~t[154]) | (~t[148] & ~t[150] & t[151] & t[152] & t[153]) | (t[151] & t[152] & ~t[153] & ~t[154]);
  assign t[116] = (t[148] & t[149] & ~t[151] & t[152] & ~t[153] & ~t[154]) | (t[149] & ~t[150] & t[151] & ~t[152] & ~t[153] & t[154]) | (~t[149] & ~t[150] & ~t[151] & ~t[152] & t[153]) | (~t[148] & ~t[151] & ~t[152] & t[153] & ~t[154]) | (~t[148] & ~t[149] & ~t[150] & t[153] & ~t[154]) | (~t[149] & t[150] & ~t[151] & t[152] & t[153]) | (t[150] & ~t[152] & t[153] & ~t[154]);
  assign t[117] = (t[148] & t[149] & ~t[150] & t[151] & ~t[152] & ~t[154]) | (t[148] & ~t[150] & ~t[151] & t[152] & ~t[153] & t[154]) | (~t[149] & t[150] & ~t[151] & ~t[152] & ~t[154]) | (~t[148] & t[150] & ~t[151] & ~t[152] & ~t[153]) | (~t[148] & ~t[149] & t[150] & ~t[153] & ~t[154]) | (~t[148] & t[150] & t[151] & ~t[152] & t[153]) | (t[150] & ~t[151] & t[153] & ~t[154]);
  assign t[118] = (t[155] & ~t[157] & ~t[158] & ~t[159] & ~t[160]) | (t[155] & ~t[156] & ~t[158] & ~t[159] & ~t[161]) | (t[155] & ~t[156] & ~t[157] & ~t[160] & ~t[161]) | (~t[155] & t[156] & t[157] & t[158] & ~t[161]) | (~t[155] & t[156] & t[159] & t[160] & ~t[161]) | (t[155] & ~t[157] & ~t[159] & t[161]) | (~t[155] & t[157] & t[159] & t[161]);
  assign t[119] = (t[155] & t[156] & ~t[157] & ~t[159] & t[160] & ~t[161]) | (t[155] & t[157] & ~t[158] & ~t[159] & ~t[160] & t[161]) | (~t[156] & ~t[157] & t[159] & ~t[160] & ~t[161]) | (~t[155] & ~t[157] & ~t[158] & t[159] & ~t[160]) | (~t[155] & ~t[156] & ~t[158] & t[159] & ~t[161]) | (~t[155] & ~t[157] & t[158] & t[159] & t[160]) | (t[158] & t[159] & ~t[160] & ~t[161]);
  assign t[11] = t[52] ^ t[53];
  assign t[120] = t[162] ^ x[8];
  assign t[121] = t[163] ^ x[9];
  assign t[122] = t[164] ^ x[6];
  assign t[123] = t[165] ^ x[10];
  assign t[124] = t[166] ^ x[11];
  assign t[125] = t[167] ^ x[12];
  assign t[126] = t[168] ^ x[7];
  assign t[127] = t[169] ^ x[19];
  assign t[128] = t[170] ^ x[14];
  assign t[129] = t[171] ^ x[15];
  assign t[12] = t[16] & t[17];
  assign t[130] = t[172] ^ x[16];
  assign t[131] = t[173] ^ x[20];
  assign t[132] = t[174] ^ x[17];
  assign t[133] = t[175] ^ x[18];
  assign t[134] = t[176] ^ x[26];
  assign t[135] = t[177] ^ x[27];
  assign t[136] = t[178] ^ x[41];
  assign t[137] = t[179] ^ x[28];
  assign t[138] = t[180] ^ x[29];
  assign t[139] = t[181] ^ x[30];
  assign t[13] = t[54] ^ t[55];
  assign t[140] = t[182] ^ x[25];
  assign t[141] = t[183] ^ x[36];
  assign t[142] = t[184] ^ x[37];
  assign t[143] = t[185] ^ x[42];
  assign t[144] = t[186] ^ x[38];
  assign t[145] = t[187] ^ x[39];
  assign t[146] = t[188] ^ x[40];
  assign t[147] = t[189] ^ x[35];
  assign t[148] = t[190] ^ x[48];
  assign t[149] = t[191] ^ x[49];
  assign t[14] = t[18] & t[19];
  assign t[150] = t[192] ^ x[53];
  assign t[151] = t[193] ^ x[50];
  assign t[152] = t[194] ^ x[51];
  assign t[153] = t[195] ^ x[52];
  assign t[154] = t[196] ^ x[47];
  assign t[155] = t[197] ^ x[61];
  assign t[156] = t[198] ^ x[56];
  assign t[157] = t[199] ^ x[57];
  assign t[158] = t[200] ^ x[58];
  assign t[159] = t[201] ^ x[62];
  assign t[15] = ~(t[20]);
  assign t[160] = t[202] ^ x[59];
  assign t[161] = t[203] ^ x[60];
  assign t[162] = (x[2] & ~x[3] & ~x[4]) | (~x[2] & x[3] & ~x[4]) | (~x[2] & ~x[3] & x[4]) | (x[2] & x[3] & x[4]);
  assign t[163] = (x[2] & ~x[3] & ~x[5]) | (~x[2] & x[3] & ~x[5]) | (~x[2] & ~x[3] & x[5]) | (x[2] & x[3] & x[5]);
  assign t[164] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[165] = (x[2] & ~x[5]) | (~x[2] & x[5]);
  assign t[166] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[167] = (x[3] & ~x[5]) | (~x[3] & x[5]);
  assign t[168] = (x[4] & ~x[5]) | (~x[4] & x[5]);
  assign t[169] = (x[13] & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0);
  assign t[16] = ~(t[52]);
  assign t[170] = (x[13] & ~1'b0 & ~1'b0) | (~x[13] & 1'b0 & ~1'b0) | (~x[13] & ~1'b0 & 1'b0) | (x[13] & 1'b0 & 1'b0);
  assign t[171] = (x[13] & ~1'b0) | (~x[13] & 1'b0);
  assign t[172] = (x[13] & ~1'b0) | (~x[13] & 1'b0);
  assign t[173] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[174] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[175] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[176] = (x[21] & ~x[22] & ~x[23]) | (~x[21] & x[22] & ~x[23]) | (~x[21] & ~x[22] & x[23]) | (x[21] & x[22] & x[23]);
  assign t[177] = (x[21] & ~x[22] & ~x[24]) | (~x[21] & x[22] & ~x[24]) | (~x[21] & ~x[22] & x[24]) | (x[21] & x[22] & x[24]);
  assign t[178] = (x[21] & ~x[23]) | (~x[21] & x[23]);
  assign t[179] = (x[21] & ~x[24]) | (~x[21] & x[24]);
  assign t[17] = ~(t[56] ^ t[16]);
  assign t[180] = (x[22] & ~x[23]) | (~x[22] & x[23]);
  assign t[181] = (x[22] & ~x[24]) | (~x[22] & x[24]);
  assign t[182] = (x[23] & ~x[24]) | (~x[23] & x[24]);
  assign t[183] = (x[31] & ~x[32] & ~x[33]) | (~x[31] & x[32] & ~x[33]) | (~x[31] & ~x[32] & x[33]) | (x[31] & x[32] & x[33]);
  assign t[184] = (x[31] & ~x[32] & ~x[34]) | (~x[31] & x[32] & ~x[34]) | (~x[31] & ~x[32] & x[34]) | (x[31] & x[32] & x[34]);
  assign t[185] = (x[31] & ~x[33]) | (~x[31] & x[33]);
  assign t[186] = (x[31] & ~x[34]) | (~x[31] & x[34]);
  assign t[187] = (x[32] & ~x[33]) | (~x[32] & x[33]);
  assign t[188] = (x[32] & ~x[34]) | (~x[32] & x[34]);
  assign t[189] = (x[33] & ~x[34]) | (~x[33] & x[34]);
  assign t[18] = ~(t[54]);
  assign t[190] = (x[43] & ~x[44] & ~x[45]) | (~x[43] & x[44] & ~x[45]) | (~x[43] & ~x[44] & x[45]) | (x[43] & x[44] & x[45]);
  assign t[191] = (x[43] & ~x[44] & ~x[46]) | (~x[43] & x[44] & ~x[46]) | (~x[43] & ~x[44] & x[46]) | (x[43] & x[44] & x[46]);
  assign t[192] = (x[43] & ~x[45]) | (~x[43] & x[45]);
  assign t[193] = (x[43] & ~x[46]) | (~x[43] & x[46]);
  assign t[194] = (x[44] & ~x[45]) | (~x[44] & x[45]);
  assign t[195] = (x[44] & ~x[46]) | (~x[44] & x[46]);
  assign t[196] = (x[45] & ~x[46]) | (~x[45] & x[46]);
  assign t[197] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[198] = (x[55] & ~1'b0 & ~1'b0) | (~x[55] & 1'b0 & ~1'b0) | (~x[55] & ~1'b0 & 1'b0) | (x[55] & 1'b0 & 1'b0);
  assign t[199] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[19] = ~(t[57] ^ t[18]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[200] = (x[55] & ~1'b0) | (~x[55] & 1'b0);
  assign t[201] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[202] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[203] = (1'b0 & ~1'b0) | (~1'b0 & 1'b0);
  assign t[20] = t[21] ^ t[22];
  assign t[21] = t[58] ^ t[59];
  assign t[22] = t[23] & t[24];
  assign t[23] = ~(t[58]);
  assign t[24] = ~(t[60] ^ t[23]);
  assign t[25] = x[0] ? x[54] : t[26];
  assign t[26] = ~(t[27] ^ t[28]);
  assign t[27] = ~(t[29] ^ t[61]);
  assign t[28] = ~(t[30] ^ t[31]);
  assign t[29] = ~t[32];
  assign t[2] = ~(t[4] ^ t[50]);
  assign t[30] = ~(t[33]);
  assign t[31] = ~(t[34]);
  assign t[32] = ~(t[35] ^ t[62]);
  assign t[33] = t[36] ^ t[12];
  assign t[34] = t[37] ^ t[14];
  assign t[35] = ~t[38];
  assign t[36] = t[39] ^ t[40];
  assign t[37] = t[41] ^ t[42];
  assign t[38] = ~(t[43]);
  assign t[39] = t[63] ^ t[52];
  assign t[3] = ~(t[5] ^ t[6]);
  assign t[40] = t[16] & t[44];
  assign t[41] = t[64] ^ t[54];
  assign t[42] = t[18] & t[45];
  assign t[43] = t[46] ^ t[22];
  assign t[44] = t[56] ^ t[11];
  assign t[45] = t[57] ^ t[13];
  assign t[46] = t[47] ^ t[48];
  assign t[47] = t[65] ^ t[58];
  assign t[48] = t[23] & t[49];
  assign t[49] = t[60] ^ t[21];
  assign t[4] = ~t[7];
  assign t[50] = (t[66] & ~t[68] & ~t[70]) | (~t[67] & t[68] & ~t[69]) | (~t[66] & ~t[68] & t[70]) | (t[67] & t[68] & t[69]);
  assign t[51] = (t[71] & ~t[72]) | (~t[71] & t[72]);
  assign t[52] = (t[73] & ~t[75] & ~t[77]) | (~t[74] & t[75] & ~t[76]) | (~t[73] & ~t[75] & t[77]) | (t[74] & t[75] & t[76]);
  assign t[53] = (t[73] & ~t[75] & ~t[76]) | (~t[74] & t[75] & ~t[77]) | (~t[73] & ~t[75] & t[76]) | (t[74] & t[75] & t[77]);
  assign t[54] = (t[78] & ~t[80] & ~t[82]) | (~t[79] & t[80] & ~t[81]) | (~t[78] & ~t[80] & t[82]) | (t[79] & t[80] & t[81]);
  assign t[55] = (t[78] & ~t[80] & ~t[81]) | (~t[79] & t[80] & ~t[82]) | (~t[78] & ~t[80] & t[81]) | (t[79] & t[80] & t[82]);
  assign t[56] = (t[73] & ~t[83]) | (~t[73] & t[83]);
  assign t[57] = (t[78] & ~t[84]) | (~t[78] & t[84]);
  assign t[58] = (t[85] & ~t[87] & ~t[89]) | (~t[86] & t[87] & ~t[88]) | (~t[85] & ~t[87] & t[89]) | (t[86] & t[87] & t[88]);
  assign t[59] = (t[85] & ~t[87] & ~t[88]) | (~t[86] & t[87] & ~t[89]) | (~t[85] & ~t[87] & t[88]) | (t[86] & t[87] & t[89]);
  assign t[5] = ~(t[8]);
  assign t[60] = (t[85] & ~t[90]) | (~t[85] & t[90]);
  assign t[61] = (t[66] & ~t[68] & ~t[69]) | (~t[67] & t[68] & ~t[70]) | (~t[66] & ~t[68] & t[69]) | (t[67] & t[68] & t[70]);
  assign t[62] = (t[91] & ~t[92]) | (~t[91] & t[92]);
  assign t[63] = (t[73] & ~t[76]) | (~t[73] & t[76]);
  assign t[64] = (t[78] & ~t[81]) | (~t[78] & t[81]);
  assign t[65] = (t[85] & ~t[88]) | (~t[85] & t[88]);
  assign t[66] = t[93] ^ x[8];
  assign t[67] = t[94] ^ x[9];
  assign t[68] = t[95] ^ x[10];
  assign t[69] = t[96] ^ x[11];
  assign t[6] = ~(t[9]);
  assign t[70] = t[97] ^ x[12];
  assign t[71] = t[98] ^ x[19];
  assign t[72] = t[99] ^ x[20];
  assign t[73] = t[100] ^ x[26];
  assign t[74] = t[101] ^ x[27];
  assign t[75] = t[102] ^ x[28];
  assign t[76] = t[103] ^ x[29];
  assign t[77] = t[104] ^ x[30];
  assign t[78] = t[105] ^ x[36];
  assign t[79] = t[106] ^ x[37];
  assign t[7] = ~(t[10] ^ t[51]);
  assign t[80] = t[107] ^ x[38];
  assign t[81] = t[108] ^ x[39];
  assign t[82] = t[109] ^ x[40];
  assign t[83] = t[110] ^ x[41];
  assign t[84] = t[111] ^ x[42];
  assign t[85] = t[112] ^ x[48];
  assign t[86] = t[113] ^ x[49];
  assign t[87] = t[114] ^ x[50];
  assign t[88] = t[115] ^ x[51];
  assign t[89] = t[116] ^ x[52];
  assign t[8] = t[11] ^ t[12];
  assign t[90] = t[117] ^ x[53];
  assign t[91] = t[118] ^ x[61];
  assign t[92] = t[119] ^ x[62];
  assign t[93] = (t[120] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (t[120] & ~t[121] & ~t[123] & ~t[124] & ~t[126]) | (t[120] & ~t[121] & ~t[122] & ~t[125] & ~t[126]) | (~t[120] & t[121] & t[122] & t[123] & ~t[126]) | (~t[120] & t[121] & t[124] & t[125] & ~t[126]) | (t[120] & ~t[122] & ~t[124] & t[126]) | (~t[120] & t[122] & t[124] & t[126]);
  assign t[94] = (t[121] & ~t[122] & ~t[123] & ~t[124] & ~t[125]) | (~t[120] & t[121] & ~t[123] & ~t[124] & ~t[126]) | (~t[120] & t[121] & ~t[122] & ~t[125] & ~t[126]) | (t[120] & ~t[121] & t[122] & t[123] & ~t[126]) | (t[120] & ~t[121] & t[124] & t[125] & ~t[126]) | (t[121] & ~t[123] & ~t[125] & t[126]) | (~t[121] & t[123] & t[125] & t[126]);
  assign t[95] = (t[120] & t[121] & t[122] & ~t[123] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & ~t[123] & ~t[124] & t[125] & t[126]) | (~t[121] & ~t[122] & t[123] & ~t[124] & ~t[125]) | (~t[120] & ~t[122] & t[123] & ~t[125] & ~t[126]) | (~t[120] & ~t[121] & t[123] & ~t[124] & ~t[126]) | (~t[121] & t[122] & t[123] & t[124] & ~t[125]) | (~t[122] & t[123] & t[124] & ~t[126]);
  assign t[96] = (t[120] & t[121] & ~t[122] & ~t[124] & t[125] & ~t[126]) | (t[120] & t[122] & ~t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & t[124] & ~t[125] & ~t[126]) | (~t[120] & ~t[122] & ~t[123] & t[124] & ~t[125]) | (~t[120] & ~t[121] & ~t[123] & t[124] & ~t[126]) | (~t[120] & ~t[122] & t[123] & t[124] & t[125]) | (t[123] & t[124] & ~t[125] & ~t[126]);
  assign t[97] = (t[120] & t[121] & ~t[123] & t[124] & ~t[125] & ~t[126]) | (t[121] & ~t[122] & t[123] & ~t[124] & ~t[125] & t[126]) | (~t[121] & ~t[122] & ~t[123] & ~t[124] & t[125]) | (~t[120] & ~t[123] & ~t[124] & t[125] & ~t[126]) | (~t[120] & ~t[121] & ~t[122] & t[125] & ~t[126]) | (~t[121] & t[122] & ~t[123] & t[124] & t[125]) | (t[122] & ~t[124] & t[125] & ~t[126]);
  assign t[98] = (t[127] & ~t[129] & ~t[130] & ~t[131] & ~t[132]) | (t[127] & ~t[128] & ~t[130] & ~t[131] & ~t[133]) | (t[127] & ~t[128] & ~t[129] & ~t[132] & ~t[133]) | (~t[127] & t[128] & t[129] & t[130] & ~t[133]) | (~t[127] & t[128] & t[131] & t[132] & ~t[133]) | (t[127] & ~t[129] & ~t[131] & t[133]) | (~t[127] & t[129] & t[131] & t[133]);
  assign t[99] = (t[127] & t[128] & ~t[129] & ~t[131] & t[132] & ~t[133]) | (t[127] & t[129] & ~t[130] & ~t[131] & ~t[132] & t[133]) | (~t[128] & ~t[129] & t[131] & ~t[132] & ~t[133]) | (~t[127] & ~t[129] & ~t[130] & t[131] & ~t[132]) | (~t[127] & ~t[128] & ~t[130] & t[131] & ~t[133]) | (~t[127] & ~t[129] & t[130] & t[131] & t[132]) | (t[130] & t[131] & ~t[132] & ~t[133]);
  assign t[9] = t[13] ^ t[14];
  assign y = (t[0] & ~t[25]) | (~t[0] & t[25]);
endmodule

module R2ind168(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind169(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind170(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind171(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind172(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind173(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind174(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind175(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind176(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind177(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind178(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind179(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind180(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind181(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind182(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind183(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind184(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind185(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind186(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind187(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind188(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind189(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind190(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind191(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind192(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind193(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind194(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind195(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind196(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind197(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind198(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind199(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind200(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind201(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind202(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind203(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind204(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind205(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind206(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind207(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind208(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind209(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind210(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind211(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind212(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind213(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind214(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind215(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind216(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind217(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind218(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind219(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind220(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind221(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind222(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind223(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind224(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind225(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind226(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind227(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind228(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind229(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind230(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind231(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind232(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind233(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind234(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind235(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind236(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind237(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind238(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind239(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind240(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind241(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind242(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind243(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind244(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind245(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind246(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind247(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind248(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind249(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind250(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind251(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind252(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind253(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind254(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind255(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind256(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind257(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind258(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind259(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind260(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind261(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind262(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind263(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind264(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind265(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind266(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind267(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind268(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind269(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind270(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind271(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind272(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind273(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[11]) | (~t[9] & t[10] & ~t[7]) | (~t[6] & ~t[10] & t[11]) | (t[9] & t[10] & t[7]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind274(x, y);
 input [14:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = x[0] ? x[8] : t[3];
  assign t[10] = t[16] ^ x[12];
  assign t[11] = t[17] ^ x[13];
  assign t[12] = (t[18] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (t[18] & ~t[19] & ~t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[19] & ~t[20] & ~t[23] & ~t[24]) | (~t[18] & t[19] & t[20] & t[21] & ~t[24]) | (~t[18] & t[19] & t[22] & t[23] & ~t[24]) | (t[18] & ~t[20] & ~t[22] & t[24]) | (~t[18] & t[20] & t[22] & t[24]);
  assign t[13] = (t[18] & t[19] & ~t[20] & ~t[22] & t[23] & ~t[24]) | (t[18] & t[20] & ~t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & t[22] & ~t[23] & ~t[24]) | (~t[18] & ~t[20] & ~t[21] & t[22] & ~t[23]) | (~t[18] & ~t[19] & ~t[21] & t[22] & ~t[24]) | (~t[18] & ~t[20] & t[21] & t[22] & t[23]) | (t[21] & t[22] & ~t[23] & ~t[24]);
  assign t[14] = (t[18] & t[19] & ~t[20] & t[21] & ~t[22] & ~t[24]) | (t[18] & ~t[20] & ~t[21] & t[22] & ~t[23] & t[24]) | (~t[19] & t[20] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[19] & t[20] & ~t[23] & ~t[24]) | (~t[18] & t[20] & t[21] & ~t[22] & t[23]) | (t[20] & ~t[21] & t[23] & ~t[24]);
  assign t[15] = (t[19] & ~t[20] & ~t[21] & ~t[22] & ~t[23]) | (~t[18] & t[19] & ~t[21] & ~t[22] & ~t[24]) | (~t[18] & t[19] & ~t[20] & ~t[23] & ~t[24]) | (t[18] & ~t[19] & t[20] & t[21] & ~t[24]) | (t[18] & ~t[19] & t[22] & t[23] & ~t[24]) | (t[19] & ~t[21] & ~t[23] & t[24]) | (~t[19] & t[21] & t[23] & t[24]);
  assign t[16] = (t[18] & t[19] & t[20] & ~t[21] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & ~t[21] & ~t[22] & t[23] & t[24]) | (~t[19] & ~t[20] & t[21] & ~t[22] & ~t[23]) | (~t[18] & ~t[20] & t[21] & ~t[23] & ~t[24]) | (~t[18] & ~t[19] & t[21] & ~t[22] & ~t[24]) | (~t[19] & t[20] & t[21] & t[22] & ~t[23]) | (~t[20] & t[21] & t[22] & ~t[24]);
  assign t[17] = (t[18] & t[19] & ~t[21] & t[22] & ~t[23] & ~t[24]) | (t[19] & ~t[20] & t[21] & ~t[22] & ~t[23] & t[24]) | (~t[19] & ~t[20] & ~t[21] & ~t[22] & t[23]) | (~t[18] & ~t[21] & ~t[22] & t[23] & ~t[24]) | (~t[18] & ~t[19] & ~t[20] & t[23] & ~t[24]) | (~t[19] & t[20] & ~t[21] & t[22] & t[23]) | (t[20] & ~t[22] & t[23] & ~t[24]);
  assign t[18] = t[25] ^ x[6];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[10] : t[4];
  assign t[20] = t[27] ^ x[9];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[7];
  assign t[23] = t[30] ^ x[13];
  assign t[24] = t[31] ^ x[5];
  assign t[25] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[26] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[27] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[28] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[29] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[2] = x[0] ? x[14] : t[5];
  assign t[30] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[31] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[3] = (t[6] & ~t[7]) | (~t[6] & t[7]);
  assign t[4] = (t[6] & ~t[8]) | (~t[6] & t[8]);
  assign t[5] = (t[6] & ~t[10] & ~t[7]) | (~t[9] & t[10] & ~t[11]) | (~t[6] & ~t[10] & t[7]) | (t[9] & t[10] & t[11]);
  assign t[6] = t[12] ^ x[6];
  assign t[7] = t[13] ^ x[7];
  assign t[8] = t[14] ^ x[9];
  assign t[9] = t[15] ^ x[11];
  assign y = (t[0] & ~t[1] & ~t[2]) | (~t[0] & t[1] & ~t[2]) | (~t[0] & ~t[1] & t[2]) | (t[0] & t[1] & t[2]);
endmodule

module R2ind275(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[5]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[5]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind276(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[9] : t[2];
  assign t[10] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[11] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[12] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[10];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[11];
  assign t[18] = t[25] ^ x[8];
  assign t[19] = t[26] ^ x[12];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[5]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[5]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[10];
  assign t[7] = t[12] ^ x[11];
  assign t[8] = t[13] ^ x[12];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind277(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[9]) | (~t[6] & t[7] & ~t[8]) | (~t[4] & ~t[7] & t[9]) | (t[6] & t[7] & t[8]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind278(x, y);
 input [13:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = x[0] ? x[8] : t[2];
  assign t[10] = (t[16] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (t[16] & ~t[17] & ~t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[17] & ~t[18] & ~t[21] & ~t[22]) | (~t[16] & t[17] & t[18] & t[19] & ~t[22]) | (~t[16] & t[17] & t[20] & t[21] & ~t[22]) | (t[16] & ~t[18] & ~t[20] & t[22]) | (~t[16] & t[18] & t[20] & t[22]);
  assign t[11] = (t[16] & t[17] & ~t[18] & t[19] & ~t[20] & ~t[22]) | (t[16] & ~t[18] & ~t[19] & t[20] & ~t[21] & t[22]) | (~t[17] & t[18] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[17] & t[18] & ~t[21] & ~t[22]) | (~t[16] & t[18] & t[19] & ~t[20] & t[21]) | (t[18] & ~t[19] & t[21] & ~t[22]);
  assign t[12] = (t[17] & ~t[18] & ~t[19] & ~t[20] & ~t[21]) | (~t[16] & t[17] & ~t[19] & ~t[20] & ~t[22]) | (~t[16] & t[17] & ~t[18] & ~t[21] & ~t[22]) | (t[16] & ~t[17] & t[18] & t[19] & ~t[22]) | (t[16] & ~t[17] & t[20] & t[21] & ~t[22]) | (t[17] & ~t[19] & ~t[21] & t[22]) | (~t[17] & t[19] & t[21] & t[22]);
  assign t[13] = (t[16] & t[17] & t[18] & ~t[19] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & ~t[19] & ~t[20] & t[21] & t[22]) | (~t[17] & ~t[18] & t[19] & ~t[20] & ~t[21]) | (~t[16] & ~t[18] & t[19] & ~t[21] & ~t[22]) | (~t[16] & ~t[17] & t[19] & ~t[20] & ~t[22]) | (~t[17] & t[18] & t[19] & t[20] & ~t[21]) | (~t[18] & t[19] & t[20] & ~t[22]);
  assign t[14] = (t[16] & t[17] & ~t[18] & ~t[20] & t[21] & ~t[22]) | (t[16] & t[18] & ~t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & t[20] & ~t[21] & ~t[22]) | (~t[16] & ~t[18] & ~t[19] & t[20] & ~t[21]) | (~t[16] & ~t[17] & ~t[19] & t[20] & ~t[22]) | (~t[16] & ~t[18] & t[19] & t[20] & t[21]) | (t[19] & t[20] & ~t[21] & ~t[22]);
  assign t[15] = (t[16] & t[17] & ~t[19] & t[20] & ~t[21] & ~t[22]) | (t[17] & ~t[18] & t[19] & ~t[20] & ~t[21] & t[22]) | (~t[17] & ~t[18] & ~t[19] & ~t[20] & t[21]) | (~t[16] & ~t[19] & ~t[20] & t[21] & ~t[22]) | (~t[16] & ~t[17] & ~t[18] & t[21] & ~t[22]) | (~t[17] & t[18] & ~t[19] & t[20] & t[21]) | (t[18] & ~t[20] & t[21] & ~t[22]);
  assign t[16] = t[23] ^ x[6];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[7];
  assign t[19] = t[26] ^ x[10];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[11];
  assign t[21] = t[28] ^ x[12];
  assign t[22] = t[29] ^ x[5];
  assign t[23] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[24] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[25] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[26] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[27] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[28] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[29] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[5]) | (~t[4] & t[5]);
  assign t[3] = (t[4] & ~t[7] & ~t[8]) | (~t[6] & t[7] & ~t[9]) | (~t[4] & ~t[7] & t[8]) | (t[6] & t[7] & t[9]);
  assign t[4] = t[10] ^ x[6];
  assign t[5] = t[11] ^ x[7];
  assign t[6] = t[12] ^ x[9];
  assign t[7] = t[13] ^ x[10];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[12];
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2ind279(x, y);
 input [13:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = x[0] ? x[12] : t[2];
  assign t[10] = (t[15] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (~t[14] & t[15] & ~t[17] & ~t[18] & ~t[20]) | (~t[14] & t[15] & ~t[16] & ~t[19] & ~t[20]) | (t[14] & ~t[15] & t[16] & t[17] & ~t[20]) | (t[14] & ~t[15] & t[18] & t[19] & ~t[20]) | (t[15] & ~t[17] & ~t[19] & t[20]) | (~t[15] & t[17] & t[19] & t[20]);
  assign t[11] = (t[14] & t[15] & t[16] & ~t[17] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & ~t[17] & ~t[18] & t[19] & t[20]) | (~t[15] & ~t[16] & t[17] & ~t[18] & ~t[19]) | (~t[14] & ~t[16] & t[17] & ~t[19] & ~t[20]) | (~t[14] & ~t[15] & t[17] & ~t[18] & ~t[20]) | (~t[15] & t[16] & t[17] & t[18] & ~t[19]) | (~t[16] & t[17] & t[18] & ~t[20]);
  assign t[12] = (t[14] & t[15] & ~t[16] & ~t[18] & t[19] & ~t[20]) | (t[14] & t[16] & ~t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & t[18] & ~t[19] & ~t[20]) | (~t[14] & ~t[16] & ~t[17] & t[18] & ~t[19]) | (~t[14] & ~t[15] & ~t[17] & t[18] & ~t[20]) | (~t[14] & ~t[16] & t[17] & t[18] & t[19]) | (t[17] & t[18] & ~t[19] & ~t[20]);
  assign t[13] = (t[14] & t[15] & ~t[17] & t[18] & ~t[19] & ~t[20]) | (t[15] & ~t[16] & t[17] & ~t[18] & ~t[19] & t[20]) | (~t[15] & ~t[16] & ~t[17] & ~t[18] & t[19]) | (~t[14] & ~t[17] & ~t[18] & t[19] & ~t[20]) | (~t[14] & ~t[15] & ~t[16] & t[19] & ~t[20]) | (~t[15] & t[16] & ~t[17] & t[18] & t[19]) | (t[16] & ~t[18] & t[19] & ~t[20]);
  assign t[14] = t[21] ^ x[7];
  assign t[15] = t[22] ^ x[8];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[9];
  assign t[18] = t[25] ^ x[10];
  assign t[19] = t[26] ^ x[11];
  assign t[1] = x[0] ? x[13] : t[3];
  assign t[20] = t[27] ^ x[6];
  assign t[21] = (x[1] & ~x[2] & ~x[3]) | (~x[1] & x[2] & ~x[3]) | (~x[1] & ~x[2] & x[3]) | (x[1] & x[2] & x[3]);
  assign t[22] = (x[1] & ~x[2] & ~x[4]) | (~x[1] & x[2] & ~x[4]) | (~x[1] & ~x[2] & x[4]) | (x[1] & x[2] & x[4]);
  assign t[23] = (x[1] & ~x[3]) | (~x[1] & x[3]);
  assign t[24] = (x[1] & ~x[4]) | (~x[1] & x[4]);
  assign t[25] = (x[2] & ~x[3]) | (~x[2] & x[3]);
  assign t[26] = (x[2] & ~x[4]) | (~x[2] & x[4]);
  assign t[27] = (x[3] & ~x[4]) | (~x[3] & x[4]);
  assign t[2] = (t[4] & ~t[6] & ~t[8]) | (~t[5] & t[6] & ~t[7]) | (~t[4] & ~t[6] & t[8]) | (t[5] & t[6] & t[7]);
  assign t[3] = (t[4] & ~t[6] & ~t[7]) | (~t[5] & t[6] & ~t[8]) | (~t[4] & ~t[6] & t[7]) | (t[5] & t[6] & t[8]);
  assign t[4] = t[9] ^ x[7];
  assign t[5] = t[10] ^ x[8];
  assign t[6] = t[11] ^ x[9];
  assign t[7] = t[12] ^ x[10];
  assign t[8] = t[13] ^ x[11];
  assign t[9] = (t[14] & ~t[16] & ~t[17] & ~t[18] & ~t[19]) | (t[14] & ~t[15] & ~t[17] & ~t[18] & ~t[20]) | (t[14] & ~t[15] & ~t[16] & ~t[19] & ~t[20]) | (~t[14] & t[15] & t[16] & t[17] & ~t[20]) | (~t[14] & t[15] & t[18] & t[19] & ~t[20]) | (t[14] & ~t[16] & ~t[18] & t[20]) | (~t[14] & t[16] & t[18] & t[20]);
  assign y = (t[0] & ~t[1]) | (~t[0] & t[1]);
endmodule

module R2_ind(x, y);
 input [536:0] x;
 output [279:0] y;

  R2ind0 R2ind0_inst(.x({x[7], x[6], x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[6], x[5], x[4], x[3], x[2], x[7], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[6], x[5], x[4], x[3], x[1], x[7], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[6], x[5], x[4], x[2], x[1], x[7], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[6], x[5], x[3], x[2], x[1], x[7], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[5], x[6], x[4], x[3], x[2], x[1], x[7], x[0]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[6], x[5], x[4], x[3], x[2], x[1], x[7], x[0]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.y(y[19]));
  R2ind20 R2ind20_inst(.y(y[20]));
  R2ind21 R2ind21_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[56]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[56]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[56]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[56]}), .y(y[24]));
  R2ind25 R2ind25_inst(.y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[56]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[56]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[56]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[56]}), .y(y[31]));
  R2ind32 R2ind32_inst(.y(y[32]));
  R2ind33 R2ind33_inst(.y(y[33]));
  R2ind34 R2ind34_inst(.y(y[34]));
  R2ind35 R2ind35_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[56]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[56]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[56]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[56]}), .y(y[38]));
  R2ind39 R2ind39_inst(.y(y[39]));
  R2ind40 R2ind40_inst(.y(y[40]));
  R2ind41 R2ind41_inst(.y(y[41]));
  R2ind42 R2ind42_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[56]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[56]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[56]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[56]}), .y(y[45]));
  R2ind46 R2ind46_inst(.y(y[46]));
  R2ind47 R2ind47_inst(.y(y[47]));
  R2ind48 R2ind48_inst(.y(y[48]));
  R2ind49 R2ind49_inst(.x({x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[56]}), .y(y[52]));
  R2ind53 R2ind53_inst(.y(y[53]));
  R2ind54 R2ind54_inst(.y(y[54]));
  R2ind55 R2ind55_inst(.y(y[55]));
  R2ind56 R2ind56_inst(.x({x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[92], x[91], x[90], x[93], x[88], x[87], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[92], x[91], x[90], x[89], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[57], x[56]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[92], x[91], x[90], x[93], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[57], x[56]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[92], x[64], x[91], x[90], x[89], x[86], x[84], x[83], x[85], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[73], x[72], x[74], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[87], x[56]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[92], x[64], x[91], x[90], x[93], x[86], x[84], x[83], x[85], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[73], x[72], x[74], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[87], x[56]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[93], x[82], x[86], x[85], x[84], x[83], x[81], x[80], x[79], x[78], x[77], x[76], x[71], x[75], x[74], x[73], x[72], x[70], x[69], x[68], x[67], x[66], x[65], x[92], x[64], x[91], x[90], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[89], x[56]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[56]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[129], x[128], x[127], x[130], x[125], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[56]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[129], x[128], x[127], x[126], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[94], x[56]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[129], x[128], x[127], x[130], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[94], x[56]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[129], x[101], x[128], x[127], x[126], x[123], x[121], x[120], x[122], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[110], x[109], x[111], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[124], x[56]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[129], x[101], x[128], x[127], x[130], x[123], x[121], x[120], x[122], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[110], x[109], x[111], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[124], x[56]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[130], x[119], x[123], x[122], x[121], x[120], x[118], x[117], x[116], x[115], x[114], x[113], x[108], x[112], x[111], x[110], x[109], x[107], x[106], x[105], x[104], x[103], x[102], x[129], x[101], x[128], x[127], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[126], x[56]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[56]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[166], x[165], x[164], x[167], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[56]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[166], x[165], x[164], x[163], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[131], x[56]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[166], x[165], x[164], x[167], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[131], x[56]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[166], x[138], x[165], x[164], x[163], x[160], x[158], x[157], x[159], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[147], x[146], x[148], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[161], x[56]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[166], x[138], x[165], x[164], x[167], x[160], x[158], x[157], x[159], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[147], x[146], x[148], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[161], x[56]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[167], x[156], x[160], x[159], x[158], x[157], x[155], x[154], x[153], x[152], x[151], x[150], x[145], x[149], x[148], x[147], x[146], x[144], x[143], x[142], x[141], x[140], x[139], x[166], x[138], x[165], x[164], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[163], x[56]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[202], x[201], x[200], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[56]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[202], x[201], x[204], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[168], x[56]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[202], x[201], x[200], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[168], x[56]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[202], x[201], x[204], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[183], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[168], x[56]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[175], x[202], x[201], x[200], x[197], x[195], x[194], x[196], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[184], x[183], x[185], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[198], x[56]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[175], x[202], x[201], x[204], x[197], x[195], x[194], x[196], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[186], x[184], x[183], x[185], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[198], x[56]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[204], x[193], x[197], x[196], x[195], x[194], x[192], x[191], x[190], x[189], x[188], x[187], x[182], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[203], x[175], x[202], x[201], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[200], x[56]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[56]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[229], x[228], x[227], x[230], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[56]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[229], x[228], x[227], x[226], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[212], x[211], x[210], x[225], x[209], x[208], x[207], x[206], x[205], x[56]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[229], x[228], x[227], x[230], x[223], x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[212], x[211], x[210], x[225], x[209], x[208], x[207], x[206], x[205], x[56]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[229], x[212], x[228], x[227], x[226], x[223], x[221], x[220], x[222], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[75], x[73], x[72], x[74], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[225], x[211], x[210], x[209], x[208], x[207], x[206], x[224], x[56]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[229], x[212], x[228], x[227], x[230], x[223], x[221], x[220], x[222], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[75], x[73], x[72], x[74], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[225], x[211], x[210], x[209], x[208], x[207], x[206], x[224], x[56]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[230], x[219], x[223], x[222], x[221], x[220], x[218], x[217], x[216], x[215], x[214], x[213], x[71], x[75], x[74], x[73], x[72], x[70], x[69], x[68], x[67], x[66], x[65], x[229], x[212], x[228], x[227], x[211], x[210], x[225], x[209], x[208], x[207], x[206], x[226], x[56]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[56]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[255], x[254], x[253], x[256], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[56]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[255], x[254], x[253], x[252], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[238], x[237], x[236], x[251], x[235], x[234], x[233], x[232], x[231], x[56]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[255], x[254], x[253], x[256], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[238], x[237], x[236], x[251], x[235], x[234], x[233], x[232], x[231], x[56]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[255], x[238], x[254], x[253], x[252], x[249], x[247], x[246], x[248], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[112], x[110], x[109], x[111], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[251], x[237], x[236], x[235], x[234], x[233], x[232], x[250], x[56]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[255], x[238], x[254], x[253], x[256], x[249], x[247], x[246], x[248], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[112], x[110], x[109], x[111], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[251], x[237], x[236], x[235], x[234], x[233], x[232], x[250], x[56]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[256], x[245], x[249], x[248], x[247], x[246], x[244], x[243], x[242], x[241], x[240], x[239], x[108], x[112], x[111], x[110], x[109], x[107], x[106], x[105], x[104], x[103], x[102], x[255], x[238], x[254], x[253], x[237], x[236], x[251], x[235], x[234], x[233], x[232], x[252], x[56]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[281], x[280], x[279], x[278], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[277], x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[149], x[148], x[147], x[146], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[56]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[281], x[280], x[279], x[282], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[277], x[276], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[149], x[148], x[147], x[146], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257], x[56]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[281], x[280], x[279], x[278], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[149], x[148], x[147], x[146], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[264], x[263], x[262], x[277], x[261], x[260], x[259], x[258], x[257], x[56]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[281], x[280], x[279], x[282], x[275], x[274], x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[149], x[148], x[147], x[146], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[264], x[263], x[262], x[277], x[261], x[260], x[259], x[258], x[257], x[56]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[281], x[264], x[280], x[279], x[278], x[275], x[273], x[272], x[274], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[149], x[147], x[146], x[148], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[277], x[263], x[262], x[261], x[260], x[259], x[258], x[276], x[56]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[281], x[264], x[280], x[279], x[282], x[275], x[273], x[272], x[274], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[149], x[147], x[146], x[148], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[277], x[263], x[262], x[261], x[260], x[259], x[258], x[276], x[56]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[282], x[271], x[275], x[274], x[273], x[272], x[270], x[269], x[268], x[267], x[266], x[265], x[145], x[149], x[148], x[147], x[146], x[144], x[143], x[142], x[141], x[140], x[139], x[281], x[264], x[280], x[279], x[263], x[262], x[277], x[261], x[260], x[259], x[258], x[278], x[56]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[307], x[306], x[305], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[56]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[307], x[306], x[305], x[308], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[56]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[307], x[306], x[305], x[304], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[290], x[289], x[288], x[303], x[287], x[286], x[285], x[284], x[283], x[56]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[307], x[306], x[305], x[308], x[301], x[300], x[299], x[298], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[290], x[289], x[288], x[303], x[287], x[286], x[285], x[284], x[283], x[56]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[307], x[290], x[306], x[305], x[304], x[301], x[299], x[298], x[300], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[186], x[184], x[183], x[185], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[303], x[289], x[288], x[287], x[286], x[285], x[284], x[302], x[56]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[307], x[290], x[306], x[305], x[308], x[301], x[299], x[298], x[300], x[297], x[296], x[295], x[294], x[293], x[292], x[291], x[186], x[184], x[183], x[185], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[303], x[289], x[288], x[287], x[286], x[285], x[284], x[302], x[56]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[308], x[297], x[301], x[300], x[299], x[298], x[296], x[295], x[294], x[293], x[292], x[291], x[182], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[307], x[290], x[306], x[305], x[289], x[288], x[303], x[287], x[286], x[285], x[284], x[304], x[56]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[92], x[91], x[90], x[311], x[88], x[310], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[309], x[56]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[92], x[91], x[90], x[312], x[88], x[310], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[309], x[56]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[92], x[91], x[90], x[311], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[309], x[56]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[92], x[91], x[90], x[312], x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[309], x[56]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[92], x[64], x[91], x[90], x[311], x[86], x[84], x[83], x[85], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[310], x[56]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[92], x[64], x[91], x[90], x[312], x[86], x[84], x[83], x[85], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[310], x[56]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[312], x[82], x[86], x[85], x[84], x[83], x[81], x[80], x[79], x[78], x[77], x[76], x[92], x[64], x[91], x[90], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[311], x[56]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[129], x[128], x[127], x[315], x[125], x[314], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[313], x[56]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[129], x[128], x[127], x[316], x[125], x[314], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[313], x[56]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[129], x[128], x[127], x[315], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[313], x[56]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[129], x[128], x[127], x[316], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[313], x[56]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[129], x[101], x[128], x[127], x[315], x[123], x[121], x[120], x[122], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[314], x[56]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[129], x[101], x[128], x[127], x[316], x[123], x[121], x[120], x[122], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[314], x[56]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[316], x[119], x[123], x[122], x[121], x[120], x[118], x[117], x[116], x[115], x[114], x[113], x[129], x[101], x[128], x[127], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[315], x[56]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[166], x[165], x[164], x[319], x[162], x[318], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[317], x[56]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[166], x[165], x[164], x[320], x[162], x[318], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[317], x[56]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[166], x[165], x[164], x[319], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[317], x[56]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[166], x[165], x[164], x[320], x[160], x[159], x[158], x[157], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[317], x[56]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[166], x[138], x[165], x[164], x[319], x[160], x[158], x[157], x[159], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[318], x[56]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[166], x[138], x[165], x[164], x[320], x[160], x[158], x[157], x[159], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[318], x[56]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[320], x[156], x[160], x[159], x[158], x[157], x[155], x[154], x[153], x[152], x[151], x[150], x[166], x[138], x[165], x[164], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[319], x[56]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[202], x[201], x[323], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[322], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[321], x[56]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[202], x[201], x[324], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[322], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[321], x[56]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[202], x[201], x[323], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[321], x[56]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[202], x[201], x[324], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[321], x[56]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[175], x[202], x[201], x[323], x[197], x[195], x[194], x[196], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[322], x[56]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[175], x[202], x[201], x[324], x[197], x[195], x[194], x[196], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[322], x[56]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[324], x[193], x[197], x[196], x[195], x[194], x[192], x[191], x[190], x[189], x[188], x[187], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[175], x[202], x[201], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[323], x[56]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[92], x[91], x[90], x[338], x[88], x[337], x[86], x[85], x[84], x[83], x[336], x[335], x[334], x[333], x[75], x[74], x[73], x[72], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[325], x[56]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[92], x[91], x[90], x[339], x[88], x[337], x[86], x[85], x[84], x[83], x[336], x[335], x[334], x[333], x[75], x[74], x[73], x[72], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[325], x[56]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[92], x[91], x[90], x[338], x[86], x[85], x[84], x[83], x[336], x[335], x[334], x[333], x[75], x[74], x[73], x[72], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[325], x[56]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[92], x[91], x[90], x[339], x[86], x[85], x[84], x[83], x[336], x[335], x[334], x[333], x[75], x[74], x[73], x[72], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[325], x[56]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[92], x[64], x[91], x[90], x[338], x[86], x[84], x[83], x[85], x[336], x[334], x[333], x[335], x[75], x[73], x[72], x[74], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[337], x[56]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[92], x[64], x[91], x[90], x[339], x[86], x[84], x[83], x[85], x[336], x[334], x[333], x[335], x[75], x[73], x[72], x[74], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[337], x[56]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[339], x[82], x[332], x[71], x[86], x[85], x[84], x[83], x[81], x[80], x[79], x[78], x[77], x[76], x[336], x[335], x[334], x[333], x[331], x[330], x[329], x[328], x[327], x[326], x[75], x[74], x[73], x[72], x[70], x[69], x[68], x[67], x[66], x[65], x[92], x[64], x[91], x[90], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[338], x[56]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[129], x[128], x[127], x[353], x[125], x[352], x[123], x[122], x[121], x[120], x[351], x[350], x[349], x[348], x[112], x[111], x[110], x[109], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[340], x[56]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[129], x[128], x[127], x[354], x[125], x[352], x[123], x[122], x[121], x[120], x[351], x[350], x[349], x[348], x[112], x[111], x[110], x[109], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[340], x[56]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[129], x[128], x[127], x[353], x[123], x[122], x[121], x[120], x[351], x[350], x[349], x[348], x[112], x[111], x[110], x[109], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[340], x[56]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[129], x[128], x[127], x[354], x[123], x[122], x[121], x[120], x[351], x[350], x[349], x[348], x[112], x[111], x[110], x[109], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[340], x[56]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[129], x[101], x[128], x[127], x[353], x[112], x[110], x[109], x[111], x[123], x[121], x[120], x[122], x[351], x[349], x[348], x[350], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[352], x[56]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[129], x[101], x[128], x[127], x[354], x[112], x[110], x[109], x[111], x[123], x[121], x[120], x[122], x[351], x[349], x[348], x[350], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[347], x[346], x[345], x[344], x[343], x[342], x[341], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[352], x[56]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[354], x[119], x[347], x[108], x[123], x[122], x[121], x[120], x[118], x[117], x[116], x[115], x[114], x[113], x[351], x[350], x[349], x[348], x[346], x[345], x[344], x[343], x[342], x[341], x[112], x[111], x[110], x[109], x[107], x[106], x[105], x[104], x[103], x[102], x[129], x[101], x[128], x[127], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[353], x[56]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[166], x[165], x[164], x[368], x[162], x[367], x[160], x[159], x[158], x[157], x[366], x[365], x[364], x[363], x[149], x[148], x[147], x[146], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[355], x[56]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[166], x[165], x[164], x[369], x[162], x[367], x[160], x[159], x[158], x[157], x[366], x[365], x[364], x[363], x[149], x[148], x[147], x[146], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[355], x[56]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[166], x[165], x[164], x[368], x[160], x[159], x[158], x[157], x[366], x[365], x[364], x[363], x[149], x[148], x[147], x[146], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[355], x[56]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[166], x[165], x[164], x[369], x[160], x[159], x[158], x[157], x[366], x[365], x[364], x[363], x[149], x[148], x[147], x[146], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[355], x[56]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[166], x[138], x[165], x[164], x[368], x[160], x[158], x[157], x[159], x[366], x[364], x[363], x[365], x[149], x[147], x[146], x[148], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[367], x[56]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[166], x[138], x[165], x[164], x[369], x[160], x[158], x[157], x[159], x[366], x[364], x[363], x[365], x[149], x[147], x[146], x[148], x[156], x[155], x[154], x[153], x[152], x[151], x[150], x[362], x[361], x[360], x[359], x[358], x[357], x[356], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[367], x[56]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[369], x[156], x[362], x[145], x[160], x[159], x[158], x[157], x[155], x[154], x[153], x[152], x[151], x[150], x[366], x[365], x[364], x[363], x[361], x[360], x[359], x[358], x[357], x[356], x[149], x[148], x[147], x[146], x[144], x[143], x[142], x[141], x[140], x[139], x[166], x[138], x[165], x[164], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[368], x[56]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[202], x[201], x[383], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[382], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[381], x[380], x[379], x[378], x[186], x[185], x[184], x[183], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[370], x[56]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[202], x[201], x[384], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[382], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[381], x[380], x[379], x[378], x[186], x[185], x[184], x[183], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[370], x[56]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[202], x[201], x[383], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[381], x[380], x[379], x[378], x[186], x[185], x[184], x[183], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[370], x[56]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[202], x[201], x[384], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[381], x[380], x[379], x[378], x[186], x[185], x[184], x[183], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[55], x[54], x[53], x[52], x[51], x[50], x[49], x[48], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[370], x[56]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[175], x[202], x[201], x[383], x[197], x[195], x[194], x[196], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[381], x[379], x[378], x[380], x[186], x[184], x[183], x[185], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[382], x[56]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[203], x[175], x[202], x[201], x[384], x[197], x[195], x[194], x[196], x[193], x[192], x[191], x[190], x[189], x[188], x[187], x[381], x[379], x[378], x[380], x[186], x[184], x[183], x[185], x[377], x[376], x[375], x[374], x[373], x[372], x[371], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[382], x[56]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[384], x[193], x[197], x[196], x[195], x[194], x[192], x[191], x[190], x[189], x[188], x[187], x[377], x[182], x[381], x[380], x[379], x[378], x[376], x[375], x[374], x[373], x[372], x[371], x[186], x[185], x[184], x[183], x[181], x[180], x[179], x[178], x[177], x[176], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[203], x[175], x[202], x[201], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[383], x[56]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[387], x[307], x[306], x[305], x[386], x[303], x[385], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[56]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[388], x[307], x[306], x[305], x[386], x[303], x[385], x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[56]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[387], x[307], x[306], x[305], x[385], x[290], x[289], x[288], x[303], x[287], x[286], x[285], x[284], x[56]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[388], x[307], x[306], x[305], x[385], x[290], x[289], x[288], x[303], x[287], x[286], x[285], x[284], x[56]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[387], x[307], x[290], x[306], x[305], x[386], x[303], x[289], x[288], x[287], x[286], x[285], x[284], x[56]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[388], x[307], x[290], x[306], x[305], x[386], x[303], x[289], x[288], x[287], x[286], x[285], x[284], x[56]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[388], x[387], x[307], x[290], x[306], x[305], x[289], x[288], x[303], x[287], x[286], x[285], x[284], x[56]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[391], x[229], x[228], x[227], x[390], x[225], x[389], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[56]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[392], x[229], x[228], x[227], x[390], x[225], x[389], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[56]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[391], x[229], x[228], x[227], x[389], x[212], x[211], x[210], x[225], x[209], x[208], x[207], x[206], x[56]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[392], x[229], x[228], x[227], x[389], x[212], x[211], x[210], x[225], x[209], x[208], x[207], x[206], x[56]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[391], x[229], x[212], x[228], x[227], x[390], x[225], x[211], x[210], x[209], x[208], x[207], x[206], x[56]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[392], x[229], x[212], x[228], x[227], x[390], x[225], x[211], x[210], x[209], x[208], x[207], x[206], x[56]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[392], x[391], x[229], x[212], x[228], x[227], x[211], x[210], x[225], x[209], x[208], x[207], x[206], x[56]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[395], x[255], x[254], x[253], x[394], x[251], x[393], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[56]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[396], x[255], x[254], x[253], x[394], x[251], x[393], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[56]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[395], x[255], x[254], x[253], x[393], x[238], x[237], x[236], x[251], x[235], x[234], x[233], x[232], x[56]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[396], x[255], x[254], x[253], x[393], x[238], x[237], x[236], x[251], x[235], x[234], x[233], x[232], x[56]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[395], x[255], x[238], x[254], x[253], x[394], x[251], x[237], x[236], x[235], x[234], x[233], x[232], x[56]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[396], x[255], x[238], x[254], x[253], x[394], x[251], x[237], x[236], x[235], x[234], x[233], x[232], x[56]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[396], x[395], x[255], x[238], x[254], x[253], x[237], x[236], x[251], x[235], x[234], x[233], x[232], x[56]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[399], x[281], x[280], x[279], x[398], x[277], x[397], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[56]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[400], x[281], x[280], x[279], x[398], x[277], x[397], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[56]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[399], x[281], x[280], x[279], x[397], x[264], x[263], x[262], x[277], x[261], x[260], x[259], x[258], x[56]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[400], x[281], x[280], x[279], x[397], x[264], x[263], x[262], x[277], x[261], x[260], x[259], x[258], x[56]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[399], x[281], x[264], x[280], x[279], x[398], x[277], x[263], x[262], x[261], x[260], x[259], x[258], x[56]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[400], x[281], x[264], x[280], x[279], x[398], x[277], x[263], x[262], x[261], x[260], x[259], x[258], x[56]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[400], x[399], x[281], x[264], x[280], x[279], x[263], x[262], x[277], x[261], x[260], x[259], x[258], x[56]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[403], x[92], x[91], x[90], x[402], x[88], x[401], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[56]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[404], x[92], x[91], x[90], x[402], x[88], x[401], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[56]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[403], x[92], x[91], x[90], x[401], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[56]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[404], x[92], x[91], x[90], x[401], x[64], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[56]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[403], x[92], x[64], x[91], x[90], x[402], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[56]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[404], x[92], x[64], x[91], x[90], x[402], x[88], x[63], x[62], x[61], x[60], x[59], x[58], x[56]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[404], x[403], x[92], x[64], x[91], x[90], x[63], x[62], x[88], x[61], x[60], x[59], x[58], x[56]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[407], x[129], x[128], x[127], x[406], x[125], x[405], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[56]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[408], x[129], x[128], x[127], x[406], x[125], x[405], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[56]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[407], x[129], x[128], x[127], x[405], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[56]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[408], x[129], x[128], x[127], x[405], x[101], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[56]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[407], x[129], x[101], x[128], x[127], x[406], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[56]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[408], x[129], x[101], x[128], x[127], x[406], x[125], x[100], x[99], x[98], x[97], x[96], x[95], x[56]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[408], x[407], x[129], x[101], x[128], x[127], x[100], x[99], x[125], x[98], x[97], x[96], x[95], x[56]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[411], x[166], x[165], x[164], x[410], x[162], x[409], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[56]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[412], x[166], x[165], x[164], x[410], x[162], x[409], x[138], x[137], x[136], x[135], x[134], x[133], x[132], x[56]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[411], x[166], x[165], x[164], x[409], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[56]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[412], x[166], x[165], x[164], x[409], x[138], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[56]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[411], x[166], x[138], x[165], x[164], x[410], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[56]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[412], x[166], x[138], x[165], x[164], x[410], x[162], x[137], x[136], x[135], x[134], x[133], x[132], x[56]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[412], x[411], x[166], x[138], x[165], x[164], x[137], x[136], x[162], x[135], x[134], x[133], x[132], x[56]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[415], x[203], x[202], x[201], x[414], x[199], x[413], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[56]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[416], x[203], x[202], x[201], x[414], x[199], x[413], x[175], x[174], x[173], x[172], x[171], x[170], x[169], x[56]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[415], x[203], x[202], x[201], x[413], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[56]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[416], x[203], x[202], x[201], x[413], x[175], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[56]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[415], x[203], x[175], x[202], x[201], x[414], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[56]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[416], x[203], x[175], x[202], x[201], x[414], x[199], x[174], x[173], x[172], x[171], x[170], x[169], x[56]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[416], x[415], x[203], x[175], x[202], x[201], x[174], x[173], x[199], x[172], x[171], x[170], x[169], x[56]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418], x[417], x[56]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[431], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[418], x[417], x[56]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[430], x[429], x[428], x[427], x[424], x[423], x[422], x[421], x[425], x[420], x[419], x[418], x[417], x[56]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[431], x[429], x[428], x[427], x[424], x[423], x[422], x[421], x[425], x[420], x[419], x[418], x[417], x[56]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[430], x[429], x[423], x[428], x[427], x[426], x[425], x[422], x[421], x[420], x[419], x[418], x[417], x[56]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[431], x[429], x[423], x[428], x[427], x[426], x[425], x[422], x[421], x[420], x[419], x[418], x[417], x[56]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[431], x[430], x[429], x[423], x[428], x[427], x[422], x[421], x[425], x[420], x[419], x[418], x[417], x[56]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[56]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[446], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[56]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[445], x[444], x[443], x[442], x[439], x[438], x[437], x[436], x[440], x[435], x[434], x[433], x[432], x[56]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[446], x[444], x[443], x[442], x[439], x[438], x[437], x[436], x[440], x[435], x[434], x[433], x[432], x[56]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[445], x[444], x[438], x[443], x[442], x[441], x[440], x[437], x[436], x[435], x[434], x[433], x[432], x[56]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[446], x[444], x[438], x[443], x[442], x[441], x[440], x[437], x[436], x[435], x[434], x[433], x[432], x[56]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[446], x[445], x[444], x[438], x[443], x[442], x[437], x[436], x[440], x[435], x[434], x[433], x[432], x[56]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[460], x[459], x[458], x[457], x[456], x[455], x[454], x[453], x[452], x[451], x[450], x[449], x[448], x[447], x[56]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[461], x[459], x[458], x[457], x[456], x[455], x[454], x[453], x[452], x[451], x[450], x[449], x[448], x[447], x[56]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[460], x[459], x[458], x[457], x[454], x[453], x[452], x[451], x[455], x[450], x[449], x[448], x[447], x[56]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[461], x[459], x[458], x[457], x[454], x[453], x[452], x[451], x[455], x[450], x[449], x[448], x[447], x[56]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[460], x[459], x[453], x[458], x[457], x[456], x[455], x[452], x[451], x[450], x[449], x[448], x[447], x[56]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[461], x[459], x[453], x[458], x[457], x[456], x[455], x[452], x[451], x[450], x[449], x[448], x[447], x[56]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[461], x[460], x[459], x[453], x[458], x[457], x[452], x[451], x[455], x[450], x[449], x[448], x[447], x[56]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[467], x[466], x[465], x[464], x[463], x[462], x[56]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[476], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[467], x[466], x[465], x[464], x[463], x[462], x[56]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[475], x[474], x[473], x[472], x[469], x[468], x[467], x[466], x[470], x[465], x[464], x[463], x[462], x[56]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[476], x[474], x[473], x[472], x[469], x[468], x[467], x[466], x[470], x[465], x[464], x[463], x[462], x[56]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[475], x[474], x[468], x[473], x[472], x[471], x[470], x[467], x[466], x[465], x[464], x[463], x[462], x[56]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[476], x[474], x[468], x[473], x[472], x[471], x[470], x[467], x[466], x[465], x[464], x[463], x[462], x[56]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[476], x[475], x[474], x[468], x[473], x[472], x[467], x[466], x[470], x[465], x[464], x[463], x[462], x[56]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[490], x[489], x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[56]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[491], x[489], x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479], x[478], x[477], x[56]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[490], x[489], x[488], x[487], x[484], x[483], x[482], x[481], x[485], x[480], x[479], x[478], x[477], x[56]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[491], x[489], x[488], x[487], x[484], x[483], x[482], x[481], x[485], x[480], x[479], x[478], x[477], x[56]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[490], x[489], x[483], x[488], x[487], x[486], x[485], x[482], x[481], x[480], x[479], x[478], x[477], x[56]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[491], x[489], x[483], x[488], x[487], x[486], x[485], x[482], x[481], x[480], x[479], x[478], x[477], x[56]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[491], x[490], x[489], x[483], x[488], x[487], x[482], x[481], x[485], x[480], x[479], x[478], x[477], x[56]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[505], x[504], x[503], x[502], x[501], x[500], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[56]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[506], x[504], x[503], x[502], x[501], x[500], x[499], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[56]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[505], x[504], x[503], x[502], x[499], x[498], x[497], x[496], x[500], x[495], x[494], x[493], x[492], x[56]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[506], x[504], x[503], x[502], x[499], x[498], x[497], x[496], x[500], x[495], x[494], x[493], x[492], x[56]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[505], x[504], x[498], x[503], x[502], x[501], x[500], x[497], x[496], x[495], x[494], x[493], x[492], x[56]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[506], x[504], x[498], x[503], x[502], x[501], x[500], x[497], x[496], x[495], x[494], x[493], x[492], x[56]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[506], x[505], x[504], x[498], x[503], x[502], x[497], x[496], x[500], x[495], x[494], x[493], x[492], x[56]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[520], x[519], x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[511], x[510], x[509], x[508], x[507], x[56]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[521], x[519], x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[511], x[510], x[509], x[508], x[507], x[56]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[520], x[519], x[518], x[517], x[514], x[513], x[512], x[511], x[515], x[510], x[509], x[508], x[507], x[56]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[521], x[519], x[518], x[517], x[514], x[513], x[512], x[511], x[515], x[510], x[509], x[508], x[507], x[56]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[520], x[519], x[513], x[518], x[517], x[516], x[515], x[512], x[511], x[510], x[509], x[508], x[507], x[56]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[521], x[519], x[513], x[518], x[517], x[516], x[515], x[512], x[511], x[510], x[509], x[508], x[507], x[56]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[521], x[520], x[519], x[513], x[518], x[517], x[512], x[511], x[515], x[510], x[509], x[508], x[507], x[56]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[535], x[534], x[533], x[532], x[531], x[530], x[529], x[528], x[527], x[526], x[525], x[524], x[523], x[522], x[56]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[536], x[534], x[533], x[532], x[531], x[530], x[529], x[528], x[527], x[526], x[525], x[524], x[523], x[522], x[56]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[535], x[534], x[533], x[532], x[529], x[528], x[527], x[526], x[530], x[525], x[524], x[523], x[522], x[56]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[536], x[534], x[533], x[532], x[529], x[528], x[527], x[526], x[530], x[525], x[524], x[523], x[522], x[56]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[535], x[534], x[528], x[533], x[532], x[531], x[530], x[527], x[526], x[525], x[524], x[523], x[522], x[56]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[536], x[534], x[528], x[533], x[532], x[531], x[530], x[527], x[526], x[525], x[524], x[523], x[522], x[56]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[536], x[535], x[534], x[528], x[533], x[532], x[527], x[526], x[530], x[525], x[524], x[523], x[522], x[56]}), .y(y[279]));
endmodule

