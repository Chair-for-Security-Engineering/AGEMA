/* modified netlist. Source: module CRAFT in file Designs/CRAFT_round-based/AGEMA/CRAFT.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module CRAFT_HPC2_BDDcudd_Pipeline_d1 (plaintext_s0, key_s0, clk, rst, key_s1, plaintext_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [63:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input rst ;
    input [127:0] key_s1 ;
    input [63:0] plaintext_s1 ;
    input [228:0] Fresh ;
    output [63:0] ciphertext_s0 ;
    output done ;
    output [63:0] ciphertext_s1 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_275 ;
    wire signal_276 ;
    wire signal_277 ;
    wire signal_278 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_281 ;
    wire signal_282 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_285 ;
    wire signal_286 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_291 ;
    wire signal_292 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_295 ;
    wire signal_296 ;
    wire signal_297 ;
    wire signal_298 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_305 ;
    wire signal_306 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1185 ;
    wire signal_1187 ;
    wire signal_1189 ;
    wire signal_1191 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1196 ;
    wire signal_1198 ;
    wire signal_1200 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1205 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1223 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1228 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1238 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1244 ;
    wire signal_1247 ;
    wire signal_1250 ;
    wire signal_1253 ;
    wire signal_1256 ;
    wire signal_1259 ;
    wire signal_1262 ;
    wire signal_1265 ;
    wire signal_1268 ;
    wire signal_1271 ;
    wire signal_1274 ;
    wire signal_1277 ;
    wire signal_1280 ;
    wire signal_1283 ;
    wire signal_1286 ;
    wire signal_1289 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1294 ;
    wire signal_1296 ;
    wire signal_1298 ;
    wire signal_1300 ;
    wire signal_1302 ;
    wire signal_1304 ;
    wire signal_1306 ;
    wire signal_1308 ;
    wire signal_1310 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1404 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1427 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1451 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1492 ;
    wire signal_1494 ;
    wire signal_1496 ;
    wire signal_1498 ;
    wire signal_1500 ;
    wire signal_1502 ;
    wire signal_1504 ;
    wire signal_1506 ;
    wire signal_1508 ;
    wire signal_1510 ;
    wire signal_1512 ;
    wire signal_1514 ;
    wire signal_1516 ;
    wire signal_1518 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1524 ;
    wire signal_1526 ;
    wire signal_1528 ;
    wire signal_1530 ;
    wire signal_1532 ;
    wire signal_1534 ;
    wire signal_1536 ;
    wire signal_1538 ;
    wire signal_1540 ;
    wire signal_1542 ;
    wire signal_1544 ;
    wire signal_1546 ;
    wire signal_1548 ;
    wire signal_1550 ;
    wire signal_1552 ;
    wire signal_1554 ;
    wire signal_1556 ;
    wire signal_1559 ;
    wire signal_1562 ;
    wire signal_1565 ;
    wire signal_1568 ;
    wire signal_1571 ;
    wire signal_1574 ;
    wire signal_1577 ;
    wire signal_1580 ;
    wire signal_1583 ;
    wire signal_1586 ;
    wire signal_1589 ;
    wire signal_1592 ;
    wire signal_1595 ;
    wire signal_1598 ;
    wire signal_1601 ;
    wire signal_1604 ;
    wire signal_1607 ;
    wire signal_1610 ;
    wire signal_1613 ;
    wire signal_1616 ;
    wire signal_1619 ;
    wire signal_1622 ;
    wire signal_1625 ;
    wire signal_1628 ;
    wire signal_1631 ;
    wire signal_1634 ;
    wire signal_1637 ;
    wire signal_1640 ;
    wire signal_1643 ;
    wire signal_1646 ;
    wire signal_1649 ;
    wire signal_1652 ;
    wire signal_1655 ;
    wire signal_1658 ;
    wire signal_1661 ;
    wire signal_1664 ;
    wire signal_1667 ;
    wire signal_1670 ;
    wire signal_1673 ;
    wire signal_1676 ;
    wire signal_1679 ;
    wire signal_1682 ;
    wire signal_1685 ;
    wire signal_1688 ;
    wire signal_1691 ;
    wire signal_1694 ;
    wire signal_1697 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1734 ;
    wire signal_1736 ;
    wire signal_1738 ;
    wire signal_1740 ;
    wire signal_1742 ;
    wire signal_1744 ;
    wire signal_1746 ;
    wire signal_1748 ;
    wire signal_1750 ;
    wire signal_1752 ;
    wire signal_1754 ;
    wire signal_1756 ;
    wire signal_1758 ;
    wire signal_1760 ;
    wire signal_1762 ;
    wire signal_1764 ;
    wire signal_1766 ;
    wire signal_1768 ;
    wire signal_1770 ;
    wire signal_1772 ;
    wire signal_1774 ;
    wire signal_1776 ;
    wire signal_1778 ;
    wire signal_1780 ;
    wire signal_1782 ;
    wire signal_1784 ;
    wire signal_1786 ;
    wire signal_1788 ;
    wire signal_1790 ;
    wire signal_1792 ;
    wire signal_1794 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2392 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2395 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2398 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2401 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2404 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_3858 ;
    wire signal_3859 ;
    wire signal_3860 ;
    wire signal_3861 ;
    wire signal_3862 ;
    wire signal_3863 ;
    wire signal_3864 ;
    wire signal_3865 ;
    wire signal_3866 ;
    wire signal_3867 ;
    wire signal_3868 ;
    wire signal_3869 ;
    wire signal_3870 ;
    wire signal_3871 ;
    wire signal_3872 ;
    wire signal_3873 ;
    wire signal_3874 ;
    wire signal_3875 ;
    wire signal_3876 ;
    wire signal_3877 ;
    wire signal_3878 ;
    wire signal_3879 ;
    wire signal_3880 ;
    wire signal_3881 ;
    wire signal_3882 ;
    wire signal_3883 ;
    wire signal_3884 ;
    wire signal_3885 ;
    wire signal_3886 ;
    wire signal_3887 ;
    wire signal_3888 ;
    wire signal_3889 ;
    wire signal_3890 ;
    wire signal_3891 ;
    wire signal_3892 ;
    wire signal_3893 ;
    wire signal_3894 ;
    wire signal_3895 ;
    wire signal_3896 ;
    wire signal_3897 ;
    wire signal_3898 ;
    wire signal_3899 ;
    wire signal_3900 ;
    wire signal_3901 ;
    wire signal_3902 ;
    wire signal_3903 ;
    wire signal_3904 ;
    wire signal_3905 ;
    wire signal_3906 ;
    wire signal_3907 ;
    wire signal_3908 ;
    wire signal_3909 ;
    wire signal_3910 ;
    wire signal_3911 ;
    wire signal_3912 ;
    wire signal_3913 ;
    wire signal_3914 ;
    wire signal_3915 ;
    wire signal_3916 ;
    wire signal_3917 ;
    wire signal_3918 ;
    wire signal_3919 ;
    wire signal_3920 ;
    wire signal_3921 ;
    wire signal_3922 ;
    wire signal_3923 ;
    wire signal_3924 ;
    wire signal_3925 ;
    wire signal_3926 ;
    wire signal_3927 ;
    wire signal_3928 ;
    wire signal_3929 ;
    wire signal_3930 ;
    wire signal_3931 ;
    wire signal_3932 ;
    wire signal_3933 ;
    wire signal_3934 ;
    wire signal_3935 ;
    wire signal_3936 ;
    wire signal_3937 ;
    wire signal_3938 ;
    wire signal_3939 ;
    wire signal_3940 ;
    wire signal_3941 ;
    wire signal_3942 ;
    wire signal_3943 ;
    wire signal_3944 ;
    wire signal_3945 ;
    wire signal_3946 ;
    wire signal_3947 ;
    wire signal_3948 ;
    wire signal_3949 ;
    wire signal_3950 ;
    wire signal_3951 ;
    wire signal_3952 ;
    wire signal_3953 ;
    wire signal_3954 ;
    wire signal_3955 ;
    wire signal_3956 ;
    wire signal_3957 ;
    wire signal_3958 ;
    wire signal_3959 ;
    wire signal_3960 ;
    wire signal_3961 ;
    wire signal_3962 ;
    wire signal_3963 ;
    wire signal_3964 ;
    wire signal_3965 ;
    wire signal_3966 ;
    wire signal_3967 ;
    wire signal_3968 ;
    wire signal_3969 ;
    wire signal_3970 ;
    wire signal_3971 ;
    wire signal_3972 ;
    wire signal_3973 ;
    wire signal_3974 ;
    wire signal_3975 ;
    wire signal_3976 ;
    wire signal_3977 ;
    wire signal_3978 ;
    wire signal_3979 ;
    wire signal_3980 ;
    wire signal_3981 ;
    wire signal_3982 ;
    wire signal_3983 ;
    wire signal_3984 ;
    wire signal_3985 ;
    wire signal_3986 ;
    wire signal_3987 ;
    wire signal_3988 ;
    wire signal_3989 ;
    wire signal_3990 ;
    wire signal_3991 ;
    wire signal_3992 ;
    wire signal_3993 ;
    wire signal_3994 ;
    wire signal_3995 ;
    wire signal_3996 ;
    wire signal_3997 ;
    wire signal_3998 ;
    wire signal_3999 ;
    wire signal_4000 ;
    wire signal_4001 ;
    wire signal_4002 ;
    wire signal_4003 ;
    wire signal_4004 ;
    wire signal_4005 ;
    wire signal_4006 ;
    wire signal_4007 ;
    wire signal_4008 ;
    wire signal_4009 ;
    wire signal_4010 ;
    wire signal_4011 ;
    wire signal_4012 ;
    wire signal_4013 ;
    wire signal_4014 ;
    wire signal_4015 ;
    wire signal_4016 ;
    wire signal_4017 ;
    wire signal_4018 ;
    wire signal_4019 ;
    wire signal_4020 ;
    wire signal_4021 ;
    wire signal_4022 ;
    wire signal_4023 ;
    wire signal_4024 ;
    wire signal_4025 ;
    wire signal_4026 ;
    wire signal_4027 ;
    wire signal_4028 ;
    wire signal_4029 ;
    wire signal_4030 ;
    wire signal_4031 ;
    wire signal_4032 ;
    wire signal_4033 ;
    wire signal_4034 ;
    wire signal_4035 ;
    wire signal_4036 ;
    wire signal_4037 ;
    wire signal_4038 ;
    wire signal_4039 ;
    wire signal_4040 ;
    wire signal_4041 ;
    wire signal_4042 ;
    wire signal_4043 ;
    wire signal_4044 ;
    wire signal_4045 ;
    wire signal_4046 ;
    wire signal_4047 ;
    wire signal_4048 ;
    wire signal_4049 ;
    wire signal_4050 ;
    wire signal_4051 ;
    wire signal_4052 ;
    wire signal_4053 ;
    wire signal_4054 ;
    wire signal_4055 ;
    wire signal_4056 ;
    wire signal_4057 ;
    wire signal_4058 ;
    wire signal_4059 ;
    wire signal_4060 ;
    wire signal_4061 ;
    wire signal_4062 ;
    wire signal_4063 ;
    wire signal_4064 ;
    wire signal_4065 ;
    wire signal_4066 ;
    wire signal_4067 ;
    wire signal_4068 ;
    wire signal_4069 ;
    wire signal_4070 ;
    wire signal_4071 ;
    wire signal_4072 ;
    wire signal_4073 ;
    wire signal_4074 ;
    wire signal_4075 ;
    wire signal_4076 ;
    wire signal_4077 ;
    wire signal_4078 ;
    wire signal_4079 ;
    wire signal_4080 ;
    wire signal_4081 ;
    wire signal_4082 ;
    wire signal_4083 ;
    wire signal_4084 ;
    wire signal_4085 ;
    wire signal_4086 ;
    wire signal_4087 ;
    wire signal_4088 ;
    wire signal_4089 ;
    wire signal_4090 ;
    wire signal_4091 ;
    wire signal_4092 ;
    wire signal_4093 ;
    wire signal_4094 ;
    wire signal_4095 ;
    wire signal_4096 ;
    wire signal_4097 ;
    wire signal_4098 ;
    wire signal_4099 ;
    wire signal_4100 ;
    wire signal_4101 ;
    wire signal_4102 ;
    wire signal_4103 ;
    wire signal_4104 ;
    wire signal_4105 ;
    wire signal_4106 ;
    wire signal_4107 ;
    wire signal_4108 ;
    wire signal_4109 ;
    wire signal_4110 ;
    wire signal_4111 ;
    wire signal_4112 ;
    wire signal_4113 ;
    wire signal_4114 ;
    wire signal_4115 ;
    wire signal_4116 ;
    wire signal_4117 ;
    wire signal_4118 ;
    wire signal_4119 ;
    wire signal_4120 ;
    wire signal_4121 ;
    wire signal_4122 ;
    wire signal_4123 ;
    wire signal_4124 ;
    wire signal_4125 ;
    wire signal_4126 ;
    wire signal_4127 ;
    wire signal_4128 ;
    wire signal_4129 ;
    wire signal_4130 ;
    wire signal_4131 ;
    wire signal_4132 ;
    wire signal_4133 ;
    wire signal_4134 ;
    wire signal_4135 ;
    wire signal_4136 ;
    wire signal_4137 ;
    wire signal_4138 ;
    wire signal_4139 ;
    wire signal_4140 ;
    wire signal_4141 ;
    wire signal_4142 ;
    wire signal_4143 ;
    wire signal_4144 ;
    wire signal_4145 ;
    wire signal_4146 ;
    wire signal_4147 ;
    wire signal_4148 ;
    wire signal_4149 ;
    wire signal_4150 ;
    wire signal_4151 ;
    wire signal_4152 ;
    wire signal_4153 ;
    wire signal_4154 ;
    wire signal_4155 ;
    wire signal_4156 ;
    wire signal_4157 ;
    wire signal_4158 ;
    wire signal_4159 ;
    wire signal_4160 ;
    wire signal_4161 ;
    wire signal_4162 ;
    wire signal_4163 ;
    wire signal_4164 ;
    wire signal_4165 ;
    wire signal_4166 ;
    wire signal_4167 ;
    wire signal_4168 ;
    wire signal_4169 ;
    wire signal_4170 ;
    wire signal_4171 ;
    wire signal_4172 ;
    wire signal_4173 ;
    wire signal_4174 ;
    wire signal_4175 ;
    wire signal_4176 ;
    wire signal_4177 ;
    wire signal_4178 ;
    wire signal_4179 ;
    wire signal_4180 ;
    wire signal_4181 ;
    wire signal_4182 ;
    wire signal_4183 ;
    wire signal_4184 ;
    wire signal_4185 ;
    wire signal_4186 ;
    wire signal_4187 ;
    wire signal_4188 ;
    wire signal_4189 ;
    wire signal_4190 ;
    wire signal_4191 ;
    wire signal_4192 ;
    wire signal_4193 ;
    wire signal_4194 ;
    wire signal_4195 ;
    wire signal_4196 ;
    wire signal_4197 ;
    wire signal_4198 ;
    wire signal_4199 ;
    wire signal_4200 ;
    wire signal_4201 ;
    wire signal_4202 ;
    wire signal_4203 ;
    wire signal_4204 ;
    wire signal_4205 ;
    wire signal_4206 ;
    wire signal_4207 ;
    wire signal_4208 ;
    wire signal_4209 ;
    wire signal_4210 ;
    wire signal_4211 ;
    wire signal_4212 ;
    wire signal_4213 ;
    wire signal_4214 ;
    wire signal_4215 ;
    wire signal_4216 ;
    wire signal_4217 ;
    wire signal_4218 ;
    wire signal_4219 ;
    wire signal_4220 ;
    wire signal_4221 ;
    wire signal_4222 ;
    wire signal_4223 ;
    wire signal_4224 ;
    wire signal_4225 ;
    wire signal_4226 ;
    wire signal_4227 ;
    wire signal_4228 ;
    wire signal_4229 ;
    wire signal_4230 ;
    wire signal_4231 ;
    wire signal_4232 ;
    wire signal_4233 ;
    wire signal_4234 ;
    wire signal_4235 ;
    wire signal_4236 ;
    wire signal_4237 ;
    wire signal_4238 ;
    wire signal_4239 ;
    wire signal_4240 ;
    wire signal_4241 ;
    wire signal_4242 ;
    wire signal_4243 ;
    wire signal_4244 ;
    wire signal_4245 ;
    wire signal_4246 ;
    wire signal_4247 ;
    wire signal_4248 ;
    wire signal_4249 ;
    wire signal_4250 ;
    wire signal_4251 ;
    wire signal_4252 ;
    wire signal_4253 ;
    wire signal_4254 ;
    wire signal_4255 ;
    wire signal_4256 ;
    wire signal_4257 ;
    wire signal_4258 ;
    wire signal_4259 ;
    wire signal_4260 ;
    wire signal_4261 ;
    wire signal_4262 ;
    wire signal_4263 ;
    wire signal_4264 ;
    wire signal_4265 ;
    wire signal_4266 ;
    wire signal_4267 ;
    wire signal_4268 ;
    wire signal_4269 ;
    wire signal_4270 ;
    wire signal_4271 ;
    wire signal_4272 ;
    wire signal_4273 ;
    wire signal_4274 ;
    wire signal_4275 ;
    wire signal_4276 ;
    wire signal_4277 ;
    wire signal_4278 ;
    wire signal_4279 ;
    wire signal_4280 ;
    wire signal_4281 ;
    wire signal_4282 ;
    wire signal_4283 ;
    wire signal_4284 ;
    wire signal_4285 ;
    wire signal_4286 ;
    wire signal_4287 ;
    wire signal_4288 ;
    wire signal_4289 ;
    wire signal_4290 ;
    wire signal_4291 ;
    wire signal_4292 ;
    wire signal_4293 ;
    wire signal_4294 ;
    wire signal_4295 ;
    wire signal_4296 ;
    wire signal_4297 ;
    wire signal_4298 ;
    wire signal_4299 ;
    wire signal_4300 ;
    wire signal_4301 ;
    wire signal_4302 ;
    wire signal_4303 ;
    wire signal_4304 ;
    wire signal_4305 ;
    wire signal_4306 ;
    wire signal_4307 ;
    wire signal_4308 ;
    wire signal_4309 ;
    wire signal_4310 ;
    wire signal_4311 ;
    wire signal_4312 ;
    wire signal_4313 ;
    wire signal_4314 ;
    wire signal_4315 ;
    wire signal_4316 ;
    wire signal_4317 ;
    wire signal_4318 ;
    wire signal_4319 ;
    wire signal_4320 ;
    wire signal_4321 ;
    wire signal_4322 ;
    wire signal_4323 ;
    wire signal_4324 ;
    wire signal_4325 ;
    wire signal_4326 ;
    wire signal_4327 ;
    wire signal_4328 ;
    wire signal_4329 ;
    wire signal_4330 ;
    wire signal_4331 ;
    wire signal_4332 ;
    wire signal_4333 ;
    wire signal_4334 ;
    wire signal_4335 ;
    wire signal_4336 ;
    wire signal_4337 ;
    wire signal_4338 ;
    wire signal_4339 ;
    wire signal_4340 ;
    wire signal_4341 ;
    wire signal_4342 ;
    wire signal_4343 ;
    wire signal_4344 ;
    wire signal_4345 ;
    wire signal_4346 ;
    wire signal_4347 ;
    wire signal_4348 ;
    wire signal_4349 ;
    wire signal_4350 ;
    wire signal_4351 ;
    wire signal_4352 ;
    wire signal_4353 ;
    wire signal_4354 ;
    wire signal_4355 ;
    wire signal_4356 ;
    wire signal_4357 ;
    wire signal_4358 ;
    wire signal_4359 ;
    wire signal_4360 ;
    wire signal_4361 ;
    wire signal_4362 ;
    wire signal_4363 ;
    wire signal_4364 ;
    wire signal_4365 ;
    wire signal_4366 ;
    wire signal_4367 ;
    wire signal_4368 ;
    wire signal_4369 ;
    wire signal_4370 ;
    wire signal_4371 ;
    wire signal_4372 ;
    wire signal_4373 ;
    wire signal_4374 ;
    wire signal_4375 ;
    wire signal_4376 ;
    wire signal_4377 ;
    wire signal_4378 ;
    wire signal_4379 ;
    wire signal_4380 ;
    wire signal_4381 ;
    wire signal_4382 ;
    wire signal_4383 ;
    wire signal_4384 ;
    wire signal_4385 ;
    wire signal_4386 ;
    wire signal_4387 ;
    wire signal_4388 ;
    wire signal_4389 ;
    wire signal_4390 ;
    wire signal_4391 ;
    wire signal_4392 ;
    wire signal_4393 ;
    wire signal_4394 ;
    wire signal_4395 ;
    wire signal_4396 ;
    wire signal_4397 ;
    wire signal_4398 ;
    wire signal_4399 ;
    wire signal_4400 ;
    wire signal_4401 ;
    wire signal_4402 ;
    wire signal_4403 ;
    wire signal_4404 ;
    wire signal_4405 ;
    wire signal_4406 ;
    wire signal_4407 ;
    wire signal_4408 ;
    wire signal_4409 ;
    wire signal_4410 ;
    wire signal_4411 ;
    wire signal_4412 ;
    wire signal_4413 ;
    wire signal_4414 ;
    wire signal_4415 ;
    wire signal_4416 ;
    wire signal_4417 ;
    wire signal_4418 ;
    wire signal_4419 ;
    wire signal_4420 ;
    wire signal_4421 ;
    wire signal_4422 ;
    wire signal_4423 ;
    wire signal_4424 ;
    wire signal_4425 ;
    wire signal_4426 ;
    wire signal_4427 ;
    wire signal_4428 ;
    wire signal_4429 ;
    wire signal_4430 ;
    wire signal_4431 ;
    wire signal_4432 ;
    wire signal_4433 ;
    wire signal_4434 ;
    wire signal_4435 ;
    wire signal_4436 ;
    wire signal_4437 ;
    wire signal_4438 ;
    wire signal_4439 ;
    wire signal_4440 ;
    wire signal_4441 ;
    wire signal_4442 ;
    wire signal_4443 ;
    wire signal_4444 ;
    wire signal_4445 ;
    wire signal_4446 ;
    wire signal_4447 ;
    wire signal_4448 ;
    wire signal_4449 ;
    wire signal_4450 ;
    wire signal_4451 ;
    wire signal_4452 ;
    wire signal_4453 ;
    wire signal_4454 ;
    wire signal_4455 ;
    wire signal_4456 ;
    wire signal_4457 ;
    wire signal_4458 ;
    wire signal_4459 ;
    wire signal_4460 ;
    wire signal_4461 ;
    wire signal_4462 ;
    wire signal_4463 ;
    wire signal_4464 ;
    wire signal_4465 ;
    wire signal_4466 ;
    wire signal_4467 ;
    wire signal_4468 ;
    wire signal_4469 ;
    wire signal_4470 ;
    wire signal_4471 ;
    wire signal_4472 ;
    wire signal_4473 ;
    wire signal_4474 ;
    wire signal_4475 ;
    wire signal_4476 ;
    wire signal_4477 ;
    wire signal_4478 ;
    wire signal_4479 ;
    wire signal_4480 ;
    wire signal_4481 ;
    wire signal_4482 ;
    wire signal_4483 ;
    wire signal_4484 ;
    wire signal_4485 ;
    wire signal_4486 ;
    wire signal_4487 ;
    wire signal_4488 ;
    wire signal_4489 ;
    wire signal_4490 ;
    wire signal_4491 ;
    wire signal_4492 ;
    wire signal_4493 ;
    wire signal_4494 ;
    wire signal_4495 ;
    wire signal_4496 ;
    wire signal_4497 ;
    wire signal_4498 ;
    wire signal_4499 ;
    wire signal_4500 ;
    wire signal_4501 ;
    wire signal_4502 ;
    wire signal_4503 ;
    wire signal_4504 ;
    wire signal_4505 ;
    wire signal_4506 ;
    wire signal_4507 ;
    wire signal_4508 ;
    wire signal_4509 ;
    wire signal_4510 ;
    wire signal_4511 ;
    wire signal_4512 ;
    wire signal_4513 ;
    wire signal_4514 ;
    wire signal_4515 ;
    wire signal_4516 ;
    wire signal_4517 ;
    wire signal_4518 ;
    wire signal_4519 ;
    wire signal_4520 ;
    wire signal_4521 ;
    wire signal_4522 ;
    wire signal_4523 ;
    wire signal_4524 ;
    wire signal_4525 ;
    wire signal_4526 ;
    wire signal_4527 ;
    wire signal_4528 ;
    wire signal_4529 ;
    wire signal_4530 ;
    wire signal_4531 ;
    wire signal_4532 ;
    wire signal_4533 ;
    wire signal_4534 ;
    wire signal_4535 ;
    wire signal_4536 ;
    wire signal_4537 ;
    wire signal_4538 ;
    wire signal_4539 ;
    wire signal_4540 ;
    wire signal_4541 ;
    wire signal_4542 ;
    wire signal_4543 ;
    wire signal_4544 ;
    wire signal_4545 ;
    wire signal_4546 ;
    wire signal_4547 ;
    wire signal_4548 ;
    wire signal_4549 ;
    wire signal_4550 ;
    wire signal_4551 ;
    wire signal_4552 ;
    wire signal_4553 ;
    wire signal_4554 ;
    wire signal_4555 ;
    wire signal_4556 ;
    wire signal_4557 ;
    wire signal_4558 ;
    wire signal_4559 ;
    wire signal_4560 ;
    wire signal_4561 ;
    wire signal_4562 ;
    wire signal_4563 ;
    wire signal_4564 ;
    wire signal_4565 ;
    wire signal_4566 ;
    wire signal_4567 ;
    wire signal_4568 ;
    wire signal_4569 ;
    wire signal_4570 ;
    wire signal_4571 ;
    wire signal_4572 ;
    wire signal_4573 ;
    wire signal_4574 ;
    wire signal_4575 ;
    wire signal_4576 ;
    wire signal_4577 ;
    wire signal_4578 ;
    wire signal_4579 ;
    wire signal_4580 ;
    wire signal_4581 ;
    wire signal_4582 ;
    wire signal_4583 ;
    wire signal_4584 ;
    wire signal_4585 ;
    wire signal_4586 ;
    wire signal_4587 ;
    wire signal_4588 ;
    wire signal_4589 ;
    wire signal_4590 ;
    wire signal_4591 ;
    wire signal_4592 ;
    wire signal_4593 ;
    wire signal_4594 ;
    wire signal_4595 ;
    wire signal_4596 ;
    wire signal_4597 ;
    wire signal_4598 ;
    wire signal_4599 ;
    wire signal_4600 ;
    wire signal_4601 ;
    wire signal_4602 ;
    wire signal_4603 ;
    wire signal_4604 ;
    wire signal_4605 ;
    wire signal_4606 ;
    wire signal_4607 ;
    wire signal_4608 ;
    wire signal_4609 ;
    wire signal_4610 ;
    wire signal_4611 ;
    wire signal_4612 ;
    wire signal_4613 ;
    wire signal_4614 ;
    wire signal_4615 ;
    wire signal_4616 ;
    wire signal_4617 ;
    wire signal_4618 ;
    wire signal_4619 ;
    wire signal_4620 ;
    wire signal_4621 ;
    wire signal_4622 ;
    wire signal_4623 ;
    wire signal_4624 ;
    wire signal_4625 ;
    wire signal_4626 ;
    wire signal_4627 ;
    wire signal_4628 ;
    wire signal_4629 ;
    wire signal_4630 ;
    wire signal_4631 ;
    wire signal_4632 ;
    wire signal_4633 ;
    wire signal_4634 ;
    wire signal_4635 ;
    wire signal_4636 ;
    wire signal_4637 ;
    wire signal_4638 ;
    wire signal_4639 ;
    wire signal_4640 ;
    wire signal_4641 ;
    wire signal_4642 ;
    wire signal_4643 ;
    wire signal_4644 ;
    wire signal_4645 ;
    wire signal_4646 ;
    wire signal_4647 ;
    wire signal_4648 ;
    wire signal_4649 ;
    wire signal_4650 ;
    wire signal_4651 ;
    wire signal_4652 ;
    wire signal_4653 ;
    wire signal_4654 ;
    wire signal_4655 ;
    wire signal_4656 ;
    wire signal_4657 ;
    wire signal_4658 ;
    wire signal_4659 ;
    wire signal_4660 ;
    wire signal_4661 ;
    wire signal_4662 ;
    wire signal_4663 ;
    wire signal_4664 ;
    wire signal_4665 ;
    wire signal_4666 ;
    wire signal_4667 ;
    wire signal_4668 ;
    wire signal_4669 ;
    wire signal_4670 ;
    wire signal_4671 ;
    wire signal_4672 ;
    wire signal_4673 ;
    wire signal_4674 ;
    wire signal_4675 ;
    wire signal_4676 ;
    wire signal_4677 ;
    wire signal_4678 ;
    wire signal_4679 ;
    wire signal_4680 ;
    wire signal_4681 ;
    wire signal_4682 ;
    wire signal_4683 ;
    wire signal_4684 ;
    wire signal_4685 ;
    wire signal_4686 ;
    wire signal_4687 ;
    wire signal_4688 ;
    wire signal_4689 ;
    wire signal_4690 ;
    wire signal_4691 ;
    wire signal_4692 ;
    wire signal_4693 ;
    wire signal_4694 ;
    wire signal_4695 ;
    wire signal_4696 ;
    wire signal_4697 ;
    wire signal_4698 ;
    wire signal_4699 ;
    wire signal_4700 ;
    wire signal_4701 ;
    wire signal_4702 ;
    wire signal_4703 ;
    wire signal_4704 ;
    wire signal_4705 ;
    wire signal_4706 ;
    wire signal_4707 ;
    wire signal_4708 ;
    wire signal_4709 ;
    wire signal_4710 ;
    wire signal_4711 ;
    wire signal_4712 ;
    wire signal_4713 ;
    wire signal_4714 ;
    wire signal_4715 ;
    wire signal_4716 ;
    wire signal_4717 ;
    wire signal_4718 ;
    wire signal_4719 ;
    wire signal_4720 ;
    wire signal_4721 ;
    wire signal_4722 ;
    wire signal_4723 ;
    wire signal_4724 ;
    wire signal_4725 ;
    wire signal_4726 ;
    wire signal_4727 ;
    wire signal_4728 ;
    wire signal_4729 ;
    wire signal_4730 ;
    wire signal_4731 ;
    wire signal_4732 ;
    wire signal_4733 ;
    wire signal_4734 ;
    wire signal_4735 ;
    wire signal_4736 ;
    wire signal_4737 ;
    wire signal_4738 ;
    wire signal_4739 ;
    wire signal_4740 ;
    wire signal_4741 ;
    wire signal_4742 ;
    wire signal_4743 ;
    wire signal_4744 ;
    wire signal_4745 ;
    wire signal_4746 ;
    wire signal_4747 ;
    wire signal_4748 ;
    wire signal_4749 ;
    wire signal_4750 ;
    wire signal_4751 ;
    wire signal_4752 ;
    wire signal_4753 ;
    wire signal_4754 ;
    wire signal_4755 ;
    wire signal_4756 ;
    wire signal_4757 ;
    wire signal_4758 ;
    wire signal_4759 ;
    wire signal_4760 ;
    wire signal_4761 ;

    /* cells in depth 0 */
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_177 ( .a ({signal_1646, signal_894}), .b ({1'b0, signal_266}), .c ({signal_1821, signal_333}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_180 ( .a ({signal_1649, signal_893}), .b ({1'b0, signal_1014}), .c ({signal_1822, signal_335}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_183 ( .a ({signal_1652, signal_892}), .b ({1'b0, signal_1013}), .c ({signal_1823, signal_337}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_186 ( .a ({signal_1655, signal_891}), .b ({1'b0, 1'b0}), .c ({signal_1824, signal_339}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_189 ( .a ({signal_1658, signal_890}), .b ({1'b0, signal_265}), .c ({signal_1825, signal_341}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_192 ( .a ({signal_1661, signal_889}), .b ({1'b0, signal_1011}), .c ({signal_1826, signal_343}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_195 ( .a ({signal_1664, signal_888}), .b ({1'b0, signal_1010}), .c ({signal_1827, signal_345}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_198 ( .a ({signal_1667, signal_887}), .b ({1'b0, signal_1009}), .c ({signal_1828, signal_347}) ) ;
    INV_X1 cell_712 ( .A (signal_1000), .ZN (signal_692) ) ;
    INV_X1 cell_713 ( .A (signal_692), .ZN (signal_693) ) ;
    INV_X1 cell_714 ( .A (signal_692), .ZN (signal_694) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_715 ( .s (signal_1000), .b ({key_s1[64], key_s0[64]}), .a ({key_s1[0], key_s0[0]}), .c ({signal_1244, signal_934}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_716 ( .s (signal_693), .b ({key_s1[65], key_s0[65]}), .a ({key_s1[1], key_s0[1]}), .c ({signal_1559, signal_933}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_717 ( .s (signal_1000), .b ({key_s1[66], key_s0[66]}), .a ({key_s1[2], key_s0[2]}), .c ({signal_1247, signal_932}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_718 ( .s (signal_693), .b ({key_s1[67], key_s0[67]}), .a ({key_s1[3], key_s0[3]}), .c ({signal_1562, signal_931}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_719 ( .s (signal_693), .b ({key_s1[68], key_s0[68]}), .a ({key_s1[4], key_s0[4]}), .c ({signal_1565, signal_930}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_720 ( .s (signal_693), .b ({key_s1[69], key_s0[69]}), .a ({key_s1[5], key_s0[5]}), .c ({signal_1568, signal_929}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_721 ( .s (signal_693), .b ({key_s1[70], key_s0[70]}), .a ({key_s1[6], key_s0[6]}), .c ({signal_1571, signal_928}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_722 ( .s (signal_693), .b ({key_s1[71], key_s0[71]}), .a ({key_s1[7], key_s0[7]}), .c ({signal_1574, signal_927}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_723 ( .s (signal_693), .b ({key_s1[72], key_s0[72]}), .a ({key_s1[8], key_s0[8]}), .c ({signal_1577, signal_926}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_724 ( .s (signal_693), .b ({key_s1[73], key_s0[73]}), .a ({key_s1[9], key_s0[9]}), .c ({signal_1580, signal_925}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_725 ( .s (signal_693), .b ({key_s1[74], key_s0[74]}), .a ({key_s1[10], key_s0[10]}), .c ({signal_1583, signal_924}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_726 ( .s (signal_693), .b ({key_s1[75], key_s0[75]}), .a ({key_s1[11], key_s0[11]}), .c ({signal_1586, signal_923}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_727 ( .s (signal_693), .b ({key_s1[76], key_s0[76]}), .a ({key_s1[12], key_s0[12]}), .c ({signal_1589, signal_922}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_728 ( .s (signal_693), .b ({key_s1[77], key_s0[77]}), .a ({key_s1[13], key_s0[13]}), .c ({signal_1592, signal_921}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_729 ( .s (signal_693), .b ({key_s1[78], key_s0[78]}), .a ({key_s1[14], key_s0[14]}), .c ({signal_1595, signal_920}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_730 ( .s (signal_693), .b ({key_s1[79], key_s0[79]}), .a ({key_s1[15], key_s0[15]}), .c ({signal_1598, signal_919}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_731 ( .s (signal_693), .b ({key_s1[80], key_s0[80]}), .a ({key_s1[16], key_s0[16]}), .c ({signal_1601, signal_918}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_732 ( .s (signal_693), .b ({key_s1[81], key_s0[81]}), .a ({key_s1[17], key_s0[17]}), .c ({signal_1604, signal_917}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_733 ( .s (signal_693), .b ({key_s1[82], key_s0[82]}), .a ({key_s1[18], key_s0[18]}), .c ({signal_1607, signal_916}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_734 ( .s (signal_693), .b ({key_s1[83], key_s0[83]}), .a ({key_s1[19], key_s0[19]}), .c ({signal_1610, signal_915}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_735 ( .s (signal_693), .b ({key_s1[84], key_s0[84]}), .a ({key_s1[20], key_s0[20]}), .c ({signal_1613, signal_914}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_736 ( .s (signal_693), .b ({key_s1[85], key_s0[85]}), .a ({key_s1[21], key_s0[21]}), .c ({signal_1616, signal_913}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_737 ( .s (signal_1000), .b ({key_s1[86], key_s0[86]}), .a ({key_s1[22], key_s0[22]}), .c ({signal_1250, signal_912}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_738 ( .s (signal_1000), .b ({key_s1[87], key_s0[87]}), .a ({key_s1[23], key_s0[23]}), .c ({signal_1253, signal_911}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_739 ( .s (signal_1000), .b ({key_s1[88], key_s0[88]}), .a ({key_s1[24], key_s0[24]}), .c ({signal_1256, signal_910}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_740 ( .s (signal_1000), .b ({key_s1[89], key_s0[89]}), .a ({key_s1[25], key_s0[25]}), .c ({signal_1259, signal_909}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_741 ( .s (signal_1000), .b ({key_s1[90], key_s0[90]}), .a ({key_s1[26], key_s0[26]}), .c ({signal_1262, signal_908}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_742 ( .s (signal_1000), .b ({key_s1[91], key_s0[91]}), .a ({key_s1[27], key_s0[27]}), .c ({signal_1265, signal_907}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_743 ( .s (signal_694), .b ({key_s1[92], key_s0[92]}), .a ({key_s1[28], key_s0[28]}), .c ({signal_1619, signal_906}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_744 ( .s (signal_694), .b ({key_s1[93], key_s0[93]}), .a ({key_s1[29], key_s0[29]}), .c ({signal_1622, signal_905}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_745 ( .s (signal_694), .b ({key_s1[94], key_s0[94]}), .a ({key_s1[30], key_s0[30]}), .c ({signal_1625, signal_904}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_746 ( .s (signal_694), .b ({key_s1[95], key_s0[95]}), .a ({key_s1[31], key_s0[31]}), .c ({signal_1628, signal_903}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_747 ( .s (signal_694), .b ({key_s1[96], key_s0[96]}), .a ({key_s1[32], key_s0[32]}), .c ({signal_1631, signal_902}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_748 ( .s (signal_1000), .b ({key_s1[97], key_s0[97]}), .a ({key_s1[33], key_s0[33]}), .c ({signal_1268, signal_901}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_749 ( .s (signal_694), .b ({key_s1[98], key_s0[98]}), .a ({key_s1[34], key_s0[34]}), .c ({signal_1634, signal_900}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_750 ( .s (signal_694), .b ({key_s1[99], key_s0[99]}), .a ({key_s1[35], key_s0[35]}), .c ({signal_1637, signal_899}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_751 ( .s (signal_1000), .b ({key_s1[100], key_s0[100]}), .a ({key_s1[36], key_s0[36]}), .c ({signal_1271, signal_898}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_752 ( .s (signal_694), .b ({key_s1[101], key_s0[101]}), .a ({key_s1[37], key_s0[37]}), .c ({signal_1640, signal_897}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_753 ( .s (signal_694), .b ({key_s1[102], key_s0[102]}), .a ({key_s1[38], key_s0[38]}), .c ({signal_1643, signal_896}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_754 ( .s (signal_1000), .b ({key_s1[103], key_s0[103]}), .a ({key_s1[39], key_s0[39]}), .c ({signal_1274, signal_895}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_755 ( .s (signal_694), .b ({key_s1[104], key_s0[104]}), .a ({key_s1[40], key_s0[40]}), .c ({signal_1646, signal_894}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_756 ( .s (signal_694), .b ({key_s1[105], key_s0[105]}), .a ({key_s1[41], key_s0[41]}), .c ({signal_1649, signal_893}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_757 ( .s (signal_694), .b ({key_s1[106], key_s0[106]}), .a ({key_s1[42], key_s0[42]}), .c ({signal_1652, signal_892}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_758 ( .s (signal_694), .b ({key_s1[107], key_s0[107]}), .a ({key_s1[43], key_s0[43]}), .c ({signal_1655, signal_891}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_759 ( .s (signal_694), .b ({key_s1[108], key_s0[108]}), .a ({key_s1[44], key_s0[44]}), .c ({signal_1658, signal_890}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_760 ( .s (signal_694), .b ({key_s1[109], key_s0[109]}), .a ({key_s1[45], key_s0[45]}), .c ({signal_1661, signal_889}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_761 ( .s (signal_694), .b ({key_s1[110], key_s0[110]}), .a ({key_s1[46], key_s0[46]}), .c ({signal_1664, signal_888}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_762 ( .s (signal_694), .b ({key_s1[111], key_s0[111]}), .a ({key_s1[47], key_s0[47]}), .c ({signal_1667, signal_887}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_763 ( .s (signal_694), .b ({key_s1[112], key_s0[112]}), .a ({key_s1[48], key_s0[48]}), .c ({signal_1670, signal_886}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_764 ( .s (signal_694), .b ({key_s1[113], key_s0[113]}), .a ({key_s1[49], key_s0[49]}), .c ({signal_1673, signal_885}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_765 ( .s (signal_694), .b ({key_s1[114], key_s0[114]}), .a ({key_s1[50], key_s0[50]}), .c ({signal_1676, signal_884}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_766 ( .s (signal_694), .b ({key_s1[115], key_s0[115]}), .a ({key_s1[51], key_s0[51]}), .c ({signal_1679, signal_883}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_767 ( .s (signal_694), .b ({key_s1[116], key_s0[116]}), .a ({key_s1[52], key_s0[52]}), .c ({signal_1682, signal_882}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_768 ( .s (signal_1000), .b ({key_s1[117], key_s0[117]}), .a ({key_s1[53], key_s0[53]}), .c ({signal_1277, signal_881}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_769 ( .s (signal_1000), .b ({key_s1[118], key_s0[118]}), .a ({key_s1[54], key_s0[54]}), .c ({signal_1280, signal_880}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_770 ( .s (signal_694), .b ({key_s1[119], key_s0[119]}), .a ({key_s1[55], key_s0[55]}), .c ({signal_1685, signal_879}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_771 ( .s (signal_1000), .b ({key_s1[120], key_s0[120]}), .a ({key_s1[56], key_s0[56]}), .c ({signal_1283, signal_878}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_772 ( .s (signal_694), .b ({key_s1[121], key_s0[121]}), .a ({key_s1[57], key_s0[57]}), .c ({signal_1688, signal_877}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_773 ( .s (signal_694), .b ({key_s1[122], key_s0[122]}), .a ({key_s1[58], key_s0[58]}), .c ({signal_1691, signal_876}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_774 ( .s (signal_1000), .b ({key_s1[123], key_s0[123]}), .a ({key_s1[59], key_s0[59]}), .c ({signal_1286, signal_875}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_775 ( .s (signal_694), .b ({key_s1[124], key_s0[124]}), .a ({key_s1[60], key_s0[60]}), .c ({signal_1694, signal_874}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_776 ( .s (signal_694), .b ({key_s1[125], key_s0[125]}), .a ({key_s1[61], key_s0[61]}), .c ({signal_1697, signal_873}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_777 ( .s (signal_1000), .b ({key_s1[126], key_s0[126]}), .a ({key_s1[62], key_s0[62]}), .c ({signal_1289, signal_872}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_778 ( .s (signal_694), .b ({key_s1[127], key_s0[127]}), .a ({key_s1[63], key_s0[63]}), .c ({signal_1700, signal_871}) ) ;
    MUX2_X1 cell_779 ( .S (rst), .A (signal_1007), .B (1'b1), .Z (signal_266) ) ;
    MUX2_X1 cell_780 ( .S (rst), .A (signal_1006), .B (1'b0), .Z (signal_1014) ) ;
    MUX2_X1 cell_781 ( .S (rst), .A (signal_1005), .B (1'b0), .Z (signal_1013) ) ;
    MUX2_X1 cell_782 ( .S (rst), .A (signal_1004), .B (1'b1), .Z (signal_265) ) ;
    MUX2_X1 cell_783 ( .S (rst), .A (signal_1003), .B (1'b0), .Z (signal_1011) ) ;
    MUX2_X1 cell_784 ( .S (rst), .A (signal_1002), .B (1'b0), .Z (signal_1010) ) ;
    MUX2_X1 cell_785 ( .S (rst), .A (signal_1001), .B (1'b0), .Z (signal_1009) ) ;
    XOR2_X1 cell_786 ( .A (signal_265), .B (signal_1011), .Z (signal_1008) ) ;
    XOR2_X1 cell_787 ( .A (signal_1014), .B (signal_266), .Z (signal_1012) ) ;
    AND2_X1 cell_802 ( .A1 (signal_1009), .A2 (signal_702), .ZN (signal_267) ) ;
    NOR2_X1 cell_803 ( .A1 (signal_703), .A2 (signal_704), .ZN (signal_702) ) ;
    NAND2_X1 cell_804 ( .A1 (signal_705), .A2 (signal_706), .ZN (signal_704) ) ;
    NOR2_X1 cell_805 ( .A1 (signal_1011), .A2 (signal_1010), .ZN (signal_706) ) ;
    NOR2_X1 cell_806 ( .A1 (signal_1014), .A2 (signal_265), .ZN (signal_705) ) ;
    NAND2_X1 cell_807 ( .A1 (signal_266), .A2 (signal_1013), .ZN (signal_703) ) ;
    MUX2_X1 cell_808 ( .S (rst), .A (signal_1016), .B (1'b0), .Z (signal_1000) ) ;
    MUX2_X1 cell_809 ( .S (rst), .A (signal_1015), .B (1'b0), .Z (signal_999) ) ;
    XNOR2_X1 cell_810 ( .A (signal_707), .B (signal_999), .ZN (signal_1017) ) ;
    XNOR2_X1 cell_811 ( .A (signal_1000), .B (1'b0), .ZN (signal_707) ) ;
    INV_X1 cell_812 ( .A (signal_1000), .ZN (signal_1018) ) ;

    /* cells in depth 1 */
    buf_clk cell_1048 ( .C (clk), .D (ciphertext_s0[42]), .Q (signal_2242) ) ;
    buf_clk cell_1050 ( .C (clk), .D (ciphertext_s1[42]), .Q (signal_2244) ) ;
    buf_clk cell_1052 ( .C (clk), .D (ciphertext_s0[19]), .Q (signal_2246) ) ;
    buf_clk cell_1054 ( .C (clk), .D (ciphertext_s1[19]), .Q (signal_2248) ) ;
    buf_clk cell_1056 ( .C (clk), .D (ciphertext_s0[52]), .Q (signal_2250) ) ;
    buf_clk cell_1058 ( .C (clk), .D (ciphertext_s1[52]), .Q (signal_2252) ) ;
    buf_clk cell_1060 ( .C (clk), .D (ciphertext_s0[36]), .Q (signal_2254) ) ;
    buf_clk cell_1062 ( .C (clk), .D (ciphertext_s1[36]), .Q (signal_2256) ) ;
    buf_clk cell_1064 ( .C (clk), .D (ciphertext_s0[48]), .Q (signal_2258) ) ;
    buf_clk cell_1066 ( .C (clk), .D (ciphertext_s1[48]), .Q (signal_2260) ) ;
    buf_clk cell_1068 ( .C (clk), .D (ciphertext_s0[34]), .Q (signal_2262) ) ;
    buf_clk cell_1070 ( .C (clk), .D (ciphertext_s1[34]), .Q (signal_2264) ) ;
    buf_clk cell_1072 ( .C (clk), .D (ciphertext_s0[30]), .Q (signal_2266) ) ;
    buf_clk cell_1074 ( .C (clk), .D (ciphertext_s1[30]), .Q (signal_2268) ) ;
    buf_clk cell_1076 ( .C (clk), .D (ciphertext_s0[44]), .Q (signal_2270) ) ;
    buf_clk cell_1078 ( .C (clk), .D (ciphertext_s1[44]), .Q (signal_2272) ) ;
    buf_clk cell_1080 ( .C (clk), .D (ciphertext_s0[58]), .Q (signal_2274) ) ;
    buf_clk cell_1082 ( .C (clk), .D (ciphertext_s1[58]), .Q (signal_2276) ) ;
    buf_clk cell_1084 ( .C (clk), .D (ciphertext_s0[56]), .Q (signal_2278) ) ;
    buf_clk cell_1086 ( .C (clk), .D (ciphertext_s1[56]), .Q (signal_2280) ) ;
    buf_clk cell_1088 ( .C (clk), .D (ciphertext_s0[46]), .Q (signal_2282) ) ;
    buf_clk cell_1090 ( .C (clk), .D (ciphertext_s1[46]), .Q (signal_2284) ) ;
    buf_clk cell_1092 ( .C (clk), .D (ciphertext_s0[54]), .Q (signal_2286) ) ;
    buf_clk cell_1094 ( .C (clk), .D (ciphertext_s1[54]), .Q (signal_2288) ) ;
    buf_clk cell_1096 ( .C (clk), .D (ciphertext_s0[62]), .Q (signal_2290) ) ;
    buf_clk cell_1098 ( .C (clk), .D (ciphertext_s1[62]), .Q (signal_2292) ) ;
    buf_clk cell_1100 ( .C (clk), .D (ciphertext_s0[50]), .Q (signal_2294) ) ;
    buf_clk cell_1102 ( .C (clk), .D (ciphertext_s1[50]), .Q (signal_2296) ) ;
    buf_clk cell_1104 ( .C (clk), .D (ciphertext_s0[38]), .Q (signal_2298) ) ;
    buf_clk cell_1106 ( .C (clk), .D (ciphertext_s1[38]), .Q (signal_2300) ) ;
    buf_clk cell_1108 ( .C (clk), .D (ciphertext_s0[40]), .Q (signal_2302) ) ;
    buf_clk cell_1110 ( .C (clk), .D (ciphertext_s1[40]), .Q (signal_2304) ) ;
    buf_clk cell_1112 ( .C (clk), .D (ciphertext_s0[60]), .Q (signal_2306) ) ;
    buf_clk cell_1114 ( .C (clk), .D (ciphertext_s1[60]), .Q (signal_2308) ) ;
    buf_clk cell_1116 ( .C (clk), .D (ciphertext_s0[16]), .Q (signal_2310) ) ;
    buf_clk cell_1118 ( .C (clk), .D (ciphertext_s1[16]), .Q (signal_2312) ) ;
    buf_clk cell_1120 ( .C (clk), .D (ciphertext_s0[28]), .Q (signal_2314) ) ;
    buf_clk cell_1122 ( .C (clk), .D (ciphertext_s1[28]), .Q (signal_2316) ) ;
    buf_clk cell_1124 ( .C (clk), .D (ciphertext_s0[32]), .Q (signal_2318) ) ;
    buf_clk cell_1126 ( .C (clk), .D (ciphertext_s1[32]), .Q (signal_2320) ) ;
    buf_clk cell_1128 ( .C (clk), .D (ciphertext_s0[26]), .Q (signal_2322) ) ;
    buf_clk cell_1130 ( .C (clk), .D (ciphertext_s1[26]), .Q (signal_2324) ) ;
    buf_clk cell_1132 ( .C (clk), .D (ciphertext_s0[24]), .Q (signal_2326) ) ;
    buf_clk cell_1134 ( .C (clk), .D (ciphertext_s1[24]), .Q (signal_2328) ) ;
    buf_clk cell_1136 ( .C (clk), .D (ciphertext_s0[23]), .Q (signal_2330) ) ;
    buf_clk cell_1138 ( .C (clk), .D (ciphertext_s1[23]), .Q (signal_2332) ) ;
    buf_clk cell_1140 ( .C (clk), .D (ciphertext_s0[20]), .Q (signal_2334) ) ;
    buf_clk cell_1142 ( .C (clk), .D (ciphertext_s1[20]), .Q (signal_2336) ) ;
    buf_clk cell_1144 ( .C (clk), .D (ciphertext_s0[7]), .Q (signal_2338) ) ;
    buf_clk cell_1146 ( .C (clk), .D (ciphertext_s1[7]), .Q (signal_2340) ) ;
    buf_clk cell_1148 ( .C (clk), .D (ciphertext_s0[4]), .Q (signal_2342) ) ;
    buf_clk cell_1150 ( .C (clk), .D (ciphertext_s1[4]), .Q (signal_2344) ) ;
    buf_clk cell_1152 ( .C (clk), .D (ciphertext_s0[11]), .Q (signal_2346) ) ;
    buf_clk cell_1154 ( .C (clk), .D (ciphertext_s1[11]), .Q (signal_2348) ) ;
    buf_clk cell_1156 ( .C (clk), .D (ciphertext_s0[8]), .Q (signal_2350) ) ;
    buf_clk cell_1158 ( .C (clk), .D (ciphertext_s1[8]), .Q (signal_2352) ) ;
    buf_clk cell_1160 ( .C (clk), .D (ciphertext_s0[15]), .Q (signal_2354) ) ;
    buf_clk cell_1162 ( .C (clk), .D (ciphertext_s1[15]), .Q (signal_2356) ) ;
    buf_clk cell_1164 ( .C (clk), .D (ciphertext_s0[12]), .Q (signal_2358) ) ;
    buf_clk cell_1166 ( .C (clk), .D (ciphertext_s1[12]), .Q (signal_2360) ) ;
    buf_clk cell_1168 ( .C (clk), .D (ciphertext_s0[2]), .Q (signal_2362) ) ;
    buf_clk cell_1170 ( .C (clk), .D (ciphertext_s1[2]), .Q (signal_2364) ) ;
    buf_clk cell_1172 ( .C (clk), .D (ciphertext_s0[0]), .Q (signal_2366) ) ;
    buf_clk cell_1174 ( .C (clk), .D (ciphertext_s1[0]), .Q (signal_2368) ) ;
    buf_clk cell_1176 ( .C (clk), .D (rst), .Q (signal_2370) ) ;
    buf_clk cell_1182 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_2376) ) ;
    buf_clk cell_1188 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_2382) ) ;
    buf_clk cell_1194 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_2388) ) ;
    buf_clk cell_1200 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_2394) ) ;
    buf_clk cell_1206 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_2400) ) ;
    buf_clk cell_1212 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_2406) ) ;
    buf_clk cell_1218 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_2412) ) ;
    buf_clk cell_1224 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_2418) ) ;
    buf_clk cell_1230 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_2424) ) ;
    buf_clk cell_1236 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_2430) ) ;
    buf_clk cell_1242 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_2436) ) ;
    buf_clk cell_1248 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_2442) ) ;
    buf_clk cell_1254 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_2448) ) ;
    buf_clk cell_1260 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_2454) ) ;
    buf_clk cell_1266 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_2460) ) ;
    buf_clk cell_1272 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_2466) ) ;
    buf_clk cell_1278 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_2472) ) ;
    buf_clk cell_1284 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_2478) ) ;
    buf_clk cell_1290 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_2484) ) ;
    buf_clk cell_1296 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_2490) ) ;
    buf_clk cell_1302 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_2496) ) ;
    buf_clk cell_1308 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_2502) ) ;
    buf_clk cell_1314 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_2508) ) ;
    buf_clk cell_1320 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_2514) ) ;
    buf_clk cell_1326 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_2520) ) ;
    buf_clk cell_1332 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_2526) ) ;
    buf_clk cell_1338 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_2532) ) ;
    buf_clk cell_1344 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_2538) ) ;
    buf_clk cell_1350 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_2544) ) ;
    buf_clk cell_1356 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_2550) ) ;
    buf_clk cell_1362 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_2556) ) ;
    buf_clk cell_1368 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_2562) ) ;
    buf_clk cell_1374 ( .C (clk), .D (plaintext_s0[33]), .Q (signal_2568) ) ;
    buf_clk cell_1380 ( .C (clk), .D (plaintext_s1[33]), .Q (signal_2574) ) ;
    buf_clk cell_1386 ( .C (clk), .D (plaintext_s0[35]), .Q (signal_2580) ) ;
    buf_clk cell_1392 ( .C (clk), .D (plaintext_s1[35]), .Q (signal_2586) ) ;
    buf_clk cell_1398 ( .C (clk), .D (plaintext_s0[37]), .Q (signal_2592) ) ;
    buf_clk cell_1404 ( .C (clk), .D (plaintext_s1[37]), .Q (signal_2598) ) ;
    buf_clk cell_1410 ( .C (clk), .D (plaintext_s0[39]), .Q (signal_2604) ) ;
    buf_clk cell_1416 ( .C (clk), .D (plaintext_s1[39]), .Q (signal_2610) ) ;
    buf_clk cell_1422 ( .C (clk), .D (plaintext_s0[41]), .Q (signal_2616) ) ;
    buf_clk cell_1428 ( .C (clk), .D (plaintext_s1[41]), .Q (signal_2622) ) ;
    buf_clk cell_1434 ( .C (clk), .D (plaintext_s0[43]), .Q (signal_2628) ) ;
    buf_clk cell_1440 ( .C (clk), .D (plaintext_s1[43]), .Q (signal_2634) ) ;
    buf_clk cell_1446 ( .C (clk), .D (plaintext_s0[45]), .Q (signal_2640) ) ;
    buf_clk cell_1452 ( .C (clk), .D (plaintext_s1[45]), .Q (signal_2646) ) ;
    buf_clk cell_1458 ( .C (clk), .D (plaintext_s0[47]), .Q (signal_2652) ) ;
    buf_clk cell_1464 ( .C (clk), .D (plaintext_s1[47]), .Q (signal_2658) ) ;
    buf_clk cell_1470 ( .C (clk), .D (plaintext_s0[49]), .Q (signal_2664) ) ;
    buf_clk cell_1476 ( .C (clk), .D (plaintext_s1[49]), .Q (signal_2670) ) ;
    buf_clk cell_1482 ( .C (clk), .D (plaintext_s0[51]), .Q (signal_2676) ) ;
    buf_clk cell_1488 ( .C (clk), .D (plaintext_s1[51]), .Q (signal_2682) ) ;
    buf_clk cell_1494 ( .C (clk), .D (plaintext_s0[53]), .Q (signal_2688) ) ;
    buf_clk cell_1500 ( .C (clk), .D (plaintext_s1[53]), .Q (signal_2694) ) ;
    buf_clk cell_1506 ( .C (clk), .D (plaintext_s0[55]), .Q (signal_2700) ) ;
    buf_clk cell_1512 ( .C (clk), .D (plaintext_s1[55]), .Q (signal_2706) ) ;
    buf_clk cell_1518 ( .C (clk), .D (plaintext_s0[57]), .Q (signal_2712) ) ;
    buf_clk cell_1524 ( .C (clk), .D (plaintext_s1[57]), .Q (signal_2718) ) ;
    buf_clk cell_1530 ( .C (clk), .D (plaintext_s0[59]), .Q (signal_2724) ) ;
    buf_clk cell_1536 ( .C (clk), .D (plaintext_s1[59]), .Q (signal_2730) ) ;
    buf_clk cell_1542 ( .C (clk), .D (plaintext_s0[61]), .Q (signal_2736) ) ;
    buf_clk cell_1548 ( .C (clk), .D (plaintext_s1[61]), .Q (signal_2742) ) ;
    buf_clk cell_1554 ( .C (clk), .D (plaintext_s0[63]), .Q (signal_2748) ) ;
    buf_clk cell_1560 ( .C (clk), .D (plaintext_s1[63]), .Q (signal_2754) ) ;
    buf_clk cell_1566 ( .C (clk), .D (signal_885), .Q (signal_2760) ) ;
    buf_clk cell_1572 ( .C (clk), .D (signal_1673), .Q (signal_2766) ) ;
    buf_clk cell_1578 ( .C (clk), .D (signal_883), .Q (signal_2772) ) ;
    buf_clk cell_1584 ( .C (clk), .D (signal_1679), .Q (signal_2778) ) ;
    buf_clk cell_1590 ( .C (clk), .D (signal_881), .Q (signal_2784) ) ;
    buf_clk cell_1596 ( .C (clk), .D (signal_1277), .Q (signal_2790) ) ;
    buf_clk cell_1602 ( .C (clk), .D (signal_879), .Q (signal_2796) ) ;
    buf_clk cell_1608 ( .C (clk), .D (signal_1685), .Q (signal_2802) ) ;
    buf_clk cell_1614 ( .C (clk), .D (signal_877), .Q (signal_2808) ) ;
    buf_clk cell_1620 ( .C (clk), .D (signal_1688), .Q (signal_2814) ) ;
    buf_clk cell_1626 ( .C (clk), .D (signal_875), .Q (signal_2820) ) ;
    buf_clk cell_1632 ( .C (clk), .D (signal_1286), .Q (signal_2826) ) ;
    buf_clk cell_1638 ( .C (clk), .D (signal_873), .Q (signal_2832) ) ;
    buf_clk cell_1644 ( .C (clk), .D (signal_1697), .Q (signal_2838) ) ;
    buf_clk cell_1650 ( .C (clk), .D (signal_871), .Q (signal_2844) ) ;
    buf_clk cell_1656 ( .C (clk), .D (signal_1700), .Q (signal_2850) ) ;
    buf_clk cell_1662 ( .C (clk), .D (signal_335), .Q (signal_2856) ) ;
    buf_clk cell_1668 ( .C (clk), .D (signal_1822), .Q (signal_2862) ) ;
    buf_clk cell_1674 ( .C (clk), .D (signal_339), .Q (signal_2868) ) ;
    buf_clk cell_1680 ( .C (clk), .D (signal_1824), .Q (signal_2874) ) ;
    buf_clk cell_1686 ( .C (clk), .D (signal_343), .Q (signal_2880) ) ;
    buf_clk cell_1692 ( .C (clk), .D (signal_1826), .Q (signal_2886) ) ;
    buf_clk cell_1698 ( .C (clk), .D (signal_347), .Q (signal_2892) ) ;
    buf_clk cell_1704 ( .C (clk), .D (signal_1828), .Q (signal_2898) ) ;
    buf_clk cell_1710 ( .C (clk), .D (signal_933), .Q (signal_2904) ) ;
    buf_clk cell_1716 ( .C (clk), .D (signal_1559), .Q (signal_2910) ) ;
    buf_clk cell_1722 ( .C (clk), .D (signal_931), .Q (signal_2916) ) ;
    buf_clk cell_1728 ( .C (clk), .D (signal_1562), .Q (signal_2922) ) ;
    buf_clk cell_1734 ( .C (clk), .D (signal_929), .Q (signal_2928) ) ;
    buf_clk cell_1740 ( .C (clk), .D (signal_1568), .Q (signal_2934) ) ;
    buf_clk cell_1746 ( .C (clk), .D (signal_927), .Q (signal_2940) ) ;
    buf_clk cell_1752 ( .C (clk), .D (signal_1574), .Q (signal_2946) ) ;
    buf_clk cell_1758 ( .C (clk), .D (signal_925), .Q (signal_2952) ) ;
    buf_clk cell_1764 ( .C (clk), .D (signal_1580), .Q (signal_2958) ) ;
    buf_clk cell_1770 ( .C (clk), .D (signal_923), .Q (signal_2964) ) ;
    buf_clk cell_1776 ( .C (clk), .D (signal_1586), .Q (signal_2970) ) ;
    buf_clk cell_1782 ( .C (clk), .D (signal_921), .Q (signal_2976) ) ;
    buf_clk cell_1788 ( .C (clk), .D (signal_1592), .Q (signal_2982) ) ;
    buf_clk cell_1794 ( .C (clk), .D (signal_919), .Q (signal_2988) ) ;
    buf_clk cell_1800 ( .C (clk), .D (signal_1598), .Q (signal_2994) ) ;
    buf_clk cell_1806 ( .C (clk), .D (signal_917), .Q (signal_3000) ) ;
    buf_clk cell_1812 ( .C (clk), .D (signal_1604), .Q (signal_3006) ) ;
    buf_clk cell_1818 ( .C (clk), .D (signal_915), .Q (signal_3012) ) ;
    buf_clk cell_1824 ( .C (clk), .D (signal_1610), .Q (signal_3018) ) ;
    buf_clk cell_1830 ( .C (clk), .D (signal_913), .Q (signal_3024) ) ;
    buf_clk cell_1836 ( .C (clk), .D (signal_1616), .Q (signal_3030) ) ;
    buf_clk cell_1842 ( .C (clk), .D (signal_911), .Q (signal_3036) ) ;
    buf_clk cell_1848 ( .C (clk), .D (signal_1253), .Q (signal_3042) ) ;
    buf_clk cell_1854 ( .C (clk), .D (signal_909), .Q (signal_3048) ) ;
    buf_clk cell_1860 ( .C (clk), .D (signal_1259), .Q (signal_3054) ) ;
    buf_clk cell_1866 ( .C (clk), .D (signal_907), .Q (signal_3060) ) ;
    buf_clk cell_1872 ( .C (clk), .D (signal_1265), .Q (signal_3066) ) ;
    buf_clk cell_1878 ( .C (clk), .D (signal_905), .Q (signal_3072) ) ;
    buf_clk cell_1884 ( .C (clk), .D (signal_1622), .Q (signal_3078) ) ;
    buf_clk cell_1890 ( .C (clk), .D (signal_903), .Q (signal_3084) ) ;
    buf_clk cell_1896 ( .C (clk), .D (signal_1628), .Q (signal_3090) ) ;
    buf_clk cell_1902 ( .C (clk), .D (signal_901), .Q (signal_3096) ) ;
    buf_clk cell_1908 ( .C (clk), .D (signal_1268), .Q (signal_3102) ) ;
    buf_clk cell_1914 ( .C (clk), .D (signal_899), .Q (signal_3108) ) ;
    buf_clk cell_1920 ( .C (clk), .D (signal_1637), .Q (signal_3114) ) ;
    buf_clk cell_1926 ( .C (clk), .D (signal_897), .Q (signal_3120) ) ;
    buf_clk cell_1932 ( .C (clk), .D (signal_1640), .Q (signal_3126) ) ;
    buf_clk cell_1938 ( .C (clk), .D (signal_895), .Q (signal_3132) ) ;
    buf_clk cell_1944 ( .C (clk), .D (signal_1274), .Q (signal_3138) ) ;
    buf_clk cell_1954 ( .C (clk), .D (ciphertext_s0[45]), .Q (signal_3148) ) ;
    buf_clk cell_1958 ( .C (clk), .D (ciphertext_s1[45]), .Q (signal_3152) ) ;
    buf_clk cell_1986 ( .C (clk), .D (ciphertext_s0[37]), .Q (signal_3180) ) ;
    buf_clk cell_1990 ( .C (clk), .D (ciphertext_s1[37]), .Q (signal_3184) ) ;
    buf_clk cell_1994 ( .C (clk), .D (ciphertext_s0[53]), .Q (signal_3188) ) ;
    buf_clk cell_1998 ( .C (clk), .D (ciphertext_s1[53]), .Q (signal_3192) ) ;
    buf_clk cell_2010 ( .C (clk), .D (ciphertext_s0[17]), .Q (signal_3204) ) ;
    buf_clk cell_2014 ( .C (clk), .D (ciphertext_s1[17]), .Q (signal_3208) ) ;
    buf_clk cell_2018 ( .C (clk), .D (ciphertext_s0[29]), .Q (signal_3212) ) ;
    buf_clk cell_2022 ( .C (clk), .D (ciphertext_s1[29]), .Q (signal_3216) ) ;
    buf_clk cell_2030 ( .C (clk), .D (ciphertext_s0[61]), .Q (signal_3224) ) ;
    buf_clk cell_2034 ( .C (clk), .D (ciphertext_s1[61]), .Q (signal_3228) ) ;
    buf_clk cell_2038 ( .C (clk), .D (ciphertext_s0[33]), .Q (signal_3232) ) ;
    buf_clk cell_2042 ( .C (clk), .D (ciphertext_s1[33]), .Q (signal_3236) ) ;
    buf_clk cell_2046 ( .C (clk), .D (ciphertext_s0[41]), .Q (signal_3240) ) ;
    buf_clk cell_2050 ( .C (clk), .D (ciphertext_s1[41]), .Q (signal_3244) ) ;
    buf_clk cell_2054 ( .C (clk), .D (ciphertext_s0[57]), .Q (signal_3248) ) ;
    buf_clk cell_2058 ( .C (clk), .D (ciphertext_s1[57]), .Q (signal_3252) ) ;
    buf_clk cell_2062 ( .C (clk), .D (ciphertext_s0[49]), .Q (signal_3256) ) ;
    buf_clk cell_2066 ( .C (clk), .D (ciphertext_s1[49]), .Q (signal_3260) ) ;
    buf_clk cell_2074 ( .C (clk), .D (ciphertext_s0[25]), .Q (signal_3268) ) ;
    buf_clk cell_2078 ( .C (clk), .D (ciphertext_s1[25]), .Q (signal_3272) ) ;
    buf_clk cell_2086 ( .C (clk), .D (ciphertext_s0[21]), .Q (signal_3280) ) ;
    buf_clk cell_2090 ( .C (clk), .D (ciphertext_s1[21]), .Q (signal_3284) ) ;
    buf_clk cell_2098 ( .C (clk), .D (ciphertext_s0[5]), .Q (signal_3292) ) ;
    buf_clk cell_2102 ( .C (clk), .D (ciphertext_s1[5]), .Q (signal_3296) ) ;
    buf_clk cell_2110 ( .C (clk), .D (ciphertext_s0[9]), .Q (signal_3304) ) ;
    buf_clk cell_2114 ( .C (clk), .D (ciphertext_s1[9]), .Q (signal_3308) ) ;
    buf_clk cell_2122 ( .C (clk), .D (ciphertext_s0[13]), .Q (signal_3316) ) ;
    buf_clk cell_2126 ( .C (clk), .D (ciphertext_s1[13]), .Q (signal_3320) ) ;
    buf_clk cell_2134 ( .C (clk), .D (ciphertext_s0[1]), .Q (signal_3328) ) ;
    buf_clk cell_2138 ( .C (clk), .D (ciphertext_s1[1]), .Q (signal_3332) ) ;
    buf_clk cell_2144 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_3338) ) ;
    buf_clk cell_2152 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_3346) ) ;
    buf_clk cell_2160 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_3354) ) ;
    buf_clk cell_2168 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_3362) ) ;
    buf_clk cell_2176 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_3370) ) ;
    buf_clk cell_2184 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_3378) ) ;
    buf_clk cell_2192 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_3386) ) ;
    buf_clk cell_2200 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_3394) ) ;
    buf_clk cell_2208 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_3402) ) ;
    buf_clk cell_2216 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_3410) ) ;
    buf_clk cell_2224 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_3418) ) ;
    buf_clk cell_2232 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_3426) ) ;
    buf_clk cell_2240 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_3434) ) ;
    buf_clk cell_2248 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_3442) ) ;
    buf_clk cell_2256 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_3450) ) ;
    buf_clk cell_2264 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_3458) ) ;
    buf_clk cell_2272 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_3466) ) ;
    buf_clk cell_2280 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_3474) ) ;
    buf_clk cell_2288 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_3482) ) ;
    buf_clk cell_2296 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_3490) ) ;
    buf_clk cell_2304 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_3498) ) ;
    buf_clk cell_2312 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_3506) ) ;
    buf_clk cell_2320 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_3514) ) ;
    buf_clk cell_2328 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_3522) ) ;
    buf_clk cell_2336 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_3530) ) ;
    buf_clk cell_2344 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_3538) ) ;
    buf_clk cell_2352 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_3546) ) ;
    buf_clk cell_2360 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_3554) ) ;
    buf_clk cell_2368 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_3562) ) ;
    buf_clk cell_2376 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_3570) ) ;
    buf_clk cell_2384 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_3578) ) ;
    buf_clk cell_2392 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_3586) ) ;
    buf_clk cell_2400 ( .C (clk), .D (plaintext_s0[32]), .Q (signal_3594) ) ;
    buf_clk cell_2408 ( .C (clk), .D (plaintext_s1[32]), .Q (signal_3602) ) ;
    buf_clk cell_2416 ( .C (clk), .D (plaintext_s0[34]), .Q (signal_3610) ) ;
    buf_clk cell_2424 ( .C (clk), .D (plaintext_s1[34]), .Q (signal_3618) ) ;
    buf_clk cell_2432 ( .C (clk), .D (plaintext_s0[36]), .Q (signal_3626) ) ;
    buf_clk cell_2440 ( .C (clk), .D (plaintext_s1[36]), .Q (signal_3634) ) ;
    buf_clk cell_2448 ( .C (clk), .D (plaintext_s0[38]), .Q (signal_3642) ) ;
    buf_clk cell_2456 ( .C (clk), .D (plaintext_s1[38]), .Q (signal_3650) ) ;
    buf_clk cell_2464 ( .C (clk), .D (plaintext_s0[40]), .Q (signal_3658) ) ;
    buf_clk cell_2472 ( .C (clk), .D (plaintext_s1[40]), .Q (signal_3666) ) ;
    buf_clk cell_2480 ( .C (clk), .D (plaintext_s0[42]), .Q (signal_3674) ) ;
    buf_clk cell_2488 ( .C (clk), .D (plaintext_s1[42]), .Q (signal_3682) ) ;
    buf_clk cell_2496 ( .C (clk), .D (plaintext_s0[44]), .Q (signal_3690) ) ;
    buf_clk cell_2504 ( .C (clk), .D (plaintext_s1[44]), .Q (signal_3698) ) ;
    buf_clk cell_2512 ( .C (clk), .D (plaintext_s0[46]), .Q (signal_3706) ) ;
    buf_clk cell_2520 ( .C (clk), .D (plaintext_s1[46]), .Q (signal_3714) ) ;
    buf_clk cell_2528 ( .C (clk), .D (plaintext_s0[48]), .Q (signal_3722) ) ;
    buf_clk cell_2536 ( .C (clk), .D (plaintext_s1[48]), .Q (signal_3730) ) ;
    buf_clk cell_2544 ( .C (clk), .D (plaintext_s0[50]), .Q (signal_3738) ) ;
    buf_clk cell_2552 ( .C (clk), .D (plaintext_s1[50]), .Q (signal_3746) ) ;
    buf_clk cell_2560 ( .C (clk), .D (plaintext_s0[52]), .Q (signal_3754) ) ;
    buf_clk cell_2568 ( .C (clk), .D (plaintext_s1[52]), .Q (signal_3762) ) ;
    buf_clk cell_2576 ( .C (clk), .D (plaintext_s0[54]), .Q (signal_3770) ) ;
    buf_clk cell_2584 ( .C (clk), .D (plaintext_s1[54]), .Q (signal_3778) ) ;
    buf_clk cell_2592 ( .C (clk), .D (plaintext_s0[56]), .Q (signal_3786) ) ;
    buf_clk cell_2600 ( .C (clk), .D (plaintext_s1[56]), .Q (signal_3794) ) ;
    buf_clk cell_2608 ( .C (clk), .D (plaintext_s0[58]), .Q (signal_3802) ) ;
    buf_clk cell_2616 ( .C (clk), .D (plaintext_s1[58]), .Q (signal_3810) ) ;
    buf_clk cell_2624 ( .C (clk), .D (plaintext_s0[60]), .Q (signal_3818) ) ;
    buf_clk cell_2632 ( .C (clk), .D (plaintext_s1[60]), .Q (signal_3826) ) ;
    buf_clk cell_2640 ( .C (clk), .D (plaintext_s0[62]), .Q (signal_3834) ) ;
    buf_clk cell_2648 ( .C (clk), .D (plaintext_s1[62]), .Q (signal_3842) ) ;
    buf_clk cell_2656 ( .C (clk), .D (signal_886), .Q (signal_3850) ) ;
    buf_clk cell_2664 ( .C (clk), .D (signal_1670), .Q (signal_3858) ) ;
    buf_clk cell_2672 ( .C (clk), .D (signal_884), .Q (signal_3866) ) ;
    buf_clk cell_2680 ( .C (clk), .D (signal_1676), .Q (signal_3874) ) ;
    buf_clk cell_2688 ( .C (clk), .D (signal_882), .Q (signal_3882) ) ;
    buf_clk cell_2696 ( .C (clk), .D (signal_1682), .Q (signal_3890) ) ;
    buf_clk cell_2704 ( .C (clk), .D (signal_880), .Q (signal_3898) ) ;
    buf_clk cell_2712 ( .C (clk), .D (signal_1280), .Q (signal_3906) ) ;
    buf_clk cell_2720 ( .C (clk), .D (signal_878), .Q (signal_3914) ) ;
    buf_clk cell_2728 ( .C (clk), .D (signal_1283), .Q (signal_3922) ) ;
    buf_clk cell_2736 ( .C (clk), .D (signal_876), .Q (signal_3930) ) ;
    buf_clk cell_2744 ( .C (clk), .D (signal_1691), .Q (signal_3938) ) ;
    buf_clk cell_2752 ( .C (clk), .D (signal_874), .Q (signal_3946) ) ;
    buf_clk cell_2760 ( .C (clk), .D (signal_1694), .Q (signal_3954) ) ;
    buf_clk cell_2768 ( .C (clk), .D (signal_872), .Q (signal_3962) ) ;
    buf_clk cell_2776 ( .C (clk), .D (signal_1289), .Q (signal_3970) ) ;
    buf_clk cell_2784 ( .C (clk), .D (signal_333), .Q (signal_3978) ) ;
    buf_clk cell_2792 ( .C (clk), .D (signal_1821), .Q (signal_3986) ) ;
    buf_clk cell_2800 ( .C (clk), .D (signal_337), .Q (signal_3994) ) ;
    buf_clk cell_2808 ( .C (clk), .D (signal_1823), .Q (signal_4002) ) ;
    buf_clk cell_2816 ( .C (clk), .D (signal_341), .Q (signal_4010) ) ;
    buf_clk cell_2824 ( .C (clk), .D (signal_1825), .Q (signal_4018) ) ;
    buf_clk cell_2832 ( .C (clk), .D (signal_345), .Q (signal_4026) ) ;
    buf_clk cell_2840 ( .C (clk), .D (signal_1827), .Q (signal_4034) ) ;
    buf_clk cell_2848 ( .C (clk), .D (signal_934), .Q (signal_4042) ) ;
    buf_clk cell_2856 ( .C (clk), .D (signal_1244), .Q (signal_4050) ) ;
    buf_clk cell_2864 ( .C (clk), .D (signal_932), .Q (signal_4058) ) ;
    buf_clk cell_2872 ( .C (clk), .D (signal_1247), .Q (signal_4066) ) ;
    buf_clk cell_2880 ( .C (clk), .D (signal_930), .Q (signal_4074) ) ;
    buf_clk cell_2888 ( .C (clk), .D (signal_1565), .Q (signal_4082) ) ;
    buf_clk cell_2896 ( .C (clk), .D (signal_928), .Q (signal_4090) ) ;
    buf_clk cell_2904 ( .C (clk), .D (signal_1571), .Q (signal_4098) ) ;
    buf_clk cell_2912 ( .C (clk), .D (signal_926), .Q (signal_4106) ) ;
    buf_clk cell_2920 ( .C (clk), .D (signal_1577), .Q (signal_4114) ) ;
    buf_clk cell_2928 ( .C (clk), .D (signal_924), .Q (signal_4122) ) ;
    buf_clk cell_2936 ( .C (clk), .D (signal_1583), .Q (signal_4130) ) ;
    buf_clk cell_2944 ( .C (clk), .D (signal_922), .Q (signal_4138) ) ;
    buf_clk cell_2952 ( .C (clk), .D (signal_1589), .Q (signal_4146) ) ;
    buf_clk cell_2960 ( .C (clk), .D (signal_920), .Q (signal_4154) ) ;
    buf_clk cell_2968 ( .C (clk), .D (signal_1595), .Q (signal_4162) ) ;
    buf_clk cell_2976 ( .C (clk), .D (signal_918), .Q (signal_4170) ) ;
    buf_clk cell_2984 ( .C (clk), .D (signal_1601), .Q (signal_4178) ) ;
    buf_clk cell_2992 ( .C (clk), .D (signal_916), .Q (signal_4186) ) ;
    buf_clk cell_3000 ( .C (clk), .D (signal_1607), .Q (signal_4194) ) ;
    buf_clk cell_3008 ( .C (clk), .D (signal_914), .Q (signal_4202) ) ;
    buf_clk cell_3016 ( .C (clk), .D (signal_1613), .Q (signal_4210) ) ;
    buf_clk cell_3024 ( .C (clk), .D (signal_912), .Q (signal_4218) ) ;
    buf_clk cell_3032 ( .C (clk), .D (signal_1250), .Q (signal_4226) ) ;
    buf_clk cell_3040 ( .C (clk), .D (signal_910), .Q (signal_4234) ) ;
    buf_clk cell_3048 ( .C (clk), .D (signal_1256), .Q (signal_4242) ) ;
    buf_clk cell_3056 ( .C (clk), .D (signal_908), .Q (signal_4250) ) ;
    buf_clk cell_3064 ( .C (clk), .D (signal_1262), .Q (signal_4258) ) ;
    buf_clk cell_3072 ( .C (clk), .D (signal_906), .Q (signal_4266) ) ;
    buf_clk cell_3080 ( .C (clk), .D (signal_1619), .Q (signal_4274) ) ;
    buf_clk cell_3088 ( .C (clk), .D (signal_904), .Q (signal_4282) ) ;
    buf_clk cell_3096 ( .C (clk), .D (signal_1625), .Q (signal_4290) ) ;
    buf_clk cell_3104 ( .C (clk), .D (signal_902), .Q (signal_4298) ) ;
    buf_clk cell_3112 ( .C (clk), .D (signal_1631), .Q (signal_4306) ) ;
    buf_clk cell_3120 ( .C (clk), .D (signal_900), .Q (signal_4314) ) ;
    buf_clk cell_3128 ( .C (clk), .D (signal_1634), .Q (signal_4322) ) ;
    buf_clk cell_3136 ( .C (clk), .D (signal_898), .Q (signal_4330) ) ;
    buf_clk cell_3144 ( .C (clk), .D (signal_1271), .Q (signal_4338) ) ;
    buf_clk cell_3152 ( .C (clk), .D (signal_896), .Q (signal_4346) ) ;
    buf_clk cell_3160 ( .C (clk), .D (signal_1643), .Q (signal_4354) ) ;
    buf_clk cell_3488 ( .C (clk), .D (signal_1008), .Q (signal_4682) ) ;
    buf_clk cell_3496 ( .C (clk), .D (signal_1009), .Q (signal_4690) ) ;
    buf_clk cell_3504 ( .C (clk), .D (signal_1010), .Q (signal_4698) ) ;
    buf_clk cell_3512 ( .C (clk), .D (signal_1011), .Q (signal_4706) ) ;
    buf_clk cell_3520 ( .C (clk), .D (signal_1012), .Q (signal_4714) ) ;
    buf_clk cell_3528 ( .C (clk), .D (signal_1013), .Q (signal_4722) ) ;
    buf_clk cell_3536 ( .C (clk), .D (signal_1014), .Q (signal_4730) ) ;
    buf_clk cell_3544 ( .C (clk), .D (signal_1017), .Q (signal_4738) ) ;
    buf_clk cell_3552 ( .C (clk), .D (signal_1018), .Q (signal_4746) ) ;
    buf_clk cell_3560 ( .C (clk), .D (signal_267), .Q (signal_4754) ) ;

    /* cells in depth 2 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_819 ( .s ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[0]), .c ({signal_1185, signal_1019}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_820 ( .s ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[1]), .c ({signal_1187, signal_1020}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_821 ( .s ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[2]), .c ({signal_1189, signal_1021}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_822 ( .s ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[3]), .c ({signal_1191, signal_1022}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_823 ( .s ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[4]), .c ({signal_1193, signal_1023}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_824 ( .s ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[5]), .c ({signal_1194, signal_1024}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_825 ( .s ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[6]), .c ({signal_1196, signal_1025}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_826 ( .s ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[7]), .c ({signal_1198, signal_1026}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_827 ( .s ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[8]), .c ({signal_1200, signal_1027}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_828 ( .s ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[9]), .c ({signal_1202, signal_1028}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_829 ( .s ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[10]), .c ({signal_1203, signal_1029}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_830 ( .s ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[11]), .c ({signal_1205, signal_1030}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_831 ( .s ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[12]), .c ({signal_1207, signal_1031}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_832 ( .s ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[13]), .c ({signal_1208, signal_1032}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_833 ( .s ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[14]), .c ({signal_1209, signal_1033}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_834 ( .s ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[15]), .c ({signal_1210, signal_1034}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_835 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[16]), .c ({signal_1212, signal_1035}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_836 ( .s ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[17]), .c ({signal_1213, signal_1036}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_837 ( .s ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[18]), .c ({signal_1214, signal_1037}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_838 ( .s ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[19]), .c ({signal_1215, signal_1038}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_839 ( .s ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[20]), .c ({signal_1216, signal_1039}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_840 ( .s ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[21]), .c ({signal_1217, signal_1040}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_841 ( .s ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[22]), .c ({signal_1218, signal_1041}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_842 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[23]), .c ({signal_1220, signal_1042}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_843 ( .s ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[24]), .c ({signal_1221, signal_1043}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_844 ( .s ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[25]), .c ({signal_1223, signal_1044}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_845 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[26]), .c ({signal_1225, signal_1045}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_846 ( .s ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[27]), .c ({signal_1226, signal_1046}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_847 ( .s ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[28]), .c ({signal_1228, signal_1047}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_848 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[29]), .c ({signal_1230, signal_1048}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_849 ( .s ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[30]), .c ({signal_1231, signal_1049}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_850 ( .s ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[31]), .c ({signal_1233, signal_1050}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_851 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[32]), .c ({signal_1235, signal_1051}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_852 ( .s ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[33]), .c ({signal_1236, signal_1052}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_853 ( .s ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[34]), .c ({signal_1238, signal_1053}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_854 ( .s ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({1'b0, 1'b0}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[35]), .c ({signal_1240, signal_1054}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_855 ( .s ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({1'b0, 1'b1}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[36]), .c ({signal_1241, signal_1055}) ) ;
    buf_clk cell_1049 ( .C (clk), .D (signal_2242), .Q (signal_2243) ) ;
    buf_clk cell_1051 ( .C (clk), .D (signal_2244), .Q (signal_2245) ) ;
    buf_clk cell_1053 ( .C (clk), .D (signal_2246), .Q (signal_2247) ) ;
    buf_clk cell_1055 ( .C (clk), .D (signal_2248), .Q (signal_2249) ) ;
    buf_clk cell_1057 ( .C (clk), .D (signal_2250), .Q (signal_2251) ) ;
    buf_clk cell_1059 ( .C (clk), .D (signal_2252), .Q (signal_2253) ) ;
    buf_clk cell_1061 ( .C (clk), .D (signal_2254), .Q (signal_2255) ) ;
    buf_clk cell_1063 ( .C (clk), .D (signal_2256), .Q (signal_2257) ) ;
    buf_clk cell_1065 ( .C (clk), .D (signal_2258), .Q (signal_2259) ) ;
    buf_clk cell_1067 ( .C (clk), .D (signal_2260), .Q (signal_2261) ) ;
    buf_clk cell_1069 ( .C (clk), .D (signal_2262), .Q (signal_2263) ) ;
    buf_clk cell_1071 ( .C (clk), .D (signal_2264), .Q (signal_2265) ) ;
    buf_clk cell_1073 ( .C (clk), .D (signal_2266), .Q (signal_2267) ) ;
    buf_clk cell_1075 ( .C (clk), .D (signal_2268), .Q (signal_2269) ) ;
    buf_clk cell_1077 ( .C (clk), .D (signal_2270), .Q (signal_2271) ) ;
    buf_clk cell_1079 ( .C (clk), .D (signal_2272), .Q (signal_2273) ) ;
    buf_clk cell_1081 ( .C (clk), .D (signal_2274), .Q (signal_2275) ) ;
    buf_clk cell_1083 ( .C (clk), .D (signal_2276), .Q (signal_2277) ) ;
    buf_clk cell_1085 ( .C (clk), .D (signal_2278), .Q (signal_2279) ) ;
    buf_clk cell_1087 ( .C (clk), .D (signal_2280), .Q (signal_2281) ) ;
    buf_clk cell_1089 ( .C (clk), .D (signal_2282), .Q (signal_2283) ) ;
    buf_clk cell_1091 ( .C (clk), .D (signal_2284), .Q (signal_2285) ) ;
    buf_clk cell_1093 ( .C (clk), .D (signal_2286), .Q (signal_2287) ) ;
    buf_clk cell_1095 ( .C (clk), .D (signal_2288), .Q (signal_2289) ) ;
    buf_clk cell_1097 ( .C (clk), .D (signal_2290), .Q (signal_2291) ) ;
    buf_clk cell_1099 ( .C (clk), .D (signal_2292), .Q (signal_2293) ) ;
    buf_clk cell_1101 ( .C (clk), .D (signal_2294), .Q (signal_2295) ) ;
    buf_clk cell_1103 ( .C (clk), .D (signal_2296), .Q (signal_2297) ) ;
    buf_clk cell_1105 ( .C (clk), .D (signal_2298), .Q (signal_2299) ) ;
    buf_clk cell_1107 ( .C (clk), .D (signal_2300), .Q (signal_2301) ) ;
    buf_clk cell_1109 ( .C (clk), .D (signal_2302), .Q (signal_2303) ) ;
    buf_clk cell_1111 ( .C (clk), .D (signal_2304), .Q (signal_2305) ) ;
    buf_clk cell_1113 ( .C (clk), .D (signal_2306), .Q (signal_2307) ) ;
    buf_clk cell_1115 ( .C (clk), .D (signal_2308), .Q (signal_2309) ) ;
    buf_clk cell_1117 ( .C (clk), .D (signal_2310), .Q (signal_2311) ) ;
    buf_clk cell_1119 ( .C (clk), .D (signal_2312), .Q (signal_2313) ) ;
    buf_clk cell_1121 ( .C (clk), .D (signal_2314), .Q (signal_2315) ) ;
    buf_clk cell_1123 ( .C (clk), .D (signal_2316), .Q (signal_2317) ) ;
    buf_clk cell_1125 ( .C (clk), .D (signal_2318), .Q (signal_2319) ) ;
    buf_clk cell_1127 ( .C (clk), .D (signal_2320), .Q (signal_2321) ) ;
    buf_clk cell_1129 ( .C (clk), .D (signal_2322), .Q (signal_2323) ) ;
    buf_clk cell_1131 ( .C (clk), .D (signal_2324), .Q (signal_2325) ) ;
    buf_clk cell_1133 ( .C (clk), .D (signal_2326), .Q (signal_2327) ) ;
    buf_clk cell_1135 ( .C (clk), .D (signal_2328), .Q (signal_2329) ) ;
    buf_clk cell_1137 ( .C (clk), .D (signal_2330), .Q (signal_2331) ) ;
    buf_clk cell_1139 ( .C (clk), .D (signal_2332), .Q (signal_2333) ) ;
    buf_clk cell_1141 ( .C (clk), .D (signal_2334), .Q (signal_2335) ) ;
    buf_clk cell_1143 ( .C (clk), .D (signal_2336), .Q (signal_2337) ) ;
    buf_clk cell_1145 ( .C (clk), .D (signal_2338), .Q (signal_2339) ) ;
    buf_clk cell_1147 ( .C (clk), .D (signal_2340), .Q (signal_2341) ) ;
    buf_clk cell_1149 ( .C (clk), .D (signal_2342), .Q (signal_2343) ) ;
    buf_clk cell_1151 ( .C (clk), .D (signal_2344), .Q (signal_2345) ) ;
    buf_clk cell_1153 ( .C (clk), .D (signal_2346), .Q (signal_2347) ) ;
    buf_clk cell_1155 ( .C (clk), .D (signal_2348), .Q (signal_2349) ) ;
    buf_clk cell_1157 ( .C (clk), .D (signal_2350), .Q (signal_2351) ) ;
    buf_clk cell_1159 ( .C (clk), .D (signal_2352), .Q (signal_2353) ) ;
    buf_clk cell_1161 ( .C (clk), .D (signal_2354), .Q (signal_2355) ) ;
    buf_clk cell_1163 ( .C (clk), .D (signal_2356), .Q (signal_2357) ) ;
    buf_clk cell_1165 ( .C (clk), .D (signal_2358), .Q (signal_2359) ) ;
    buf_clk cell_1167 ( .C (clk), .D (signal_2360), .Q (signal_2361) ) ;
    buf_clk cell_1169 ( .C (clk), .D (signal_2362), .Q (signal_2363) ) ;
    buf_clk cell_1171 ( .C (clk), .D (signal_2364), .Q (signal_2365) ) ;
    buf_clk cell_1173 ( .C (clk), .D (signal_2366), .Q (signal_2367) ) ;
    buf_clk cell_1175 ( .C (clk), .D (signal_2368), .Q (signal_2369) ) ;
    buf_clk cell_1177 ( .C (clk), .D (signal_2370), .Q (signal_2371) ) ;
    buf_clk cell_1183 ( .C (clk), .D (signal_2376), .Q (signal_2377) ) ;
    buf_clk cell_1189 ( .C (clk), .D (signal_2382), .Q (signal_2383) ) ;
    buf_clk cell_1195 ( .C (clk), .D (signal_2388), .Q (signal_2389) ) ;
    buf_clk cell_1201 ( .C (clk), .D (signal_2394), .Q (signal_2395) ) ;
    buf_clk cell_1207 ( .C (clk), .D (signal_2400), .Q (signal_2401) ) ;
    buf_clk cell_1213 ( .C (clk), .D (signal_2406), .Q (signal_2407) ) ;
    buf_clk cell_1219 ( .C (clk), .D (signal_2412), .Q (signal_2413) ) ;
    buf_clk cell_1225 ( .C (clk), .D (signal_2418), .Q (signal_2419) ) ;
    buf_clk cell_1231 ( .C (clk), .D (signal_2424), .Q (signal_2425) ) ;
    buf_clk cell_1237 ( .C (clk), .D (signal_2430), .Q (signal_2431) ) ;
    buf_clk cell_1243 ( .C (clk), .D (signal_2436), .Q (signal_2437) ) ;
    buf_clk cell_1249 ( .C (clk), .D (signal_2442), .Q (signal_2443) ) ;
    buf_clk cell_1255 ( .C (clk), .D (signal_2448), .Q (signal_2449) ) ;
    buf_clk cell_1261 ( .C (clk), .D (signal_2454), .Q (signal_2455) ) ;
    buf_clk cell_1267 ( .C (clk), .D (signal_2460), .Q (signal_2461) ) ;
    buf_clk cell_1273 ( .C (clk), .D (signal_2466), .Q (signal_2467) ) ;
    buf_clk cell_1279 ( .C (clk), .D (signal_2472), .Q (signal_2473) ) ;
    buf_clk cell_1285 ( .C (clk), .D (signal_2478), .Q (signal_2479) ) ;
    buf_clk cell_1291 ( .C (clk), .D (signal_2484), .Q (signal_2485) ) ;
    buf_clk cell_1297 ( .C (clk), .D (signal_2490), .Q (signal_2491) ) ;
    buf_clk cell_1303 ( .C (clk), .D (signal_2496), .Q (signal_2497) ) ;
    buf_clk cell_1309 ( .C (clk), .D (signal_2502), .Q (signal_2503) ) ;
    buf_clk cell_1315 ( .C (clk), .D (signal_2508), .Q (signal_2509) ) ;
    buf_clk cell_1321 ( .C (clk), .D (signal_2514), .Q (signal_2515) ) ;
    buf_clk cell_1327 ( .C (clk), .D (signal_2520), .Q (signal_2521) ) ;
    buf_clk cell_1333 ( .C (clk), .D (signal_2526), .Q (signal_2527) ) ;
    buf_clk cell_1339 ( .C (clk), .D (signal_2532), .Q (signal_2533) ) ;
    buf_clk cell_1345 ( .C (clk), .D (signal_2538), .Q (signal_2539) ) ;
    buf_clk cell_1351 ( .C (clk), .D (signal_2544), .Q (signal_2545) ) ;
    buf_clk cell_1357 ( .C (clk), .D (signal_2550), .Q (signal_2551) ) ;
    buf_clk cell_1363 ( .C (clk), .D (signal_2556), .Q (signal_2557) ) ;
    buf_clk cell_1369 ( .C (clk), .D (signal_2562), .Q (signal_2563) ) ;
    buf_clk cell_1375 ( .C (clk), .D (signal_2568), .Q (signal_2569) ) ;
    buf_clk cell_1381 ( .C (clk), .D (signal_2574), .Q (signal_2575) ) ;
    buf_clk cell_1387 ( .C (clk), .D (signal_2580), .Q (signal_2581) ) ;
    buf_clk cell_1393 ( .C (clk), .D (signal_2586), .Q (signal_2587) ) ;
    buf_clk cell_1399 ( .C (clk), .D (signal_2592), .Q (signal_2593) ) ;
    buf_clk cell_1405 ( .C (clk), .D (signal_2598), .Q (signal_2599) ) ;
    buf_clk cell_1411 ( .C (clk), .D (signal_2604), .Q (signal_2605) ) ;
    buf_clk cell_1417 ( .C (clk), .D (signal_2610), .Q (signal_2611) ) ;
    buf_clk cell_1423 ( .C (clk), .D (signal_2616), .Q (signal_2617) ) ;
    buf_clk cell_1429 ( .C (clk), .D (signal_2622), .Q (signal_2623) ) ;
    buf_clk cell_1435 ( .C (clk), .D (signal_2628), .Q (signal_2629) ) ;
    buf_clk cell_1441 ( .C (clk), .D (signal_2634), .Q (signal_2635) ) ;
    buf_clk cell_1447 ( .C (clk), .D (signal_2640), .Q (signal_2641) ) ;
    buf_clk cell_1453 ( .C (clk), .D (signal_2646), .Q (signal_2647) ) ;
    buf_clk cell_1459 ( .C (clk), .D (signal_2652), .Q (signal_2653) ) ;
    buf_clk cell_1465 ( .C (clk), .D (signal_2658), .Q (signal_2659) ) ;
    buf_clk cell_1471 ( .C (clk), .D (signal_2664), .Q (signal_2665) ) ;
    buf_clk cell_1477 ( .C (clk), .D (signal_2670), .Q (signal_2671) ) ;
    buf_clk cell_1483 ( .C (clk), .D (signal_2676), .Q (signal_2677) ) ;
    buf_clk cell_1489 ( .C (clk), .D (signal_2682), .Q (signal_2683) ) ;
    buf_clk cell_1495 ( .C (clk), .D (signal_2688), .Q (signal_2689) ) ;
    buf_clk cell_1501 ( .C (clk), .D (signal_2694), .Q (signal_2695) ) ;
    buf_clk cell_1507 ( .C (clk), .D (signal_2700), .Q (signal_2701) ) ;
    buf_clk cell_1513 ( .C (clk), .D (signal_2706), .Q (signal_2707) ) ;
    buf_clk cell_1519 ( .C (clk), .D (signal_2712), .Q (signal_2713) ) ;
    buf_clk cell_1525 ( .C (clk), .D (signal_2718), .Q (signal_2719) ) ;
    buf_clk cell_1531 ( .C (clk), .D (signal_2724), .Q (signal_2725) ) ;
    buf_clk cell_1537 ( .C (clk), .D (signal_2730), .Q (signal_2731) ) ;
    buf_clk cell_1543 ( .C (clk), .D (signal_2736), .Q (signal_2737) ) ;
    buf_clk cell_1549 ( .C (clk), .D (signal_2742), .Q (signal_2743) ) ;
    buf_clk cell_1555 ( .C (clk), .D (signal_2748), .Q (signal_2749) ) ;
    buf_clk cell_1561 ( .C (clk), .D (signal_2754), .Q (signal_2755) ) ;
    buf_clk cell_1567 ( .C (clk), .D (signal_2760), .Q (signal_2761) ) ;
    buf_clk cell_1573 ( .C (clk), .D (signal_2766), .Q (signal_2767) ) ;
    buf_clk cell_1579 ( .C (clk), .D (signal_2772), .Q (signal_2773) ) ;
    buf_clk cell_1585 ( .C (clk), .D (signal_2778), .Q (signal_2779) ) ;
    buf_clk cell_1591 ( .C (clk), .D (signal_2784), .Q (signal_2785) ) ;
    buf_clk cell_1597 ( .C (clk), .D (signal_2790), .Q (signal_2791) ) ;
    buf_clk cell_1603 ( .C (clk), .D (signal_2796), .Q (signal_2797) ) ;
    buf_clk cell_1609 ( .C (clk), .D (signal_2802), .Q (signal_2803) ) ;
    buf_clk cell_1615 ( .C (clk), .D (signal_2808), .Q (signal_2809) ) ;
    buf_clk cell_1621 ( .C (clk), .D (signal_2814), .Q (signal_2815) ) ;
    buf_clk cell_1627 ( .C (clk), .D (signal_2820), .Q (signal_2821) ) ;
    buf_clk cell_1633 ( .C (clk), .D (signal_2826), .Q (signal_2827) ) ;
    buf_clk cell_1639 ( .C (clk), .D (signal_2832), .Q (signal_2833) ) ;
    buf_clk cell_1645 ( .C (clk), .D (signal_2838), .Q (signal_2839) ) ;
    buf_clk cell_1651 ( .C (clk), .D (signal_2844), .Q (signal_2845) ) ;
    buf_clk cell_1657 ( .C (clk), .D (signal_2850), .Q (signal_2851) ) ;
    buf_clk cell_1663 ( .C (clk), .D (signal_2856), .Q (signal_2857) ) ;
    buf_clk cell_1669 ( .C (clk), .D (signal_2862), .Q (signal_2863) ) ;
    buf_clk cell_1675 ( .C (clk), .D (signal_2868), .Q (signal_2869) ) ;
    buf_clk cell_1681 ( .C (clk), .D (signal_2874), .Q (signal_2875) ) ;
    buf_clk cell_1687 ( .C (clk), .D (signal_2880), .Q (signal_2881) ) ;
    buf_clk cell_1693 ( .C (clk), .D (signal_2886), .Q (signal_2887) ) ;
    buf_clk cell_1699 ( .C (clk), .D (signal_2892), .Q (signal_2893) ) ;
    buf_clk cell_1705 ( .C (clk), .D (signal_2898), .Q (signal_2899) ) ;
    buf_clk cell_1711 ( .C (clk), .D (signal_2904), .Q (signal_2905) ) ;
    buf_clk cell_1717 ( .C (clk), .D (signal_2910), .Q (signal_2911) ) ;
    buf_clk cell_1723 ( .C (clk), .D (signal_2916), .Q (signal_2917) ) ;
    buf_clk cell_1729 ( .C (clk), .D (signal_2922), .Q (signal_2923) ) ;
    buf_clk cell_1735 ( .C (clk), .D (signal_2928), .Q (signal_2929) ) ;
    buf_clk cell_1741 ( .C (clk), .D (signal_2934), .Q (signal_2935) ) ;
    buf_clk cell_1747 ( .C (clk), .D (signal_2940), .Q (signal_2941) ) ;
    buf_clk cell_1753 ( .C (clk), .D (signal_2946), .Q (signal_2947) ) ;
    buf_clk cell_1759 ( .C (clk), .D (signal_2952), .Q (signal_2953) ) ;
    buf_clk cell_1765 ( .C (clk), .D (signal_2958), .Q (signal_2959) ) ;
    buf_clk cell_1771 ( .C (clk), .D (signal_2964), .Q (signal_2965) ) ;
    buf_clk cell_1777 ( .C (clk), .D (signal_2970), .Q (signal_2971) ) ;
    buf_clk cell_1783 ( .C (clk), .D (signal_2976), .Q (signal_2977) ) ;
    buf_clk cell_1789 ( .C (clk), .D (signal_2982), .Q (signal_2983) ) ;
    buf_clk cell_1795 ( .C (clk), .D (signal_2988), .Q (signal_2989) ) ;
    buf_clk cell_1801 ( .C (clk), .D (signal_2994), .Q (signal_2995) ) ;
    buf_clk cell_1807 ( .C (clk), .D (signal_3000), .Q (signal_3001) ) ;
    buf_clk cell_1813 ( .C (clk), .D (signal_3006), .Q (signal_3007) ) ;
    buf_clk cell_1819 ( .C (clk), .D (signal_3012), .Q (signal_3013) ) ;
    buf_clk cell_1825 ( .C (clk), .D (signal_3018), .Q (signal_3019) ) ;
    buf_clk cell_1831 ( .C (clk), .D (signal_3024), .Q (signal_3025) ) ;
    buf_clk cell_1837 ( .C (clk), .D (signal_3030), .Q (signal_3031) ) ;
    buf_clk cell_1843 ( .C (clk), .D (signal_3036), .Q (signal_3037) ) ;
    buf_clk cell_1849 ( .C (clk), .D (signal_3042), .Q (signal_3043) ) ;
    buf_clk cell_1855 ( .C (clk), .D (signal_3048), .Q (signal_3049) ) ;
    buf_clk cell_1861 ( .C (clk), .D (signal_3054), .Q (signal_3055) ) ;
    buf_clk cell_1867 ( .C (clk), .D (signal_3060), .Q (signal_3061) ) ;
    buf_clk cell_1873 ( .C (clk), .D (signal_3066), .Q (signal_3067) ) ;
    buf_clk cell_1879 ( .C (clk), .D (signal_3072), .Q (signal_3073) ) ;
    buf_clk cell_1885 ( .C (clk), .D (signal_3078), .Q (signal_3079) ) ;
    buf_clk cell_1891 ( .C (clk), .D (signal_3084), .Q (signal_3085) ) ;
    buf_clk cell_1897 ( .C (clk), .D (signal_3090), .Q (signal_3091) ) ;
    buf_clk cell_1903 ( .C (clk), .D (signal_3096), .Q (signal_3097) ) ;
    buf_clk cell_1909 ( .C (clk), .D (signal_3102), .Q (signal_3103) ) ;
    buf_clk cell_1915 ( .C (clk), .D (signal_3108), .Q (signal_3109) ) ;
    buf_clk cell_1921 ( .C (clk), .D (signal_3114), .Q (signal_3115) ) ;
    buf_clk cell_1927 ( .C (clk), .D (signal_3120), .Q (signal_3121) ) ;
    buf_clk cell_1933 ( .C (clk), .D (signal_3126), .Q (signal_3127) ) ;
    buf_clk cell_1939 ( .C (clk), .D (signal_3132), .Q (signal_3133) ) ;
    buf_clk cell_1945 ( .C (clk), .D (signal_3138), .Q (signal_3139) ) ;
    buf_clk cell_1955 ( .C (clk), .D (signal_3148), .Q (signal_3149) ) ;
    buf_clk cell_1959 ( .C (clk), .D (signal_3152), .Q (signal_3153) ) ;
    buf_clk cell_1987 ( .C (clk), .D (signal_3180), .Q (signal_3181) ) ;
    buf_clk cell_1991 ( .C (clk), .D (signal_3184), .Q (signal_3185) ) ;
    buf_clk cell_1995 ( .C (clk), .D (signal_3188), .Q (signal_3189) ) ;
    buf_clk cell_1999 ( .C (clk), .D (signal_3192), .Q (signal_3193) ) ;
    buf_clk cell_2011 ( .C (clk), .D (signal_3204), .Q (signal_3205) ) ;
    buf_clk cell_2015 ( .C (clk), .D (signal_3208), .Q (signal_3209) ) ;
    buf_clk cell_2019 ( .C (clk), .D (signal_3212), .Q (signal_3213) ) ;
    buf_clk cell_2023 ( .C (clk), .D (signal_3216), .Q (signal_3217) ) ;
    buf_clk cell_2031 ( .C (clk), .D (signal_3224), .Q (signal_3225) ) ;
    buf_clk cell_2035 ( .C (clk), .D (signal_3228), .Q (signal_3229) ) ;
    buf_clk cell_2039 ( .C (clk), .D (signal_3232), .Q (signal_3233) ) ;
    buf_clk cell_2043 ( .C (clk), .D (signal_3236), .Q (signal_3237) ) ;
    buf_clk cell_2047 ( .C (clk), .D (signal_3240), .Q (signal_3241) ) ;
    buf_clk cell_2051 ( .C (clk), .D (signal_3244), .Q (signal_3245) ) ;
    buf_clk cell_2055 ( .C (clk), .D (signal_3248), .Q (signal_3249) ) ;
    buf_clk cell_2059 ( .C (clk), .D (signal_3252), .Q (signal_3253) ) ;
    buf_clk cell_2063 ( .C (clk), .D (signal_3256), .Q (signal_3257) ) ;
    buf_clk cell_2067 ( .C (clk), .D (signal_3260), .Q (signal_3261) ) ;
    buf_clk cell_2075 ( .C (clk), .D (signal_3268), .Q (signal_3269) ) ;
    buf_clk cell_2079 ( .C (clk), .D (signal_3272), .Q (signal_3273) ) ;
    buf_clk cell_2087 ( .C (clk), .D (signal_3280), .Q (signal_3281) ) ;
    buf_clk cell_2091 ( .C (clk), .D (signal_3284), .Q (signal_3285) ) ;
    buf_clk cell_2099 ( .C (clk), .D (signal_3292), .Q (signal_3293) ) ;
    buf_clk cell_2103 ( .C (clk), .D (signal_3296), .Q (signal_3297) ) ;
    buf_clk cell_2111 ( .C (clk), .D (signal_3304), .Q (signal_3305) ) ;
    buf_clk cell_2115 ( .C (clk), .D (signal_3308), .Q (signal_3309) ) ;
    buf_clk cell_2123 ( .C (clk), .D (signal_3316), .Q (signal_3317) ) ;
    buf_clk cell_2127 ( .C (clk), .D (signal_3320), .Q (signal_3321) ) ;
    buf_clk cell_2135 ( .C (clk), .D (signal_3328), .Q (signal_3329) ) ;
    buf_clk cell_2139 ( .C (clk), .D (signal_3332), .Q (signal_3333) ) ;
    buf_clk cell_2145 ( .C (clk), .D (signal_3338), .Q (signal_3339) ) ;
    buf_clk cell_2153 ( .C (clk), .D (signal_3346), .Q (signal_3347) ) ;
    buf_clk cell_2161 ( .C (clk), .D (signal_3354), .Q (signal_3355) ) ;
    buf_clk cell_2169 ( .C (clk), .D (signal_3362), .Q (signal_3363) ) ;
    buf_clk cell_2177 ( .C (clk), .D (signal_3370), .Q (signal_3371) ) ;
    buf_clk cell_2185 ( .C (clk), .D (signal_3378), .Q (signal_3379) ) ;
    buf_clk cell_2193 ( .C (clk), .D (signal_3386), .Q (signal_3387) ) ;
    buf_clk cell_2201 ( .C (clk), .D (signal_3394), .Q (signal_3395) ) ;
    buf_clk cell_2209 ( .C (clk), .D (signal_3402), .Q (signal_3403) ) ;
    buf_clk cell_2217 ( .C (clk), .D (signal_3410), .Q (signal_3411) ) ;
    buf_clk cell_2225 ( .C (clk), .D (signal_3418), .Q (signal_3419) ) ;
    buf_clk cell_2233 ( .C (clk), .D (signal_3426), .Q (signal_3427) ) ;
    buf_clk cell_2241 ( .C (clk), .D (signal_3434), .Q (signal_3435) ) ;
    buf_clk cell_2249 ( .C (clk), .D (signal_3442), .Q (signal_3443) ) ;
    buf_clk cell_2257 ( .C (clk), .D (signal_3450), .Q (signal_3451) ) ;
    buf_clk cell_2265 ( .C (clk), .D (signal_3458), .Q (signal_3459) ) ;
    buf_clk cell_2273 ( .C (clk), .D (signal_3466), .Q (signal_3467) ) ;
    buf_clk cell_2281 ( .C (clk), .D (signal_3474), .Q (signal_3475) ) ;
    buf_clk cell_2289 ( .C (clk), .D (signal_3482), .Q (signal_3483) ) ;
    buf_clk cell_2297 ( .C (clk), .D (signal_3490), .Q (signal_3491) ) ;
    buf_clk cell_2305 ( .C (clk), .D (signal_3498), .Q (signal_3499) ) ;
    buf_clk cell_2313 ( .C (clk), .D (signal_3506), .Q (signal_3507) ) ;
    buf_clk cell_2321 ( .C (clk), .D (signal_3514), .Q (signal_3515) ) ;
    buf_clk cell_2329 ( .C (clk), .D (signal_3522), .Q (signal_3523) ) ;
    buf_clk cell_2337 ( .C (clk), .D (signal_3530), .Q (signal_3531) ) ;
    buf_clk cell_2345 ( .C (clk), .D (signal_3538), .Q (signal_3539) ) ;
    buf_clk cell_2353 ( .C (clk), .D (signal_3546), .Q (signal_3547) ) ;
    buf_clk cell_2361 ( .C (clk), .D (signal_3554), .Q (signal_3555) ) ;
    buf_clk cell_2369 ( .C (clk), .D (signal_3562), .Q (signal_3563) ) ;
    buf_clk cell_2377 ( .C (clk), .D (signal_3570), .Q (signal_3571) ) ;
    buf_clk cell_2385 ( .C (clk), .D (signal_3578), .Q (signal_3579) ) ;
    buf_clk cell_2393 ( .C (clk), .D (signal_3586), .Q (signal_3587) ) ;
    buf_clk cell_2401 ( .C (clk), .D (signal_3594), .Q (signal_3595) ) ;
    buf_clk cell_2409 ( .C (clk), .D (signal_3602), .Q (signal_3603) ) ;
    buf_clk cell_2417 ( .C (clk), .D (signal_3610), .Q (signal_3611) ) ;
    buf_clk cell_2425 ( .C (clk), .D (signal_3618), .Q (signal_3619) ) ;
    buf_clk cell_2433 ( .C (clk), .D (signal_3626), .Q (signal_3627) ) ;
    buf_clk cell_2441 ( .C (clk), .D (signal_3634), .Q (signal_3635) ) ;
    buf_clk cell_2449 ( .C (clk), .D (signal_3642), .Q (signal_3643) ) ;
    buf_clk cell_2457 ( .C (clk), .D (signal_3650), .Q (signal_3651) ) ;
    buf_clk cell_2465 ( .C (clk), .D (signal_3658), .Q (signal_3659) ) ;
    buf_clk cell_2473 ( .C (clk), .D (signal_3666), .Q (signal_3667) ) ;
    buf_clk cell_2481 ( .C (clk), .D (signal_3674), .Q (signal_3675) ) ;
    buf_clk cell_2489 ( .C (clk), .D (signal_3682), .Q (signal_3683) ) ;
    buf_clk cell_2497 ( .C (clk), .D (signal_3690), .Q (signal_3691) ) ;
    buf_clk cell_2505 ( .C (clk), .D (signal_3698), .Q (signal_3699) ) ;
    buf_clk cell_2513 ( .C (clk), .D (signal_3706), .Q (signal_3707) ) ;
    buf_clk cell_2521 ( .C (clk), .D (signal_3714), .Q (signal_3715) ) ;
    buf_clk cell_2529 ( .C (clk), .D (signal_3722), .Q (signal_3723) ) ;
    buf_clk cell_2537 ( .C (clk), .D (signal_3730), .Q (signal_3731) ) ;
    buf_clk cell_2545 ( .C (clk), .D (signal_3738), .Q (signal_3739) ) ;
    buf_clk cell_2553 ( .C (clk), .D (signal_3746), .Q (signal_3747) ) ;
    buf_clk cell_2561 ( .C (clk), .D (signal_3754), .Q (signal_3755) ) ;
    buf_clk cell_2569 ( .C (clk), .D (signal_3762), .Q (signal_3763) ) ;
    buf_clk cell_2577 ( .C (clk), .D (signal_3770), .Q (signal_3771) ) ;
    buf_clk cell_2585 ( .C (clk), .D (signal_3778), .Q (signal_3779) ) ;
    buf_clk cell_2593 ( .C (clk), .D (signal_3786), .Q (signal_3787) ) ;
    buf_clk cell_2601 ( .C (clk), .D (signal_3794), .Q (signal_3795) ) ;
    buf_clk cell_2609 ( .C (clk), .D (signal_3802), .Q (signal_3803) ) ;
    buf_clk cell_2617 ( .C (clk), .D (signal_3810), .Q (signal_3811) ) ;
    buf_clk cell_2625 ( .C (clk), .D (signal_3818), .Q (signal_3819) ) ;
    buf_clk cell_2633 ( .C (clk), .D (signal_3826), .Q (signal_3827) ) ;
    buf_clk cell_2641 ( .C (clk), .D (signal_3834), .Q (signal_3835) ) ;
    buf_clk cell_2649 ( .C (clk), .D (signal_3842), .Q (signal_3843) ) ;
    buf_clk cell_2657 ( .C (clk), .D (signal_3850), .Q (signal_3851) ) ;
    buf_clk cell_2665 ( .C (clk), .D (signal_3858), .Q (signal_3859) ) ;
    buf_clk cell_2673 ( .C (clk), .D (signal_3866), .Q (signal_3867) ) ;
    buf_clk cell_2681 ( .C (clk), .D (signal_3874), .Q (signal_3875) ) ;
    buf_clk cell_2689 ( .C (clk), .D (signal_3882), .Q (signal_3883) ) ;
    buf_clk cell_2697 ( .C (clk), .D (signal_3890), .Q (signal_3891) ) ;
    buf_clk cell_2705 ( .C (clk), .D (signal_3898), .Q (signal_3899) ) ;
    buf_clk cell_2713 ( .C (clk), .D (signal_3906), .Q (signal_3907) ) ;
    buf_clk cell_2721 ( .C (clk), .D (signal_3914), .Q (signal_3915) ) ;
    buf_clk cell_2729 ( .C (clk), .D (signal_3922), .Q (signal_3923) ) ;
    buf_clk cell_2737 ( .C (clk), .D (signal_3930), .Q (signal_3931) ) ;
    buf_clk cell_2745 ( .C (clk), .D (signal_3938), .Q (signal_3939) ) ;
    buf_clk cell_2753 ( .C (clk), .D (signal_3946), .Q (signal_3947) ) ;
    buf_clk cell_2761 ( .C (clk), .D (signal_3954), .Q (signal_3955) ) ;
    buf_clk cell_2769 ( .C (clk), .D (signal_3962), .Q (signal_3963) ) ;
    buf_clk cell_2777 ( .C (clk), .D (signal_3970), .Q (signal_3971) ) ;
    buf_clk cell_2785 ( .C (clk), .D (signal_3978), .Q (signal_3979) ) ;
    buf_clk cell_2793 ( .C (clk), .D (signal_3986), .Q (signal_3987) ) ;
    buf_clk cell_2801 ( .C (clk), .D (signal_3994), .Q (signal_3995) ) ;
    buf_clk cell_2809 ( .C (clk), .D (signal_4002), .Q (signal_4003) ) ;
    buf_clk cell_2817 ( .C (clk), .D (signal_4010), .Q (signal_4011) ) ;
    buf_clk cell_2825 ( .C (clk), .D (signal_4018), .Q (signal_4019) ) ;
    buf_clk cell_2833 ( .C (clk), .D (signal_4026), .Q (signal_4027) ) ;
    buf_clk cell_2841 ( .C (clk), .D (signal_4034), .Q (signal_4035) ) ;
    buf_clk cell_2849 ( .C (clk), .D (signal_4042), .Q (signal_4043) ) ;
    buf_clk cell_2857 ( .C (clk), .D (signal_4050), .Q (signal_4051) ) ;
    buf_clk cell_2865 ( .C (clk), .D (signal_4058), .Q (signal_4059) ) ;
    buf_clk cell_2873 ( .C (clk), .D (signal_4066), .Q (signal_4067) ) ;
    buf_clk cell_2881 ( .C (clk), .D (signal_4074), .Q (signal_4075) ) ;
    buf_clk cell_2889 ( .C (clk), .D (signal_4082), .Q (signal_4083) ) ;
    buf_clk cell_2897 ( .C (clk), .D (signal_4090), .Q (signal_4091) ) ;
    buf_clk cell_2905 ( .C (clk), .D (signal_4098), .Q (signal_4099) ) ;
    buf_clk cell_2913 ( .C (clk), .D (signal_4106), .Q (signal_4107) ) ;
    buf_clk cell_2921 ( .C (clk), .D (signal_4114), .Q (signal_4115) ) ;
    buf_clk cell_2929 ( .C (clk), .D (signal_4122), .Q (signal_4123) ) ;
    buf_clk cell_2937 ( .C (clk), .D (signal_4130), .Q (signal_4131) ) ;
    buf_clk cell_2945 ( .C (clk), .D (signal_4138), .Q (signal_4139) ) ;
    buf_clk cell_2953 ( .C (clk), .D (signal_4146), .Q (signal_4147) ) ;
    buf_clk cell_2961 ( .C (clk), .D (signal_4154), .Q (signal_4155) ) ;
    buf_clk cell_2969 ( .C (clk), .D (signal_4162), .Q (signal_4163) ) ;
    buf_clk cell_2977 ( .C (clk), .D (signal_4170), .Q (signal_4171) ) ;
    buf_clk cell_2985 ( .C (clk), .D (signal_4178), .Q (signal_4179) ) ;
    buf_clk cell_2993 ( .C (clk), .D (signal_4186), .Q (signal_4187) ) ;
    buf_clk cell_3001 ( .C (clk), .D (signal_4194), .Q (signal_4195) ) ;
    buf_clk cell_3009 ( .C (clk), .D (signal_4202), .Q (signal_4203) ) ;
    buf_clk cell_3017 ( .C (clk), .D (signal_4210), .Q (signal_4211) ) ;
    buf_clk cell_3025 ( .C (clk), .D (signal_4218), .Q (signal_4219) ) ;
    buf_clk cell_3033 ( .C (clk), .D (signal_4226), .Q (signal_4227) ) ;
    buf_clk cell_3041 ( .C (clk), .D (signal_4234), .Q (signal_4235) ) ;
    buf_clk cell_3049 ( .C (clk), .D (signal_4242), .Q (signal_4243) ) ;
    buf_clk cell_3057 ( .C (clk), .D (signal_4250), .Q (signal_4251) ) ;
    buf_clk cell_3065 ( .C (clk), .D (signal_4258), .Q (signal_4259) ) ;
    buf_clk cell_3073 ( .C (clk), .D (signal_4266), .Q (signal_4267) ) ;
    buf_clk cell_3081 ( .C (clk), .D (signal_4274), .Q (signal_4275) ) ;
    buf_clk cell_3089 ( .C (clk), .D (signal_4282), .Q (signal_4283) ) ;
    buf_clk cell_3097 ( .C (clk), .D (signal_4290), .Q (signal_4291) ) ;
    buf_clk cell_3105 ( .C (clk), .D (signal_4298), .Q (signal_4299) ) ;
    buf_clk cell_3113 ( .C (clk), .D (signal_4306), .Q (signal_4307) ) ;
    buf_clk cell_3121 ( .C (clk), .D (signal_4314), .Q (signal_4315) ) ;
    buf_clk cell_3129 ( .C (clk), .D (signal_4322), .Q (signal_4323) ) ;
    buf_clk cell_3137 ( .C (clk), .D (signal_4330), .Q (signal_4331) ) ;
    buf_clk cell_3145 ( .C (clk), .D (signal_4338), .Q (signal_4339) ) ;
    buf_clk cell_3153 ( .C (clk), .D (signal_4346), .Q (signal_4347) ) ;
    buf_clk cell_3161 ( .C (clk), .D (signal_4354), .Q (signal_4355) ) ;
    buf_clk cell_3489 ( .C (clk), .D (signal_4682), .Q (signal_4683) ) ;
    buf_clk cell_3497 ( .C (clk), .D (signal_4690), .Q (signal_4691) ) ;
    buf_clk cell_3505 ( .C (clk), .D (signal_4698), .Q (signal_4699) ) ;
    buf_clk cell_3513 ( .C (clk), .D (signal_4706), .Q (signal_4707) ) ;
    buf_clk cell_3521 ( .C (clk), .D (signal_4714), .Q (signal_4715) ) ;
    buf_clk cell_3529 ( .C (clk), .D (signal_4722), .Q (signal_4723) ) ;
    buf_clk cell_3537 ( .C (clk), .D (signal_4730), .Q (signal_4731) ) ;
    buf_clk cell_3545 ( .C (clk), .D (signal_4738), .Q (signal_4739) ) ;
    buf_clk cell_3553 ( .C (clk), .D (signal_4746), .Q (signal_4747) ) ;
    buf_clk cell_3561 ( .C (clk), .D (signal_4754), .Q (signal_4755) ) ;

    /* cells in depth 3 */
    buf_clk cell_1178 ( .C (clk), .D (signal_2371), .Q (signal_2372) ) ;
    buf_clk cell_1184 ( .C (clk), .D (signal_2377), .Q (signal_2378) ) ;
    buf_clk cell_1190 ( .C (clk), .D (signal_2383), .Q (signal_2384) ) ;
    buf_clk cell_1196 ( .C (clk), .D (signal_2389), .Q (signal_2390) ) ;
    buf_clk cell_1202 ( .C (clk), .D (signal_2395), .Q (signal_2396) ) ;
    buf_clk cell_1208 ( .C (clk), .D (signal_2401), .Q (signal_2402) ) ;
    buf_clk cell_1214 ( .C (clk), .D (signal_2407), .Q (signal_2408) ) ;
    buf_clk cell_1220 ( .C (clk), .D (signal_2413), .Q (signal_2414) ) ;
    buf_clk cell_1226 ( .C (clk), .D (signal_2419), .Q (signal_2420) ) ;
    buf_clk cell_1232 ( .C (clk), .D (signal_2425), .Q (signal_2426) ) ;
    buf_clk cell_1238 ( .C (clk), .D (signal_2431), .Q (signal_2432) ) ;
    buf_clk cell_1244 ( .C (clk), .D (signal_2437), .Q (signal_2438) ) ;
    buf_clk cell_1250 ( .C (clk), .D (signal_2443), .Q (signal_2444) ) ;
    buf_clk cell_1256 ( .C (clk), .D (signal_2449), .Q (signal_2450) ) ;
    buf_clk cell_1262 ( .C (clk), .D (signal_2455), .Q (signal_2456) ) ;
    buf_clk cell_1268 ( .C (clk), .D (signal_2461), .Q (signal_2462) ) ;
    buf_clk cell_1274 ( .C (clk), .D (signal_2467), .Q (signal_2468) ) ;
    buf_clk cell_1280 ( .C (clk), .D (signal_2473), .Q (signal_2474) ) ;
    buf_clk cell_1286 ( .C (clk), .D (signal_2479), .Q (signal_2480) ) ;
    buf_clk cell_1292 ( .C (clk), .D (signal_2485), .Q (signal_2486) ) ;
    buf_clk cell_1298 ( .C (clk), .D (signal_2491), .Q (signal_2492) ) ;
    buf_clk cell_1304 ( .C (clk), .D (signal_2497), .Q (signal_2498) ) ;
    buf_clk cell_1310 ( .C (clk), .D (signal_2503), .Q (signal_2504) ) ;
    buf_clk cell_1316 ( .C (clk), .D (signal_2509), .Q (signal_2510) ) ;
    buf_clk cell_1322 ( .C (clk), .D (signal_2515), .Q (signal_2516) ) ;
    buf_clk cell_1328 ( .C (clk), .D (signal_2521), .Q (signal_2522) ) ;
    buf_clk cell_1334 ( .C (clk), .D (signal_2527), .Q (signal_2528) ) ;
    buf_clk cell_1340 ( .C (clk), .D (signal_2533), .Q (signal_2534) ) ;
    buf_clk cell_1346 ( .C (clk), .D (signal_2539), .Q (signal_2540) ) ;
    buf_clk cell_1352 ( .C (clk), .D (signal_2545), .Q (signal_2546) ) ;
    buf_clk cell_1358 ( .C (clk), .D (signal_2551), .Q (signal_2552) ) ;
    buf_clk cell_1364 ( .C (clk), .D (signal_2557), .Q (signal_2558) ) ;
    buf_clk cell_1370 ( .C (clk), .D (signal_2563), .Q (signal_2564) ) ;
    buf_clk cell_1376 ( .C (clk), .D (signal_2569), .Q (signal_2570) ) ;
    buf_clk cell_1382 ( .C (clk), .D (signal_2575), .Q (signal_2576) ) ;
    buf_clk cell_1388 ( .C (clk), .D (signal_2581), .Q (signal_2582) ) ;
    buf_clk cell_1394 ( .C (clk), .D (signal_2587), .Q (signal_2588) ) ;
    buf_clk cell_1400 ( .C (clk), .D (signal_2593), .Q (signal_2594) ) ;
    buf_clk cell_1406 ( .C (clk), .D (signal_2599), .Q (signal_2600) ) ;
    buf_clk cell_1412 ( .C (clk), .D (signal_2605), .Q (signal_2606) ) ;
    buf_clk cell_1418 ( .C (clk), .D (signal_2611), .Q (signal_2612) ) ;
    buf_clk cell_1424 ( .C (clk), .D (signal_2617), .Q (signal_2618) ) ;
    buf_clk cell_1430 ( .C (clk), .D (signal_2623), .Q (signal_2624) ) ;
    buf_clk cell_1436 ( .C (clk), .D (signal_2629), .Q (signal_2630) ) ;
    buf_clk cell_1442 ( .C (clk), .D (signal_2635), .Q (signal_2636) ) ;
    buf_clk cell_1448 ( .C (clk), .D (signal_2641), .Q (signal_2642) ) ;
    buf_clk cell_1454 ( .C (clk), .D (signal_2647), .Q (signal_2648) ) ;
    buf_clk cell_1460 ( .C (clk), .D (signal_2653), .Q (signal_2654) ) ;
    buf_clk cell_1466 ( .C (clk), .D (signal_2659), .Q (signal_2660) ) ;
    buf_clk cell_1472 ( .C (clk), .D (signal_2665), .Q (signal_2666) ) ;
    buf_clk cell_1478 ( .C (clk), .D (signal_2671), .Q (signal_2672) ) ;
    buf_clk cell_1484 ( .C (clk), .D (signal_2677), .Q (signal_2678) ) ;
    buf_clk cell_1490 ( .C (clk), .D (signal_2683), .Q (signal_2684) ) ;
    buf_clk cell_1496 ( .C (clk), .D (signal_2689), .Q (signal_2690) ) ;
    buf_clk cell_1502 ( .C (clk), .D (signal_2695), .Q (signal_2696) ) ;
    buf_clk cell_1508 ( .C (clk), .D (signal_2701), .Q (signal_2702) ) ;
    buf_clk cell_1514 ( .C (clk), .D (signal_2707), .Q (signal_2708) ) ;
    buf_clk cell_1520 ( .C (clk), .D (signal_2713), .Q (signal_2714) ) ;
    buf_clk cell_1526 ( .C (clk), .D (signal_2719), .Q (signal_2720) ) ;
    buf_clk cell_1532 ( .C (clk), .D (signal_2725), .Q (signal_2726) ) ;
    buf_clk cell_1538 ( .C (clk), .D (signal_2731), .Q (signal_2732) ) ;
    buf_clk cell_1544 ( .C (clk), .D (signal_2737), .Q (signal_2738) ) ;
    buf_clk cell_1550 ( .C (clk), .D (signal_2743), .Q (signal_2744) ) ;
    buf_clk cell_1556 ( .C (clk), .D (signal_2749), .Q (signal_2750) ) ;
    buf_clk cell_1562 ( .C (clk), .D (signal_2755), .Q (signal_2756) ) ;
    buf_clk cell_1568 ( .C (clk), .D (signal_2761), .Q (signal_2762) ) ;
    buf_clk cell_1574 ( .C (clk), .D (signal_2767), .Q (signal_2768) ) ;
    buf_clk cell_1580 ( .C (clk), .D (signal_2773), .Q (signal_2774) ) ;
    buf_clk cell_1586 ( .C (clk), .D (signal_2779), .Q (signal_2780) ) ;
    buf_clk cell_1592 ( .C (clk), .D (signal_2785), .Q (signal_2786) ) ;
    buf_clk cell_1598 ( .C (clk), .D (signal_2791), .Q (signal_2792) ) ;
    buf_clk cell_1604 ( .C (clk), .D (signal_2797), .Q (signal_2798) ) ;
    buf_clk cell_1610 ( .C (clk), .D (signal_2803), .Q (signal_2804) ) ;
    buf_clk cell_1616 ( .C (clk), .D (signal_2809), .Q (signal_2810) ) ;
    buf_clk cell_1622 ( .C (clk), .D (signal_2815), .Q (signal_2816) ) ;
    buf_clk cell_1628 ( .C (clk), .D (signal_2821), .Q (signal_2822) ) ;
    buf_clk cell_1634 ( .C (clk), .D (signal_2827), .Q (signal_2828) ) ;
    buf_clk cell_1640 ( .C (clk), .D (signal_2833), .Q (signal_2834) ) ;
    buf_clk cell_1646 ( .C (clk), .D (signal_2839), .Q (signal_2840) ) ;
    buf_clk cell_1652 ( .C (clk), .D (signal_2845), .Q (signal_2846) ) ;
    buf_clk cell_1658 ( .C (clk), .D (signal_2851), .Q (signal_2852) ) ;
    buf_clk cell_1664 ( .C (clk), .D (signal_2857), .Q (signal_2858) ) ;
    buf_clk cell_1670 ( .C (clk), .D (signal_2863), .Q (signal_2864) ) ;
    buf_clk cell_1676 ( .C (clk), .D (signal_2869), .Q (signal_2870) ) ;
    buf_clk cell_1682 ( .C (clk), .D (signal_2875), .Q (signal_2876) ) ;
    buf_clk cell_1688 ( .C (clk), .D (signal_2881), .Q (signal_2882) ) ;
    buf_clk cell_1694 ( .C (clk), .D (signal_2887), .Q (signal_2888) ) ;
    buf_clk cell_1700 ( .C (clk), .D (signal_2893), .Q (signal_2894) ) ;
    buf_clk cell_1706 ( .C (clk), .D (signal_2899), .Q (signal_2900) ) ;
    buf_clk cell_1712 ( .C (clk), .D (signal_2905), .Q (signal_2906) ) ;
    buf_clk cell_1718 ( .C (clk), .D (signal_2911), .Q (signal_2912) ) ;
    buf_clk cell_1724 ( .C (clk), .D (signal_2917), .Q (signal_2918) ) ;
    buf_clk cell_1730 ( .C (clk), .D (signal_2923), .Q (signal_2924) ) ;
    buf_clk cell_1736 ( .C (clk), .D (signal_2929), .Q (signal_2930) ) ;
    buf_clk cell_1742 ( .C (clk), .D (signal_2935), .Q (signal_2936) ) ;
    buf_clk cell_1748 ( .C (clk), .D (signal_2941), .Q (signal_2942) ) ;
    buf_clk cell_1754 ( .C (clk), .D (signal_2947), .Q (signal_2948) ) ;
    buf_clk cell_1760 ( .C (clk), .D (signal_2953), .Q (signal_2954) ) ;
    buf_clk cell_1766 ( .C (clk), .D (signal_2959), .Q (signal_2960) ) ;
    buf_clk cell_1772 ( .C (clk), .D (signal_2965), .Q (signal_2966) ) ;
    buf_clk cell_1778 ( .C (clk), .D (signal_2971), .Q (signal_2972) ) ;
    buf_clk cell_1784 ( .C (clk), .D (signal_2977), .Q (signal_2978) ) ;
    buf_clk cell_1790 ( .C (clk), .D (signal_2983), .Q (signal_2984) ) ;
    buf_clk cell_1796 ( .C (clk), .D (signal_2989), .Q (signal_2990) ) ;
    buf_clk cell_1802 ( .C (clk), .D (signal_2995), .Q (signal_2996) ) ;
    buf_clk cell_1808 ( .C (clk), .D (signal_3001), .Q (signal_3002) ) ;
    buf_clk cell_1814 ( .C (clk), .D (signal_3007), .Q (signal_3008) ) ;
    buf_clk cell_1820 ( .C (clk), .D (signal_3013), .Q (signal_3014) ) ;
    buf_clk cell_1826 ( .C (clk), .D (signal_3019), .Q (signal_3020) ) ;
    buf_clk cell_1832 ( .C (clk), .D (signal_3025), .Q (signal_3026) ) ;
    buf_clk cell_1838 ( .C (clk), .D (signal_3031), .Q (signal_3032) ) ;
    buf_clk cell_1844 ( .C (clk), .D (signal_3037), .Q (signal_3038) ) ;
    buf_clk cell_1850 ( .C (clk), .D (signal_3043), .Q (signal_3044) ) ;
    buf_clk cell_1856 ( .C (clk), .D (signal_3049), .Q (signal_3050) ) ;
    buf_clk cell_1862 ( .C (clk), .D (signal_3055), .Q (signal_3056) ) ;
    buf_clk cell_1868 ( .C (clk), .D (signal_3061), .Q (signal_3062) ) ;
    buf_clk cell_1874 ( .C (clk), .D (signal_3067), .Q (signal_3068) ) ;
    buf_clk cell_1880 ( .C (clk), .D (signal_3073), .Q (signal_3074) ) ;
    buf_clk cell_1886 ( .C (clk), .D (signal_3079), .Q (signal_3080) ) ;
    buf_clk cell_1892 ( .C (clk), .D (signal_3085), .Q (signal_3086) ) ;
    buf_clk cell_1898 ( .C (clk), .D (signal_3091), .Q (signal_3092) ) ;
    buf_clk cell_1904 ( .C (clk), .D (signal_3097), .Q (signal_3098) ) ;
    buf_clk cell_1910 ( .C (clk), .D (signal_3103), .Q (signal_3104) ) ;
    buf_clk cell_1916 ( .C (clk), .D (signal_3109), .Q (signal_3110) ) ;
    buf_clk cell_1922 ( .C (clk), .D (signal_3115), .Q (signal_3116) ) ;
    buf_clk cell_1928 ( .C (clk), .D (signal_3121), .Q (signal_3122) ) ;
    buf_clk cell_1934 ( .C (clk), .D (signal_3127), .Q (signal_3128) ) ;
    buf_clk cell_1940 ( .C (clk), .D (signal_3133), .Q (signal_3134) ) ;
    buf_clk cell_1946 ( .C (clk), .D (signal_3139), .Q (signal_3140) ) ;
    buf_clk cell_1950 ( .C (clk), .D (signal_2315), .Q (signal_3144) ) ;
    buf_clk cell_1952 ( .C (clk), .D (signal_2317), .Q (signal_3146) ) ;
    buf_clk cell_1956 ( .C (clk), .D (signal_3149), .Q (signal_3150) ) ;
    buf_clk cell_1960 ( .C (clk), .D (signal_3153), .Q (signal_3154) ) ;
    buf_clk cell_1962 ( .C (clk), .D (signal_2307), .Q (signal_3156) ) ;
    buf_clk cell_1964 ( .C (clk), .D (signal_2309), .Q (signal_3158) ) ;
    buf_clk cell_1966 ( .C (clk), .D (signal_2259), .Q (signal_3160) ) ;
    buf_clk cell_1968 ( .C (clk), .D (signal_2261), .Q (signal_3162) ) ;
    buf_clk cell_1970 ( .C (clk), .D (signal_2255), .Q (signal_3164) ) ;
    buf_clk cell_1972 ( .C (clk), .D (signal_2257), .Q (signal_3166) ) ;
    buf_clk cell_1974 ( .C (clk), .D (signal_2303), .Q (signal_3168) ) ;
    buf_clk cell_1976 ( .C (clk), .D (signal_2305), .Q (signal_3170) ) ;
    buf_clk cell_1978 ( .C (clk), .D (signal_2271), .Q (signal_3172) ) ;
    buf_clk cell_1980 ( .C (clk), .D (signal_2273), .Q (signal_3174) ) ;
    buf_clk cell_1982 ( .C (clk), .D (signal_2251), .Q (signal_3176) ) ;
    buf_clk cell_1984 ( .C (clk), .D (signal_2253), .Q (signal_3178) ) ;
    buf_clk cell_1988 ( .C (clk), .D (signal_3181), .Q (signal_3182) ) ;
    buf_clk cell_1992 ( .C (clk), .D (signal_3185), .Q (signal_3186) ) ;
    buf_clk cell_1996 ( .C (clk), .D (signal_3189), .Q (signal_3190) ) ;
    buf_clk cell_2000 ( .C (clk), .D (signal_3193), .Q (signal_3194) ) ;
    buf_clk cell_2002 ( .C (clk), .D (signal_2319), .Q (signal_3196) ) ;
    buf_clk cell_2004 ( .C (clk), .D (signal_2321), .Q (signal_3198) ) ;
    buf_clk cell_2006 ( .C (clk), .D (signal_2311), .Q (signal_3200) ) ;
    buf_clk cell_2008 ( .C (clk), .D (signal_2313), .Q (signal_3202) ) ;
    buf_clk cell_2012 ( .C (clk), .D (signal_3205), .Q (signal_3206) ) ;
    buf_clk cell_2016 ( .C (clk), .D (signal_3209), .Q (signal_3210) ) ;
    buf_clk cell_2020 ( .C (clk), .D (signal_3213), .Q (signal_3214) ) ;
    buf_clk cell_2024 ( .C (clk), .D (signal_3217), .Q (signal_3218) ) ;
    buf_clk cell_2026 ( .C (clk), .D (signal_2279), .Q (signal_3220) ) ;
    buf_clk cell_2028 ( .C (clk), .D (signal_2281), .Q (signal_3222) ) ;
    buf_clk cell_2032 ( .C (clk), .D (signal_3225), .Q (signal_3226) ) ;
    buf_clk cell_2036 ( .C (clk), .D (signal_3229), .Q (signal_3230) ) ;
    buf_clk cell_2040 ( .C (clk), .D (signal_3233), .Q (signal_3234) ) ;
    buf_clk cell_2044 ( .C (clk), .D (signal_3237), .Q (signal_3238) ) ;
    buf_clk cell_2048 ( .C (clk), .D (signal_3241), .Q (signal_3242) ) ;
    buf_clk cell_2052 ( .C (clk), .D (signal_3245), .Q (signal_3246) ) ;
    buf_clk cell_2056 ( .C (clk), .D (signal_3249), .Q (signal_3250) ) ;
    buf_clk cell_2060 ( .C (clk), .D (signal_3253), .Q (signal_3254) ) ;
    buf_clk cell_2064 ( .C (clk), .D (signal_3257), .Q (signal_3258) ) ;
    buf_clk cell_2068 ( .C (clk), .D (signal_3261), .Q (signal_3262) ) ;
    buf_clk cell_2070 ( .C (clk), .D (signal_2327), .Q (signal_3264) ) ;
    buf_clk cell_2072 ( .C (clk), .D (signal_2329), .Q (signal_3266) ) ;
    buf_clk cell_2076 ( .C (clk), .D (signal_3269), .Q (signal_3270) ) ;
    buf_clk cell_2080 ( .C (clk), .D (signal_3273), .Q (signal_3274) ) ;
    buf_clk cell_2082 ( .C (clk), .D (signal_2335), .Q (signal_3276) ) ;
    buf_clk cell_2084 ( .C (clk), .D (signal_2337), .Q (signal_3278) ) ;
    buf_clk cell_2088 ( .C (clk), .D (signal_3281), .Q (signal_3282) ) ;
    buf_clk cell_2092 ( .C (clk), .D (signal_3285), .Q (signal_3286) ) ;
    buf_clk cell_2094 ( .C (clk), .D (signal_2343), .Q (signal_3288) ) ;
    buf_clk cell_2096 ( .C (clk), .D (signal_2345), .Q (signal_3290) ) ;
    buf_clk cell_2100 ( .C (clk), .D (signal_3293), .Q (signal_3294) ) ;
    buf_clk cell_2104 ( .C (clk), .D (signal_3297), .Q (signal_3298) ) ;
    buf_clk cell_2106 ( .C (clk), .D (signal_2351), .Q (signal_3300) ) ;
    buf_clk cell_2108 ( .C (clk), .D (signal_2353), .Q (signal_3302) ) ;
    buf_clk cell_2112 ( .C (clk), .D (signal_3305), .Q (signal_3306) ) ;
    buf_clk cell_2116 ( .C (clk), .D (signal_3309), .Q (signal_3310) ) ;
    buf_clk cell_2118 ( .C (clk), .D (signal_2359), .Q (signal_3312) ) ;
    buf_clk cell_2120 ( .C (clk), .D (signal_2361), .Q (signal_3314) ) ;
    buf_clk cell_2124 ( .C (clk), .D (signal_3317), .Q (signal_3318) ) ;
    buf_clk cell_2128 ( .C (clk), .D (signal_3321), .Q (signal_3322) ) ;
    buf_clk cell_2130 ( .C (clk), .D (signal_2367), .Q (signal_3324) ) ;
    buf_clk cell_2132 ( .C (clk), .D (signal_2369), .Q (signal_3326) ) ;
    buf_clk cell_2136 ( .C (clk), .D (signal_3329), .Q (signal_3330) ) ;
    buf_clk cell_2140 ( .C (clk), .D (signal_3333), .Q (signal_3334) ) ;
    buf_clk cell_2146 ( .C (clk), .D (signal_3339), .Q (signal_3340) ) ;
    buf_clk cell_2154 ( .C (clk), .D (signal_3347), .Q (signal_3348) ) ;
    buf_clk cell_2162 ( .C (clk), .D (signal_3355), .Q (signal_3356) ) ;
    buf_clk cell_2170 ( .C (clk), .D (signal_3363), .Q (signal_3364) ) ;
    buf_clk cell_2178 ( .C (clk), .D (signal_3371), .Q (signal_3372) ) ;
    buf_clk cell_2186 ( .C (clk), .D (signal_3379), .Q (signal_3380) ) ;
    buf_clk cell_2194 ( .C (clk), .D (signal_3387), .Q (signal_3388) ) ;
    buf_clk cell_2202 ( .C (clk), .D (signal_3395), .Q (signal_3396) ) ;
    buf_clk cell_2210 ( .C (clk), .D (signal_3403), .Q (signal_3404) ) ;
    buf_clk cell_2218 ( .C (clk), .D (signal_3411), .Q (signal_3412) ) ;
    buf_clk cell_2226 ( .C (clk), .D (signal_3419), .Q (signal_3420) ) ;
    buf_clk cell_2234 ( .C (clk), .D (signal_3427), .Q (signal_3428) ) ;
    buf_clk cell_2242 ( .C (clk), .D (signal_3435), .Q (signal_3436) ) ;
    buf_clk cell_2250 ( .C (clk), .D (signal_3443), .Q (signal_3444) ) ;
    buf_clk cell_2258 ( .C (clk), .D (signal_3451), .Q (signal_3452) ) ;
    buf_clk cell_2266 ( .C (clk), .D (signal_3459), .Q (signal_3460) ) ;
    buf_clk cell_2274 ( .C (clk), .D (signal_3467), .Q (signal_3468) ) ;
    buf_clk cell_2282 ( .C (clk), .D (signal_3475), .Q (signal_3476) ) ;
    buf_clk cell_2290 ( .C (clk), .D (signal_3483), .Q (signal_3484) ) ;
    buf_clk cell_2298 ( .C (clk), .D (signal_3491), .Q (signal_3492) ) ;
    buf_clk cell_2306 ( .C (clk), .D (signal_3499), .Q (signal_3500) ) ;
    buf_clk cell_2314 ( .C (clk), .D (signal_3507), .Q (signal_3508) ) ;
    buf_clk cell_2322 ( .C (clk), .D (signal_3515), .Q (signal_3516) ) ;
    buf_clk cell_2330 ( .C (clk), .D (signal_3523), .Q (signal_3524) ) ;
    buf_clk cell_2338 ( .C (clk), .D (signal_3531), .Q (signal_3532) ) ;
    buf_clk cell_2346 ( .C (clk), .D (signal_3539), .Q (signal_3540) ) ;
    buf_clk cell_2354 ( .C (clk), .D (signal_3547), .Q (signal_3548) ) ;
    buf_clk cell_2362 ( .C (clk), .D (signal_3555), .Q (signal_3556) ) ;
    buf_clk cell_2370 ( .C (clk), .D (signal_3563), .Q (signal_3564) ) ;
    buf_clk cell_2378 ( .C (clk), .D (signal_3571), .Q (signal_3572) ) ;
    buf_clk cell_2386 ( .C (clk), .D (signal_3579), .Q (signal_3580) ) ;
    buf_clk cell_2394 ( .C (clk), .D (signal_3587), .Q (signal_3588) ) ;
    buf_clk cell_2402 ( .C (clk), .D (signal_3595), .Q (signal_3596) ) ;
    buf_clk cell_2410 ( .C (clk), .D (signal_3603), .Q (signal_3604) ) ;
    buf_clk cell_2418 ( .C (clk), .D (signal_3611), .Q (signal_3612) ) ;
    buf_clk cell_2426 ( .C (clk), .D (signal_3619), .Q (signal_3620) ) ;
    buf_clk cell_2434 ( .C (clk), .D (signal_3627), .Q (signal_3628) ) ;
    buf_clk cell_2442 ( .C (clk), .D (signal_3635), .Q (signal_3636) ) ;
    buf_clk cell_2450 ( .C (clk), .D (signal_3643), .Q (signal_3644) ) ;
    buf_clk cell_2458 ( .C (clk), .D (signal_3651), .Q (signal_3652) ) ;
    buf_clk cell_2466 ( .C (clk), .D (signal_3659), .Q (signal_3660) ) ;
    buf_clk cell_2474 ( .C (clk), .D (signal_3667), .Q (signal_3668) ) ;
    buf_clk cell_2482 ( .C (clk), .D (signal_3675), .Q (signal_3676) ) ;
    buf_clk cell_2490 ( .C (clk), .D (signal_3683), .Q (signal_3684) ) ;
    buf_clk cell_2498 ( .C (clk), .D (signal_3691), .Q (signal_3692) ) ;
    buf_clk cell_2506 ( .C (clk), .D (signal_3699), .Q (signal_3700) ) ;
    buf_clk cell_2514 ( .C (clk), .D (signal_3707), .Q (signal_3708) ) ;
    buf_clk cell_2522 ( .C (clk), .D (signal_3715), .Q (signal_3716) ) ;
    buf_clk cell_2530 ( .C (clk), .D (signal_3723), .Q (signal_3724) ) ;
    buf_clk cell_2538 ( .C (clk), .D (signal_3731), .Q (signal_3732) ) ;
    buf_clk cell_2546 ( .C (clk), .D (signal_3739), .Q (signal_3740) ) ;
    buf_clk cell_2554 ( .C (clk), .D (signal_3747), .Q (signal_3748) ) ;
    buf_clk cell_2562 ( .C (clk), .D (signal_3755), .Q (signal_3756) ) ;
    buf_clk cell_2570 ( .C (clk), .D (signal_3763), .Q (signal_3764) ) ;
    buf_clk cell_2578 ( .C (clk), .D (signal_3771), .Q (signal_3772) ) ;
    buf_clk cell_2586 ( .C (clk), .D (signal_3779), .Q (signal_3780) ) ;
    buf_clk cell_2594 ( .C (clk), .D (signal_3787), .Q (signal_3788) ) ;
    buf_clk cell_2602 ( .C (clk), .D (signal_3795), .Q (signal_3796) ) ;
    buf_clk cell_2610 ( .C (clk), .D (signal_3803), .Q (signal_3804) ) ;
    buf_clk cell_2618 ( .C (clk), .D (signal_3811), .Q (signal_3812) ) ;
    buf_clk cell_2626 ( .C (clk), .D (signal_3819), .Q (signal_3820) ) ;
    buf_clk cell_2634 ( .C (clk), .D (signal_3827), .Q (signal_3828) ) ;
    buf_clk cell_2642 ( .C (clk), .D (signal_3835), .Q (signal_3836) ) ;
    buf_clk cell_2650 ( .C (clk), .D (signal_3843), .Q (signal_3844) ) ;
    buf_clk cell_2658 ( .C (clk), .D (signal_3851), .Q (signal_3852) ) ;
    buf_clk cell_2666 ( .C (clk), .D (signal_3859), .Q (signal_3860) ) ;
    buf_clk cell_2674 ( .C (clk), .D (signal_3867), .Q (signal_3868) ) ;
    buf_clk cell_2682 ( .C (clk), .D (signal_3875), .Q (signal_3876) ) ;
    buf_clk cell_2690 ( .C (clk), .D (signal_3883), .Q (signal_3884) ) ;
    buf_clk cell_2698 ( .C (clk), .D (signal_3891), .Q (signal_3892) ) ;
    buf_clk cell_2706 ( .C (clk), .D (signal_3899), .Q (signal_3900) ) ;
    buf_clk cell_2714 ( .C (clk), .D (signal_3907), .Q (signal_3908) ) ;
    buf_clk cell_2722 ( .C (clk), .D (signal_3915), .Q (signal_3916) ) ;
    buf_clk cell_2730 ( .C (clk), .D (signal_3923), .Q (signal_3924) ) ;
    buf_clk cell_2738 ( .C (clk), .D (signal_3931), .Q (signal_3932) ) ;
    buf_clk cell_2746 ( .C (clk), .D (signal_3939), .Q (signal_3940) ) ;
    buf_clk cell_2754 ( .C (clk), .D (signal_3947), .Q (signal_3948) ) ;
    buf_clk cell_2762 ( .C (clk), .D (signal_3955), .Q (signal_3956) ) ;
    buf_clk cell_2770 ( .C (clk), .D (signal_3963), .Q (signal_3964) ) ;
    buf_clk cell_2778 ( .C (clk), .D (signal_3971), .Q (signal_3972) ) ;
    buf_clk cell_2786 ( .C (clk), .D (signal_3979), .Q (signal_3980) ) ;
    buf_clk cell_2794 ( .C (clk), .D (signal_3987), .Q (signal_3988) ) ;
    buf_clk cell_2802 ( .C (clk), .D (signal_3995), .Q (signal_3996) ) ;
    buf_clk cell_2810 ( .C (clk), .D (signal_4003), .Q (signal_4004) ) ;
    buf_clk cell_2818 ( .C (clk), .D (signal_4011), .Q (signal_4012) ) ;
    buf_clk cell_2826 ( .C (clk), .D (signal_4019), .Q (signal_4020) ) ;
    buf_clk cell_2834 ( .C (clk), .D (signal_4027), .Q (signal_4028) ) ;
    buf_clk cell_2842 ( .C (clk), .D (signal_4035), .Q (signal_4036) ) ;
    buf_clk cell_2850 ( .C (clk), .D (signal_4043), .Q (signal_4044) ) ;
    buf_clk cell_2858 ( .C (clk), .D (signal_4051), .Q (signal_4052) ) ;
    buf_clk cell_2866 ( .C (clk), .D (signal_4059), .Q (signal_4060) ) ;
    buf_clk cell_2874 ( .C (clk), .D (signal_4067), .Q (signal_4068) ) ;
    buf_clk cell_2882 ( .C (clk), .D (signal_4075), .Q (signal_4076) ) ;
    buf_clk cell_2890 ( .C (clk), .D (signal_4083), .Q (signal_4084) ) ;
    buf_clk cell_2898 ( .C (clk), .D (signal_4091), .Q (signal_4092) ) ;
    buf_clk cell_2906 ( .C (clk), .D (signal_4099), .Q (signal_4100) ) ;
    buf_clk cell_2914 ( .C (clk), .D (signal_4107), .Q (signal_4108) ) ;
    buf_clk cell_2922 ( .C (clk), .D (signal_4115), .Q (signal_4116) ) ;
    buf_clk cell_2930 ( .C (clk), .D (signal_4123), .Q (signal_4124) ) ;
    buf_clk cell_2938 ( .C (clk), .D (signal_4131), .Q (signal_4132) ) ;
    buf_clk cell_2946 ( .C (clk), .D (signal_4139), .Q (signal_4140) ) ;
    buf_clk cell_2954 ( .C (clk), .D (signal_4147), .Q (signal_4148) ) ;
    buf_clk cell_2962 ( .C (clk), .D (signal_4155), .Q (signal_4156) ) ;
    buf_clk cell_2970 ( .C (clk), .D (signal_4163), .Q (signal_4164) ) ;
    buf_clk cell_2978 ( .C (clk), .D (signal_4171), .Q (signal_4172) ) ;
    buf_clk cell_2986 ( .C (clk), .D (signal_4179), .Q (signal_4180) ) ;
    buf_clk cell_2994 ( .C (clk), .D (signal_4187), .Q (signal_4188) ) ;
    buf_clk cell_3002 ( .C (clk), .D (signal_4195), .Q (signal_4196) ) ;
    buf_clk cell_3010 ( .C (clk), .D (signal_4203), .Q (signal_4204) ) ;
    buf_clk cell_3018 ( .C (clk), .D (signal_4211), .Q (signal_4212) ) ;
    buf_clk cell_3026 ( .C (clk), .D (signal_4219), .Q (signal_4220) ) ;
    buf_clk cell_3034 ( .C (clk), .D (signal_4227), .Q (signal_4228) ) ;
    buf_clk cell_3042 ( .C (clk), .D (signal_4235), .Q (signal_4236) ) ;
    buf_clk cell_3050 ( .C (clk), .D (signal_4243), .Q (signal_4244) ) ;
    buf_clk cell_3058 ( .C (clk), .D (signal_4251), .Q (signal_4252) ) ;
    buf_clk cell_3066 ( .C (clk), .D (signal_4259), .Q (signal_4260) ) ;
    buf_clk cell_3074 ( .C (clk), .D (signal_4267), .Q (signal_4268) ) ;
    buf_clk cell_3082 ( .C (clk), .D (signal_4275), .Q (signal_4276) ) ;
    buf_clk cell_3090 ( .C (clk), .D (signal_4283), .Q (signal_4284) ) ;
    buf_clk cell_3098 ( .C (clk), .D (signal_4291), .Q (signal_4292) ) ;
    buf_clk cell_3106 ( .C (clk), .D (signal_4299), .Q (signal_4300) ) ;
    buf_clk cell_3114 ( .C (clk), .D (signal_4307), .Q (signal_4308) ) ;
    buf_clk cell_3122 ( .C (clk), .D (signal_4315), .Q (signal_4316) ) ;
    buf_clk cell_3130 ( .C (clk), .D (signal_4323), .Q (signal_4324) ) ;
    buf_clk cell_3138 ( .C (clk), .D (signal_4331), .Q (signal_4332) ) ;
    buf_clk cell_3146 ( .C (clk), .D (signal_4339), .Q (signal_4340) ) ;
    buf_clk cell_3154 ( .C (clk), .D (signal_4347), .Q (signal_4348) ) ;
    buf_clk cell_3162 ( .C (clk), .D (signal_4355), .Q (signal_4356) ) ;
    buf_clk cell_3490 ( .C (clk), .D (signal_4683), .Q (signal_4684) ) ;
    buf_clk cell_3498 ( .C (clk), .D (signal_4691), .Q (signal_4692) ) ;
    buf_clk cell_3506 ( .C (clk), .D (signal_4699), .Q (signal_4700) ) ;
    buf_clk cell_3514 ( .C (clk), .D (signal_4707), .Q (signal_4708) ) ;
    buf_clk cell_3522 ( .C (clk), .D (signal_4715), .Q (signal_4716) ) ;
    buf_clk cell_3530 ( .C (clk), .D (signal_4723), .Q (signal_4724) ) ;
    buf_clk cell_3538 ( .C (clk), .D (signal_4731), .Q (signal_4732) ) ;
    buf_clk cell_3546 ( .C (clk), .D (signal_4739), .Q (signal_4740) ) ;
    buf_clk cell_3554 ( .C (clk), .D (signal_4747), .Q (signal_4748) ) ;
    buf_clk cell_3562 ( .C (clk), .D (signal_4755), .Q (signal_4756) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_856 ( .s ({signal_2245, signal_2243}), .b ({signal_1214, signal_1037}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[37]), .c ({signal_1291, signal_1056}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_857 ( .s ({signal_2249, signal_2247}), .b ({signal_1217, signal_1040}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[38]), .c ({signal_1292, signal_1057}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_858 ( .s ({signal_2253, signal_2251}), .b ({signal_1193, signal_1023}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[39]), .c ({signal_1294, signal_1058}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_859 ( .s ({signal_2257, signal_2255}), .b ({signal_1196, signal_1025}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[40]), .c ({signal_1296, signal_1059}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_860 ( .s ({signal_2261, signal_2259}), .b ({signal_1209, signal_1033}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[41]), .c ({signal_1298, signal_1060}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_861 ( .s ({signal_2265, signal_2263}), .b ({signal_1185, signal_1019}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[42]), .c ({signal_1300, signal_1061}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_862 ( .s ({signal_2269, signal_2267}), .b ({signal_1202, signal_1028}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[43]), .c ({signal_1302, signal_1062}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_863 ( .s ({signal_2273, signal_2271}), .b ({signal_1191, signal_1022}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[44]), .c ({signal_1304, signal_1063}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_864 ( .s ({signal_2277, signal_2275}), .b ({signal_1216, signal_1039}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[45]), .c ({signal_1306, signal_1064}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_865 ( .s ({signal_2281, signal_2279}), .b ({signal_1200, signal_1027}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[46]), .c ({signal_1308, signal_1065}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_866 ( .s ({signal_2285, signal_2283}), .b ({1'b0, 1'b0}), .a ({signal_1191, signal_1022}), .clk (clk), .r (Fresh[47]), .c ({signal_1310, signal_1066}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_867 ( .s ({signal_2289, signal_2287}), .b ({1'b0, 1'b1}), .a ({signal_1193, signal_1023}), .clk (clk), .r (Fresh[48]), .c ({signal_1312, signal_1067}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_868 ( .s ({signal_2269, signal_2267}), .b ({1'b0, 1'b0}), .a ({signal_1203, signal_1029}), .clk (clk), .r (Fresh[49]), .c ({signal_1313, signal_1068}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_869 ( .s ({signal_2293, signal_2291}), .b ({signal_1210, signal_1034}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[50]), .c ({signal_1315, signal_1069}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_870 ( .s ({signal_2285, signal_2283}), .b ({1'b0, 1'b1}), .a ({signal_1191, signal_1022}), .clk (clk), .r (Fresh[51]), .c ({signal_1316, signal_1070}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_871 ( .s ({signal_2249, signal_2247}), .b ({1'b0, 1'b1}), .a ({signal_1212, signal_1035}), .clk (clk), .r (Fresh[52]), .c ({signal_1317, signal_1071}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_872 ( .s ({signal_2285, signal_2283}), .b ({signal_1213, signal_1036}), .a ({signal_1191, signal_1022}), .clk (clk), .r (Fresh[53]), .c ({signal_1318, signal_1072}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_873 ( .s ({signal_2265, signal_2263}), .b ({1'b0, 1'b1}), .a ({signal_1185, signal_1019}), .clk (clk), .r (Fresh[54]), .c ({signal_1319, signal_1073}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_874 ( .s ({signal_2277, signal_2275}), .b ({1'b0, 1'b1}), .a ({signal_1200, signal_1027}), .clk (clk), .r (Fresh[55]), .c ({signal_1320, signal_1074}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_875 ( .s ({signal_2289, signal_2287}), .b ({signal_1193, signal_1023}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[56]), .c ({signal_1321, signal_1075}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_876 ( .s ({signal_2293, signal_2291}), .b ({1'b0, 1'b0}), .a ({signal_1205, signal_1030}), .clk (clk), .r (Fresh[57]), .c ({signal_1322, signal_1076}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_877 ( .s ({signal_2249, signal_2247}), .b ({signal_1217, signal_1040}), .a ({signal_1212, signal_1035}), .clk (clk), .r (Fresh[58]), .c ({signal_1323, signal_1077}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_878 ( .s ({signal_2285, signal_2283}), .b ({signal_1213, signal_1036}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[59]), .c ({signal_1324, signal_1078}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_879 ( .s ({signal_2249, signal_2247}), .b ({1'b0, 1'b1}), .a ({signal_1217, signal_1040}), .clk (clk), .r (Fresh[60]), .c ({signal_1325, signal_1079}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_880 ( .s ({signal_2297, signal_2295}), .b ({1'b0, 1'b1}), .a ({signal_1209, signal_1033}), .clk (clk), .r (Fresh[61]), .c ({signal_1327, signal_1080}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_881 ( .s ({signal_2289, signal_2287}), .b ({signal_1215, signal_1038}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[62]), .c ({signal_1328, signal_1081}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_882 ( .s ({signal_2277, signal_2275}), .b ({signal_1200, signal_1027}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[63]), .c ({signal_1329, signal_1082}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_883 ( .s ({signal_2297, signal_2295}), .b ({1'b0, 1'b0}), .a ({signal_1209, signal_1033}), .clk (clk), .r (Fresh[64]), .c ({signal_1330, signal_1083}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_884 ( .s ({signal_2301, signal_2299}), .b ({signal_1208, signal_1032}), .a ({signal_1196, signal_1025}), .clk (clk), .r (Fresh[65]), .c ({signal_1332, signal_1084}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_885 ( .s ({signal_2277, signal_2275}), .b ({signal_1216, signal_1039}), .a ({signal_1200, signal_1027}), .clk (clk), .r (Fresh[66]), .c ({signal_1333, signal_1085}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_886 ( .s ({signal_2301, signal_2299}), .b ({signal_1208, signal_1032}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[67]), .c ({signal_1334, signal_1086}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_887 ( .s ({signal_2297, signal_2295}), .b ({signal_1209, signal_1033}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[68]), .c ({signal_1335, signal_1087}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_888 ( .s ({signal_2245, signal_2243}), .b ({1'b0, 1'b0}), .a ({signal_1214, signal_1037}), .clk (clk), .r (Fresh[69]), .c ({signal_1336, signal_1088}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_889 ( .s ({signal_2269, signal_2267}), .b ({1'b0, 1'b1}), .a ({signal_1203, signal_1029}), .clk (clk), .r (Fresh[70]), .c ({signal_1337, signal_1089}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_890 ( .s ({signal_2301, signal_2299}), .b ({1'b0, 1'b1}), .a ({signal_1196, signal_1025}), .clk (clk), .r (Fresh[71]), .c ({signal_1338, signal_1090}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_891 ( .s ({signal_2265, signal_2263}), .b ({signal_1194, signal_1024}), .a ({signal_1185, signal_1019}), .clk (clk), .r (Fresh[72]), .c ({signal_1339, signal_1091}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_892 ( .s ({signal_2289, signal_2287}), .b ({signal_1215, signal_1038}), .a ({signal_1193, signal_1023}), .clk (clk), .r (Fresh[73]), .c ({signal_1340, signal_1092}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_893 ( .s ({signal_2305, signal_2303}), .b ({signal_1214, signal_1037}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[74]), .c ({signal_1342, signal_1093}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_894 ( .s ({signal_2277, signal_2275}), .b ({1'b0, 1'b0}), .a ({signal_1200, signal_1027}), .clk (clk), .r (Fresh[75]), .c ({signal_1343, signal_1094}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_895 ( .s ({signal_2293, signal_2291}), .b ({1'b0, 1'b1}), .a ({signal_1205, signal_1030}), .clk (clk), .r (Fresh[76]), .c ({signal_1344, signal_1095}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_896 ( .s ({signal_2245, signal_2243}), .b ({1'b0, 1'b1}), .a ({signal_1214, signal_1037}), .clk (clk), .r (Fresh[77]), .c ({signal_1345, signal_1096}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_897 ( .s ({signal_2293, signal_2291}), .b ({signal_1205, signal_1030}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[78]), .c ({signal_1346, signal_1097}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_898 ( .s ({signal_2269, signal_2267}), .b ({signal_1202, signal_1028}), .a ({signal_1203, signal_1029}), .clk (clk), .r (Fresh[79]), .c ({signal_1347, signal_1098}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_899 ( .s ({signal_2285, signal_2283}), .b ({signal_1191, signal_1022}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[80]), .c ({signal_1348, signal_1099}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_900 ( .s ({signal_2297, signal_2295}), .b ({signal_1187, signal_1020}), .a ({signal_1209, signal_1033}), .clk (clk), .r (Fresh[81]), .c ({signal_1349, signal_1100}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_901 ( .s ({signal_2269, signal_2267}), .b ({signal_1203, signal_1029}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[82]), .c ({signal_1350, signal_1101}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_902 ( .s ({signal_2301, signal_2299}), .b ({1'b0, 1'b0}), .a ({signal_1196, signal_1025}), .clk (clk), .r (Fresh[83]), .c ({signal_1351, signal_1102}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_903 ( .s ({signal_2309, signal_2307}), .b ({signal_1205, signal_1030}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[84]), .c ({signal_1353, signal_1103}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_904 ( .s ({signal_2245, signal_2243}), .b ({signal_1198, signal_1026}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[85]), .c ({signal_1354, signal_1104}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_905 ( .s ({signal_2301, signal_2299}), .b ({signal_1196, signal_1025}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[86]), .c ({signal_1355, signal_1105}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_906 ( .s ({signal_2313, signal_2311}), .b ({signal_1189, signal_1021}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[87]), .c ({signal_1357, signal_1106}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_907 ( .s ({signal_2249, signal_2247}), .b ({signal_1217, signal_1040}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[88]), .c ({signal_1358, signal_1107}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_908 ( .s ({signal_2265, signal_2263}), .b ({1'b0, 1'b0}), .a ({signal_1185, signal_1019}), .clk (clk), .r (Fresh[89]), .c ({signal_1359, signal_1108}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_909 ( .s ({signal_2317, signal_2315}), .b ({signal_1203, signal_1029}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[90]), .c ({signal_1361, signal_1109}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_910 ( .s ({signal_2245, signal_2243}), .b ({signal_1198, signal_1026}), .a ({signal_1214, signal_1037}), .clk (clk), .r (Fresh[91]), .c ({signal_1362, signal_1110}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_911 ( .s ({signal_2297, signal_2295}), .b ({signal_1187, signal_1020}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[92]), .c ({signal_1363, signal_1111}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_912 ( .s ({signal_2289, signal_2287}), .b ({1'b0, 1'b0}), .a ({signal_1193, signal_1023}), .clk (clk), .r (Fresh[93]), .c ({signal_1364, signal_1112}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_913 ( .s ({signal_2265, signal_2263}), .b ({signal_1194, signal_1024}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[94]), .c ({signal_1365, signal_1113}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_914 ( .s ({signal_2321, signal_2319}), .b ({signal_1185, signal_1019}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[95]), .c ({signal_1367, signal_1114}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_915 ( .s ({signal_2293, signal_2291}), .b ({signal_1210, signal_1034}), .a ({signal_1205, signal_1030}), .clk (clk), .r (Fresh[96]), .c ({signal_1368, signal_1115}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_916 ( .s ({signal_2325, signal_2323}), .b ({1'b0, 1'b1}), .a ({signal_1218, signal_1041}), .clk (clk), .r (Fresh[97]), .c ({signal_1370, signal_1116}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_917 ( .s ({signal_2325, signal_2323}), .b ({signal_1207, signal_1031}), .a ({signal_1218, signal_1041}), .clk (clk), .r (Fresh[98]), .c ({signal_1371, signal_1117}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_918 ( .s ({signal_2325, signal_2323}), .b ({signal_1218, signal_1041}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[99]), .c ({signal_1372, signal_1118}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_919 ( .s ({signal_2325, signal_2323}), .b ({1'b0, 1'b0}), .a ({signal_1218, signal_1041}), .clk (clk), .r (Fresh[100]), .c ({signal_1373, signal_1119}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_920 ( .s ({signal_2325, signal_2323}), .b ({signal_1207, signal_1031}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[101]), .c ({signal_1374, signal_1120}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_921 ( .s ({signal_2329, signal_2327}), .b ({signal_1218, signal_1041}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[102]), .c ({signal_1376, signal_1121}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_922 ( .s ({signal_2333, signal_2331}), .b ({1'b0, 1'b1}), .a ({signal_1221, signal_1043}), .clk (clk), .r (Fresh[103]), .c ({signal_1377, signal_1122}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_923 ( .s ({signal_2333, signal_2331}), .b ({signal_1220, signal_1042}), .a ({signal_1221, signal_1043}), .clk (clk), .r (Fresh[104]), .c ({signal_1378, signal_1123}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_924 ( .s ({signal_2333, signal_2331}), .b ({1'b0, 1'b1}), .a ({signal_1220, signal_1042}), .clk (clk), .r (Fresh[105]), .c ({signal_1379, signal_1124}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_925 ( .s ({signal_2333, signal_2331}), .b ({signal_1220, signal_1042}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[106]), .c ({signal_1380, signal_1125}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_926 ( .s ({signal_2333, signal_2331}), .b ({signal_1220, signal_1042}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[107]), .c ({signal_1381, signal_1126}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_927 ( .s ({signal_2337, signal_2335}), .b ({signal_1223, signal_1044}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[108]), .c ({signal_1383, signal_1127}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_928 ( .s ({signal_2341, signal_2339}), .b ({1'b0, 1'b1}), .a ({signal_1226, signal_1046}), .clk (clk), .r (Fresh[109]), .c ({signal_1384, signal_1128}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_929 ( .s ({signal_2341, signal_2339}), .b ({signal_1225, signal_1045}), .a ({signal_1226, signal_1046}), .clk (clk), .r (Fresh[110]), .c ({signal_1385, signal_1129}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_930 ( .s ({signal_2341, signal_2339}), .b ({1'b0, 1'b1}), .a ({signal_1225, signal_1045}), .clk (clk), .r (Fresh[111]), .c ({signal_1386, signal_1130}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_931 ( .s ({signal_2341, signal_2339}), .b ({signal_1225, signal_1045}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[112]), .c ({signal_1387, signal_1131}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_932 ( .s ({signal_2341, signal_2339}), .b ({signal_1225, signal_1045}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[113]), .c ({signal_1388, signal_1132}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_933 ( .s ({signal_2345, signal_2343}), .b ({signal_1228, signal_1047}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[114]), .c ({signal_1390, signal_1133}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_934 ( .s ({signal_2349, signal_2347}), .b ({1'b0, 1'b1}), .a ({signal_1231, signal_1049}), .clk (clk), .r (Fresh[115]), .c ({signal_1391, signal_1134}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_935 ( .s ({signal_2349, signal_2347}), .b ({signal_1230, signal_1048}), .a ({signal_1231, signal_1049}), .clk (clk), .r (Fresh[116]), .c ({signal_1392, signal_1135}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_936 ( .s ({signal_2349, signal_2347}), .b ({1'b0, 1'b1}), .a ({signal_1230, signal_1048}), .clk (clk), .r (Fresh[117]), .c ({signal_1393, signal_1136}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_937 ( .s ({signal_2349, signal_2347}), .b ({signal_1230, signal_1048}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[118]), .c ({signal_1394, signal_1137}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_938 ( .s ({signal_2349, signal_2347}), .b ({signal_1230, signal_1048}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[119]), .c ({signal_1395, signal_1138}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_939 ( .s ({signal_2353, signal_2351}), .b ({signal_1233, signal_1050}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[120]), .c ({signal_1397, signal_1139}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_940 ( .s ({signal_2357, signal_2355}), .b ({1'b0, 1'b1}), .a ({signal_1236, signal_1052}), .clk (clk), .r (Fresh[121]), .c ({signal_1398, signal_1140}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_941 ( .s ({signal_2357, signal_2355}), .b ({signal_1235, signal_1051}), .a ({signal_1236, signal_1052}), .clk (clk), .r (Fresh[122]), .c ({signal_1399, signal_1141}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_942 ( .s ({signal_2357, signal_2355}), .b ({1'b0, 1'b1}), .a ({signal_1235, signal_1051}), .clk (clk), .r (Fresh[123]), .c ({signal_1400, signal_1142}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_943 ( .s ({signal_2357, signal_2355}), .b ({signal_1235, signal_1051}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[124]), .c ({signal_1401, signal_1143}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_944 ( .s ({signal_2357, signal_2355}), .b ({signal_1235, signal_1051}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[125]), .c ({signal_1402, signal_1144}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_945 ( .s ({signal_2361, signal_2359}), .b ({signal_1238, signal_1053}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[126]), .c ({signal_1404, signal_1145}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_946 ( .s ({signal_2365, signal_2363}), .b ({1'b0, 1'b1}), .a ({signal_1241, signal_1055}), .clk (clk), .r (Fresh[127]), .c ({signal_1406, signal_1146}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_947 ( .s ({signal_2365, signal_2363}), .b ({signal_1240, signal_1054}), .a ({signal_1241, signal_1055}), .clk (clk), .r (Fresh[128]), .c ({signal_1407, signal_1147}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_948 ( .s ({signal_2365, signal_2363}), .b ({signal_1241, signal_1055}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[129]), .c ({signal_1408, signal_1148}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_949 ( .s ({signal_2365, signal_2363}), .b ({1'b0, 1'b0}), .a ({signal_1241, signal_1055}), .clk (clk), .r (Fresh[130]), .c ({signal_1409, signal_1149}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_950 ( .s ({signal_2365, signal_2363}), .b ({signal_1240, signal_1054}), .a ({1'b0, 1'b1}), .clk (clk), .r (Fresh[131]), .c ({signal_1410, signal_1150}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_951 ( .s ({signal_2369, signal_2367}), .b ({signal_1241, signal_1055}), .a ({1'b0, 1'b0}), .clk (clk), .r (Fresh[132]), .c ({signal_1412, signal_1151}) ) ;
    buf_clk cell_1179 ( .C (clk), .D (signal_2372), .Q (signal_2373) ) ;
    buf_clk cell_1185 ( .C (clk), .D (signal_2378), .Q (signal_2379) ) ;
    buf_clk cell_1191 ( .C (clk), .D (signal_2384), .Q (signal_2385) ) ;
    buf_clk cell_1197 ( .C (clk), .D (signal_2390), .Q (signal_2391) ) ;
    buf_clk cell_1203 ( .C (clk), .D (signal_2396), .Q (signal_2397) ) ;
    buf_clk cell_1209 ( .C (clk), .D (signal_2402), .Q (signal_2403) ) ;
    buf_clk cell_1215 ( .C (clk), .D (signal_2408), .Q (signal_2409) ) ;
    buf_clk cell_1221 ( .C (clk), .D (signal_2414), .Q (signal_2415) ) ;
    buf_clk cell_1227 ( .C (clk), .D (signal_2420), .Q (signal_2421) ) ;
    buf_clk cell_1233 ( .C (clk), .D (signal_2426), .Q (signal_2427) ) ;
    buf_clk cell_1239 ( .C (clk), .D (signal_2432), .Q (signal_2433) ) ;
    buf_clk cell_1245 ( .C (clk), .D (signal_2438), .Q (signal_2439) ) ;
    buf_clk cell_1251 ( .C (clk), .D (signal_2444), .Q (signal_2445) ) ;
    buf_clk cell_1257 ( .C (clk), .D (signal_2450), .Q (signal_2451) ) ;
    buf_clk cell_1263 ( .C (clk), .D (signal_2456), .Q (signal_2457) ) ;
    buf_clk cell_1269 ( .C (clk), .D (signal_2462), .Q (signal_2463) ) ;
    buf_clk cell_1275 ( .C (clk), .D (signal_2468), .Q (signal_2469) ) ;
    buf_clk cell_1281 ( .C (clk), .D (signal_2474), .Q (signal_2475) ) ;
    buf_clk cell_1287 ( .C (clk), .D (signal_2480), .Q (signal_2481) ) ;
    buf_clk cell_1293 ( .C (clk), .D (signal_2486), .Q (signal_2487) ) ;
    buf_clk cell_1299 ( .C (clk), .D (signal_2492), .Q (signal_2493) ) ;
    buf_clk cell_1305 ( .C (clk), .D (signal_2498), .Q (signal_2499) ) ;
    buf_clk cell_1311 ( .C (clk), .D (signal_2504), .Q (signal_2505) ) ;
    buf_clk cell_1317 ( .C (clk), .D (signal_2510), .Q (signal_2511) ) ;
    buf_clk cell_1323 ( .C (clk), .D (signal_2516), .Q (signal_2517) ) ;
    buf_clk cell_1329 ( .C (clk), .D (signal_2522), .Q (signal_2523) ) ;
    buf_clk cell_1335 ( .C (clk), .D (signal_2528), .Q (signal_2529) ) ;
    buf_clk cell_1341 ( .C (clk), .D (signal_2534), .Q (signal_2535) ) ;
    buf_clk cell_1347 ( .C (clk), .D (signal_2540), .Q (signal_2541) ) ;
    buf_clk cell_1353 ( .C (clk), .D (signal_2546), .Q (signal_2547) ) ;
    buf_clk cell_1359 ( .C (clk), .D (signal_2552), .Q (signal_2553) ) ;
    buf_clk cell_1365 ( .C (clk), .D (signal_2558), .Q (signal_2559) ) ;
    buf_clk cell_1371 ( .C (clk), .D (signal_2564), .Q (signal_2565) ) ;
    buf_clk cell_1377 ( .C (clk), .D (signal_2570), .Q (signal_2571) ) ;
    buf_clk cell_1383 ( .C (clk), .D (signal_2576), .Q (signal_2577) ) ;
    buf_clk cell_1389 ( .C (clk), .D (signal_2582), .Q (signal_2583) ) ;
    buf_clk cell_1395 ( .C (clk), .D (signal_2588), .Q (signal_2589) ) ;
    buf_clk cell_1401 ( .C (clk), .D (signal_2594), .Q (signal_2595) ) ;
    buf_clk cell_1407 ( .C (clk), .D (signal_2600), .Q (signal_2601) ) ;
    buf_clk cell_1413 ( .C (clk), .D (signal_2606), .Q (signal_2607) ) ;
    buf_clk cell_1419 ( .C (clk), .D (signal_2612), .Q (signal_2613) ) ;
    buf_clk cell_1425 ( .C (clk), .D (signal_2618), .Q (signal_2619) ) ;
    buf_clk cell_1431 ( .C (clk), .D (signal_2624), .Q (signal_2625) ) ;
    buf_clk cell_1437 ( .C (clk), .D (signal_2630), .Q (signal_2631) ) ;
    buf_clk cell_1443 ( .C (clk), .D (signal_2636), .Q (signal_2637) ) ;
    buf_clk cell_1449 ( .C (clk), .D (signal_2642), .Q (signal_2643) ) ;
    buf_clk cell_1455 ( .C (clk), .D (signal_2648), .Q (signal_2649) ) ;
    buf_clk cell_1461 ( .C (clk), .D (signal_2654), .Q (signal_2655) ) ;
    buf_clk cell_1467 ( .C (clk), .D (signal_2660), .Q (signal_2661) ) ;
    buf_clk cell_1473 ( .C (clk), .D (signal_2666), .Q (signal_2667) ) ;
    buf_clk cell_1479 ( .C (clk), .D (signal_2672), .Q (signal_2673) ) ;
    buf_clk cell_1485 ( .C (clk), .D (signal_2678), .Q (signal_2679) ) ;
    buf_clk cell_1491 ( .C (clk), .D (signal_2684), .Q (signal_2685) ) ;
    buf_clk cell_1497 ( .C (clk), .D (signal_2690), .Q (signal_2691) ) ;
    buf_clk cell_1503 ( .C (clk), .D (signal_2696), .Q (signal_2697) ) ;
    buf_clk cell_1509 ( .C (clk), .D (signal_2702), .Q (signal_2703) ) ;
    buf_clk cell_1515 ( .C (clk), .D (signal_2708), .Q (signal_2709) ) ;
    buf_clk cell_1521 ( .C (clk), .D (signal_2714), .Q (signal_2715) ) ;
    buf_clk cell_1527 ( .C (clk), .D (signal_2720), .Q (signal_2721) ) ;
    buf_clk cell_1533 ( .C (clk), .D (signal_2726), .Q (signal_2727) ) ;
    buf_clk cell_1539 ( .C (clk), .D (signal_2732), .Q (signal_2733) ) ;
    buf_clk cell_1545 ( .C (clk), .D (signal_2738), .Q (signal_2739) ) ;
    buf_clk cell_1551 ( .C (clk), .D (signal_2744), .Q (signal_2745) ) ;
    buf_clk cell_1557 ( .C (clk), .D (signal_2750), .Q (signal_2751) ) ;
    buf_clk cell_1563 ( .C (clk), .D (signal_2756), .Q (signal_2757) ) ;
    buf_clk cell_1569 ( .C (clk), .D (signal_2762), .Q (signal_2763) ) ;
    buf_clk cell_1575 ( .C (clk), .D (signal_2768), .Q (signal_2769) ) ;
    buf_clk cell_1581 ( .C (clk), .D (signal_2774), .Q (signal_2775) ) ;
    buf_clk cell_1587 ( .C (clk), .D (signal_2780), .Q (signal_2781) ) ;
    buf_clk cell_1593 ( .C (clk), .D (signal_2786), .Q (signal_2787) ) ;
    buf_clk cell_1599 ( .C (clk), .D (signal_2792), .Q (signal_2793) ) ;
    buf_clk cell_1605 ( .C (clk), .D (signal_2798), .Q (signal_2799) ) ;
    buf_clk cell_1611 ( .C (clk), .D (signal_2804), .Q (signal_2805) ) ;
    buf_clk cell_1617 ( .C (clk), .D (signal_2810), .Q (signal_2811) ) ;
    buf_clk cell_1623 ( .C (clk), .D (signal_2816), .Q (signal_2817) ) ;
    buf_clk cell_1629 ( .C (clk), .D (signal_2822), .Q (signal_2823) ) ;
    buf_clk cell_1635 ( .C (clk), .D (signal_2828), .Q (signal_2829) ) ;
    buf_clk cell_1641 ( .C (clk), .D (signal_2834), .Q (signal_2835) ) ;
    buf_clk cell_1647 ( .C (clk), .D (signal_2840), .Q (signal_2841) ) ;
    buf_clk cell_1653 ( .C (clk), .D (signal_2846), .Q (signal_2847) ) ;
    buf_clk cell_1659 ( .C (clk), .D (signal_2852), .Q (signal_2853) ) ;
    buf_clk cell_1665 ( .C (clk), .D (signal_2858), .Q (signal_2859) ) ;
    buf_clk cell_1671 ( .C (clk), .D (signal_2864), .Q (signal_2865) ) ;
    buf_clk cell_1677 ( .C (clk), .D (signal_2870), .Q (signal_2871) ) ;
    buf_clk cell_1683 ( .C (clk), .D (signal_2876), .Q (signal_2877) ) ;
    buf_clk cell_1689 ( .C (clk), .D (signal_2882), .Q (signal_2883) ) ;
    buf_clk cell_1695 ( .C (clk), .D (signal_2888), .Q (signal_2889) ) ;
    buf_clk cell_1701 ( .C (clk), .D (signal_2894), .Q (signal_2895) ) ;
    buf_clk cell_1707 ( .C (clk), .D (signal_2900), .Q (signal_2901) ) ;
    buf_clk cell_1713 ( .C (clk), .D (signal_2906), .Q (signal_2907) ) ;
    buf_clk cell_1719 ( .C (clk), .D (signal_2912), .Q (signal_2913) ) ;
    buf_clk cell_1725 ( .C (clk), .D (signal_2918), .Q (signal_2919) ) ;
    buf_clk cell_1731 ( .C (clk), .D (signal_2924), .Q (signal_2925) ) ;
    buf_clk cell_1737 ( .C (clk), .D (signal_2930), .Q (signal_2931) ) ;
    buf_clk cell_1743 ( .C (clk), .D (signal_2936), .Q (signal_2937) ) ;
    buf_clk cell_1749 ( .C (clk), .D (signal_2942), .Q (signal_2943) ) ;
    buf_clk cell_1755 ( .C (clk), .D (signal_2948), .Q (signal_2949) ) ;
    buf_clk cell_1761 ( .C (clk), .D (signal_2954), .Q (signal_2955) ) ;
    buf_clk cell_1767 ( .C (clk), .D (signal_2960), .Q (signal_2961) ) ;
    buf_clk cell_1773 ( .C (clk), .D (signal_2966), .Q (signal_2967) ) ;
    buf_clk cell_1779 ( .C (clk), .D (signal_2972), .Q (signal_2973) ) ;
    buf_clk cell_1785 ( .C (clk), .D (signal_2978), .Q (signal_2979) ) ;
    buf_clk cell_1791 ( .C (clk), .D (signal_2984), .Q (signal_2985) ) ;
    buf_clk cell_1797 ( .C (clk), .D (signal_2990), .Q (signal_2991) ) ;
    buf_clk cell_1803 ( .C (clk), .D (signal_2996), .Q (signal_2997) ) ;
    buf_clk cell_1809 ( .C (clk), .D (signal_3002), .Q (signal_3003) ) ;
    buf_clk cell_1815 ( .C (clk), .D (signal_3008), .Q (signal_3009) ) ;
    buf_clk cell_1821 ( .C (clk), .D (signal_3014), .Q (signal_3015) ) ;
    buf_clk cell_1827 ( .C (clk), .D (signal_3020), .Q (signal_3021) ) ;
    buf_clk cell_1833 ( .C (clk), .D (signal_3026), .Q (signal_3027) ) ;
    buf_clk cell_1839 ( .C (clk), .D (signal_3032), .Q (signal_3033) ) ;
    buf_clk cell_1845 ( .C (clk), .D (signal_3038), .Q (signal_3039) ) ;
    buf_clk cell_1851 ( .C (clk), .D (signal_3044), .Q (signal_3045) ) ;
    buf_clk cell_1857 ( .C (clk), .D (signal_3050), .Q (signal_3051) ) ;
    buf_clk cell_1863 ( .C (clk), .D (signal_3056), .Q (signal_3057) ) ;
    buf_clk cell_1869 ( .C (clk), .D (signal_3062), .Q (signal_3063) ) ;
    buf_clk cell_1875 ( .C (clk), .D (signal_3068), .Q (signal_3069) ) ;
    buf_clk cell_1881 ( .C (clk), .D (signal_3074), .Q (signal_3075) ) ;
    buf_clk cell_1887 ( .C (clk), .D (signal_3080), .Q (signal_3081) ) ;
    buf_clk cell_1893 ( .C (clk), .D (signal_3086), .Q (signal_3087) ) ;
    buf_clk cell_1899 ( .C (clk), .D (signal_3092), .Q (signal_3093) ) ;
    buf_clk cell_1905 ( .C (clk), .D (signal_3098), .Q (signal_3099) ) ;
    buf_clk cell_1911 ( .C (clk), .D (signal_3104), .Q (signal_3105) ) ;
    buf_clk cell_1917 ( .C (clk), .D (signal_3110), .Q (signal_3111) ) ;
    buf_clk cell_1923 ( .C (clk), .D (signal_3116), .Q (signal_3117) ) ;
    buf_clk cell_1929 ( .C (clk), .D (signal_3122), .Q (signal_3123) ) ;
    buf_clk cell_1935 ( .C (clk), .D (signal_3128), .Q (signal_3129) ) ;
    buf_clk cell_1941 ( .C (clk), .D (signal_3134), .Q (signal_3135) ) ;
    buf_clk cell_1947 ( .C (clk), .D (signal_3140), .Q (signal_3141) ) ;
    buf_clk cell_1951 ( .C (clk), .D (signal_3144), .Q (signal_3145) ) ;
    buf_clk cell_1953 ( .C (clk), .D (signal_3146), .Q (signal_3147) ) ;
    buf_clk cell_1957 ( .C (clk), .D (signal_3150), .Q (signal_3151) ) ;
    buf_clk cell_1961 ( .C (clk), .D (signal_3154), .Q (signal_3155) ) ;
    buf_clk cell_1963 ( .C (clk), .D (signal_3156), .Q (signal_3157) ) ;
    buf_clk cell_1965 ( .C (clk), .D (signal_3158), .Q (signal_3159) ) ;
    buf_clk cell_1967 ( .C (clk), .D (signal_3160), .Q (signal_3161) ) ;
    buf_clk cell_1969 ( .C (clk), .D (signal_3162), .Q (signal_3163) ) ;
    buf_clk cell_1971 ( .C (clk), .D (signal_3164), .Q (signal_3165) ) ;
    buf_clk cell_1973 ( .C (clk), .D (signal_3166), .Q (signal_3167) ) ;
    buf_clk cell_1975 ( .C (clk), .D (signal_3168), .Q (signal_3169) ) ;
    buf_clk cell_1977 ( .C (clk), .D (signal_3170), .Q (signal_3171) ) ;
    buf_clk cell_1979 ( .C (clk), .D (signal_3172), .Q (signal_3173) ) ;
    buf_clk cell_1981 ( .C (clk), .D (signal_3174), .Q (signal_3175) ) ;
    buf_clk cell_1983 ( .C (clk), .D (signal_3176), .Q (signal_3177) ) ;
    buf_clk cell_1985 ( .C (clk), .D (signal_3178), .Q (signal_3179) ) ;
    buf_clk cell_1989 ( .C (clk), .D (signal_3182), .Q (signal_3183) ) ;
    buf_clk cell_1993 ( .C (clk), .D (signal_3186), .Q (signal_3187) ) ;
    buf_clk cell_1997 ( .C (clk), .D (signal_3190), .Q (signal_3191) ) ;
    buf_clk cell_2001 ( .C (clk), .D (signal_3194), .Q (signal_3195) ) ;
    buf_clk cell_2003 ( .C (clk), .D (signal_3196), .Q (signal_3197) ) ;
    buf_clk cell_2005 ( .C (clk), .D (signal_3198), .Q (signal_3199) ) ;
    buf_clk cell_2007 ( .C (clk), .D (signal_3200), .Q (signal_3201) ) ;
    buf_clk cell_2009 ( .C (clk), .D (signal_3202), .Q (signal_3203) ) ;
    buf_clk cell_2013 ( .C (clk), .D (signal_3206), .Q (signal_3207) ) ;
    buf_clk cell_2017 ( .C (clk), .D (signal_3210), .Q (signal_3211) ) ;
    buf_clk cell_2021 ( .C (clk), .D (signal_3214), .Q (signal_3215) ) ;
    buf_clk cell_2025 ( .C (clk), .D (signal_3218), .Q (signal_3219) ) ;
    buf_clk cell_2027 ( .C (clk), .D (signal_3220), .Q (signal_3221) ) ;
    buf_clk cell_2029 ( .C (clk), .D (signal_3222), .Q (signal_3223) ) ;
    buf_clk cell_2033 ( .C (clk), .D (signal_3226), .Q (signal_3227) ) ;
    buf_clk cell_2037 ( .C (clk), .D (signal_3230), .Q (signal_3231) ) ;
    buf_clk cell_2041 ( .C (clk), .D (signal_3234), .Q (signal_3235) ) ;
    buf_clk cell_2045 ( .C (clk), .D (signal_3238), .Q (signal_3239) ) ;
    buf_clk cell_2049 ( .C (clk), .D (signal_3242), .Q (signal_3243) ) ;
    buf_clk cell_2053 ( .C (clk), .D (signal_3246), .Q (signal_3247) ) ;
    buf_clk cell_2057 ( .C (clk), .D (signal_3250), .Q (signal_3251) ) ;
    buf_clk cell_2061 ( .C (clk), .D (signal_3254), .Q (signal_3255) ) ;
    buf_clk cell_2065 ( .C (clk), .D (signal_3258), .Q (signal_3259) ) ;
    buf_clk cell_2069 ( .C (clk), .D (signal_3262), .Q (signal_3263) ) ;
    buf_clk cell_2071 ( .C (clk), .D (signal_3264), .Q (signal_3265) ) ;
    buf_clk cell_2073 ( .C (clk), .D (signal_3266), .Q (signal_3267) ) ;
    buf_clk cell_2077 ( .C (clk), .D (signal_3270), .Q (signal_3271) ) ;
    buf_clk cell_2081 ( .C (clk), .D (signal_3274), .Q (signal_3275) ) ;
    buf_clk cell_2083 ( .C (clk), .D (signal_3276), .Q (signal_3277) ) ;
    buf_clk cell_2085 ( .C (clk), .D (signal_3278), .Q (signal_3279) ) ;
    buf_clk cell_2089 ( .C (clk), .D (signal_3282), .Q (signal_3283) ) ;
    buf_clk cell_2093 ( .C (clk), .D (signal_3286), .Q (signal_3287) ) ;
    buf_clk cell_2095 ( .C (clk), .D (signal_3288), .Q (signal_3289) ) ;
    buf_clk cell_2097 ( .C (clk), .D (signal_3290), .Q (signal_3291) ) ;
    buf_clk cell_2101 ( .C (clk), .D (signal_3294), .Q (signal_3295) ) ;
    buf_clk cell_2105 ( .C (clk), .D (signal_3298), .Q (signal_3299) ) ;
    buf_clk cell_2107 ( .C (clk), .D (signal_3300), .Q (signal_3301) ) ;
    buf_clk cell_2109 ( .C (clk), .D (signal_3302), .Q (signal_3303) ) ;
    buf_clk cell_2113 ( .C (clk), .D (signal_3306), .Q (signal_3307) ) ;
    buf_clk cell_2117 ( .C (clk), .D (signal_3310), .Q (signal_3311) ) ;
    buf_clk cell_2119 ( .C (clk), .D (signal_3312), .Q (signal_3313) ) ;
    buf_clk cell_2121 ( .C (clk), .D (signal_3314), .Q (signal_3315) ) ;
    buf_clk cell_2125 ( .C (clk), .D (signal_3318), .Q (signal_3319) ) ;
    buf_clk cell_2129 ( .C (clk), .D (signal_3322), .Q (signal_3323) ) ;
    buf_clk cell_2131 ( .C (clk), .D (signal_3324), .Q (signal_3325) ) ;
    buf_clk cell_2133 ( .C (clk), .D (signal_3326), .Q (signal_3327) ) ;
    buf_clk cell_2137 ( .C (clk), .D (signal_3330), .Q (signal_3331) ) ;
    buf_clk cell_2141 ( .C (clk), .D (signal_3334), .Q (signal_3335) ) ;
    buf_clk cell_2147 ( .C (clk), .D (signal_3340), .Q (signal_3341) ) ;
    buf_clk cell_2155 ( .C (clk), .D (signal_3348), .Q (signal_3349) ) ;
    buf_clk cell_2163 ( .C (clk), .D (signal_3356), .Q (signal_3357) ) ;
    buf_clk cell_2171 ( .C (clk), .D (signal_3364), .Q (signal_3365) ) ;
    buf_clk cell_2179 ( .C (clk), .D (signal_3372), .Q (signal_3373) ) ;
    buf_clk cell_2187 ( .C (clk), .D (signal_3380), .Q (signal_3381) ) ;
    buf_clk cell_2195 ( .C (clk), .D (signal_3388), .Q (signal_3389) ) ;
    buf_clk cell_2203 ( .C (clk), .D (signal_3396), .Q (signal_3397) ) ;
    buf_clk cell_2211 ( .C (clk), .D (signal_3404), .Q (signal_3405) ) ;
    buf_clk cell_2219 ( .C (clk), .D (signal_3412), .Q (signal_3413) ) ;
    buf_clk cell_2227 ( .C (clk), .D (signal_3420), .Q (signal_3421) ) ;
    buf_clk cell_2235 ( .C (clk), .D (signal_3428), .Q (signal_3429) ) ;
    buf_clk cell_2243 ( .C (clk), .D (signal_3436), .Q (signal_3437) ) ;
    buf_clk cell_2251 ( .C (clk), .D (signal_3444), .Q (signal_3445) ) ;
    buf_clk cell_2259 ( .C (clk), .D (signal_3452), .Q (signal_3453) ) ;
    buf_clk cell_2267 ( .C (clk), .D (signal_3460), .Q (signal_3461) ) ;
    buf_clk cell_2275 ( .C (clk), .D (signal_3468), .Q (signal_3469) ) ;
    buf_clk cell_2283 ( .C (clk), .D (signal_3476), .Q (signal_3477) ) ;
    buf_clk cell_2291 ( .C (clk), .D (signal_3484), .Q (signal_3485) ) ;
    buf_clk cell_2299 ( .C (clk), .D (signal_3492), .Q (signal_3493) ) ;
    buf_clk cell_2307 ( .C (clk), .D (signal_3500), .Q (signal_3501) ) ;
    buf_clk cell_2315 ( .C (clk), .D (signal_3508), .Q (signal_3509) ) ;
    buf_clk cell_2323 ( .C (clk), .D (signal_3516), .Q (signal_3517) ) ;
    buf_clk cell_2331 ( .C (clk), .D (signal_3524), .Q (signal_3525) ) ;
    buf_clk cell_2339 ( .C (clk), .D (signal_3532), .Q (signal_3533) ) ;
    buf_clk cell_2347 ( .C (clk), .D (signal_3540), .Q (signal_3541) ) ;
    buf_clk cell_2355 ( .C (clk), .D (signal_3548), .Q (signal_3549) ) ;
    buf_clk cell_2363 ( .C (clk), .D (signal_3556), .Q (signal_3557) ) ;
    buf_clk cell_2371 ( .C (clk), .D (signal_3564), .Q (signal_3565) ) ;
    buf_clk cell_2379 ( .C (clk), .D (signal_3572), .Q (signal_3573) ) ;
    buf_clk cell_2387 ( .C (clk), .D (signal_3580), .Q (signal_3581) ) ;
    buf_clk cell_2395 ( .C (clk), .D (signal_3588), .Q (signal_3589) ) ;
    buf_clk cell_2403 ( .C (clk), .D (signal_3596), .Q (signal_3597) ) ;
    buf_clk cell_2411 ( .C (clk), .D (signal_3604), .Q (signal_3605) ) ;
    buf_clk cell_2419 ( .C (clk), .D (signal_3612), .Q (signal_3613) ) ;
    buf_clk cell_2427 ( .C (clk), .D (signal_3620), .Q (signal_3621) ) ;
    buf_clk cell_2435 ( .C (clk), .D (signal_3628), .Q (signal_3629) ) ;
    buf_clk cell_2443 ( .C (clk), .D (signal_3636), .Q (signal_3637) ) ;
    buf_clk cell_2451 ( .C (clk), .D (signal_3644), .Q (signal_3645) ) ;
    buf_clk cell_2459 ( .C (clk), .D (signal_3652), .Q (signal_3653) ) ;
    buf_clk cell_2467 ( .C (clk), .D (signal_3660), .Q (signal_3661) ) ;
    buf_clk cell_2475 ( .C (clk), .D (signal_3668), .Q (signal_3669) ) ;
    buf_clk cell_2483 ( .C (clk), .D (signal_3676), .Q (signal_3677) ) ;
    buf_clk cell_2491 ( .C (clk), .D (signal_3684), .Q (signal_3685) ) ;
    buf_clk cell_2499 ( .C (clk), .D (signal_3692), .Q (signal_3693) ) ;
    buf_clk cell_2507 ( .C (clk), .D (signal_3700), .Q (signal_3701) ) ;
    buf_clk cell_2515 ( .C (clk), .D (signal_3708), .Q (signal_3709) ) ;
    buf_clk cell_2523 ( .C (clk), .D (signal_3716), .Q (signal_3717) ) ;
    buf_clk cell_2531 ( .C (clk), .D (signal_3724), .Q (signal_3725) ) ;
    buf_clk cell_2539 ( .C (clk), .D (signal_3732), .Q (signal_3733) ) ;
    buf_clk cell_2547 ( .C (clk), .D (signal_3740), .Q (signal_3741) ) ;
    buf_clk cell_2555 ( .C (clk), .D (signal_3748), .Q (signal_3749) ) ;
    buf_clk cell_2563 ( .C (clk), .D (signal_3756), .Q (signal_3757) ) ;
    buf_clk cell_2571 ( .C (clk), .D (signal_3764), .Q (signal_3765) ) ;
    buf_clk cell_2579 ( .C (clk), .D (signal_3772), .Q (signal_3773) ) ;
    buf_clk cell_2587 ( .C (clk), .D (signal_3780), .Q (signal_3781) ) ;
    buf_clk cell_2595 ( .C (clk), .D (signal_3788), .Q (signal_3789) ) ;
    buf_clk cell_2603 ( .C (clk), .D (signal_3796), .Q (signal_3797) ) ;
    buf_clk cell_2611 ( .C (clk), .D (signal_3804), .Q (signal_3805) ) ;
    buf_clk cell_2619 ( .C (clk), .D (signal_3812), .Q (signal_3813) ) ;
    buf_clk cell_2627 ( .C (clk), .D (signal_3820), .Q (signal_3821) ) ;
    buf_clk cell_2635 ( .C (clk), .D (signal_3828), .Q (signal_3829) ) ;
    buf_clk cell_2643 ( .C (clk), .D (signal_3836), .Q (signal_3837) ) ;
    buf_clk cell_2651 ( .C (clk), .D (signal_3844), .Q (signal_3845) ) ;
    buf_clk cell_2659 ( .C (clk), .D (signal_3852), .Q (signal_3853) ) ;
    buf_clk cell_2667 ( .C (clk), .D (signal_3860), .Q (signal_3861) ) ;
    buf_clk cell_2675 ( .C (clk), .D (signal_3868), .Q (signal_3869) ) ;
    buf_clk cell_2683 ( .C (clk), .D (signal_3876), .Q (signal_3877) ) ;
    buf_clk cell_2691 ( .C (clk), .D (signal_3884), .Q (signal_3885) ) ;
    buf_clk cell_2699 ( .C (clk), .D (signal_3892), .Q (signal_3893) ) ;
    buf_clk cell_2707 ( .C (clk), .D (signal_3900), .Q (signal_3901) ) ;
    buf_clk cell_2715 ( .C (clk), .D (signal_3908), .Q (signal_3909) ) ;
    buf_clk cell_2723 ( .C (clk), .D (signal_3916), .Q (signal_3917) ) ;
    buf_clk cell_2731 ( .C (clk), .D (signal_3924), .Q (signal_3925) ) ;
    buf_clk cell_2739 ( .C (clk), .D (signal_3932), .Q (signal_3933) ) ;
    buf_clk cell_2747 ( .C (clk), .D (signal_3940), .Q (signal_3941) ) ;
    buf_clk cell_2755 ( .C (clk), .D (signal_3948), .Q (signal_3949) ) ;
    buf_clk cell_2763 ( .C (clk), .D (signal_3956), .Q (signal_3957) ) ;
    buf_clk cell_2771 ( .C (clk), .D (signal_3964), .Q (signal_3965) ) ;
    buf_clk cell_2779 ( .C (clk), .D (signal_3972), .Q (signal_3973) ) ;
    buf_clk cell_2787 ( .C (clk), .D (signal_3980), .Q (signal_3981) ) ;
    buf_clk cell_2795 ( .C (clk), .D (signal_3988), .Q (signal_3989) ) ;
    buf_clk cell_2803 ( .C (clk), .D (signal_3996), .Q (signal_3997) ) ;
    buf_clk cell_2811 ( .C (clk), .D (signal_4004), .Q (signal_4005) ) ;
    buf_clk cell_2819 ( .C (clk), .D (signal_4012), .Q (signal_4013) ) ;
    buf_clk cell_2827 ( .C (clk), .D (signal_4020), .Q (signal_4021) ) ;
    buf_clk cell_2835 ( .C (clk), .D (signal_4028), .Q (signal_4029) ) ;
    buf_clk cell_2843 ( .C (clk), .D (signal_4036), .Q (signal_4037) ) ;
    buf_clk cell_2851 ( .C (clk), .D (signal_4044), .Q (signal_4045) ) ;
    buf_clk cell_2859 ( .C (clk), .D (signal_4052), .Q (signal_4053) ) ;
    buf_clk cell_2867 ( .C (clk), .D (signal_4060), .Q (signal_4061) ) ;
    buf_clk cell_2875 ( .C (clk), .D (signal_4068), .Q (signal_4069) ) ;
    buf_clk cell_2883 ( .C (clk), .D (signal_4076), .Q (signal_4077) ) ;
    buf_clk cell_2891 ( .C (clk), .D (signal_4084), .Q (signal_4085) ) ;
    buf_clk cell_2899 ( .C (clk), .D (signal_4092), .Q (signal_4093) ) ;
    buf_clk cell_2907 ( .C (clk), .D (signal_4100), .Q (signal_4101) ) ;
    buf_clk cell_2915 ( .C (clk), .D (signal_4108), .Q (signal_4109) ) ;
    buf_clk cell_2923 ( .C (clk), .D (signal_4116), .Q (signal_4117) ) ;
    buf_clk cell_2931 ( .C (clk), .D (signal_4124), .Q (signal_4125) ) ;
    buf_clk cell_2939 ( .C (clk), .D (signal_4132), .Q (signal_4133) ) ;
    buf_clk cell_2947 ( .C (clk), .D (signal_4140), .Q (signal_4141) ) ;
    buf_clk cell_2955 ( .C (clk), .D (signal_4148), .Q (signal_4149) ) ;
    buf_clk cell_2963 ( .C (clk), .D (signal_4156), .Q (signal_4157) ) ;
    buf_clk cell_2971 ( .C (clk), .D (signal_4164), .Q (signal_4165) ) ;
    buf_clk cell_2979 ( .C (clk), .D (signal_4172), .Q (signal_4173) ) ;
    buf_clk cell_2987 ( .C (clk), .D (signal_4180), .Q (signal_4181) ) ;
    buf_clk cell_2995 ( .C (clk), .D (signal_4188), .Q (signal_4189) ) ;
    buf_clk cell_3003 ( .C (clk), .D (signal_4196), .Q (signal_4197) ) ;
    buf_clk cell_3011 ( .C (clk), .D (signal_4204), .Q (signal_4205) ) ;
    buf_clk cell_3019 ( .C (clk), .D (signal_4212), .Q (signal_4213) ) ;
    buf_clk cell_3027 ( .C (clk), .D (signal_4220), .Q (signal_4221) ) ;
    buf_clk cell_3035 ( .C (clk), .D (signal_4228), .Q (signal_4229) ) ;
    buf_clk cell_3043 ( .C (clk), .D (signal_4236), .Q (signal_4237) ) ;
    buf_clk cell_3051 ( .C (clk), .D (signal_4244), .Q (signal_4245) ) ;
    buf_clk cell_3059 ( .C (clk), .D (signal_4252), .Q (signal_4253) ) ;
    buf_clk cell_3067 ( .C (clk), .D (signal_4260), .Q (signal_4261) ) ;
    buf_clk cell_3075 ( .C (clk), .D (signal_4268), .Q (signal_4269) ) ;
    buf_clk cell_3083 ( .C (clk), .D (signal_4276), .Q (signal_4277) ) ;
    buf_clk cell_3091 ( .C (clk), .D (signal_4284), .Q (signal_4285) ) ;
    buf_clk cell_3099 ( .C (clk), .D (signal_4292), .Q (signal_4293) ) ;
    buf_clk cell_3107 ( .C (clk), .D (signal_4300), .Q (signal_4301) ) ;
    buf_clk cell_3115 ( .C (clk), .D (signal_4308), .Q (signal_4309) ) ;
    buf_clk cell_3123 ( .C (clk), .D (signal_4316), .Q (signal_4317) ) ;
    buf_clk cell_3131 ( .C (clk), .D (signal_4324), .Q (signal_4325) ) ;
    buf_clk cell_3139 ( .C (clk), .D (signal_4332), .Q (signal_4333) ) ;
    buf_clk cell_3147 ( .C (clk), .D (signal_4340), .Q (signal_4341) ) ;
    buf_clk cell_3155 ( .C (clk), .D (signal_4348), .Q (signal_4349) ) ;
    buf_clk cell_3163 ( .C (clk), .D (signal_4356), .Q (signal_4357) ) ;
    buf_clk cell_3491 ( .C (clk), .D (signal_4684), .Q (signal_4685) ) ;
    buf_clk cell_3499 ( .C (clk), .D (signal_4692), .Q (signal_4693) ) ;
    buf_clk cell_3507 ( .C (clk), .D (signal_4700), .Q (signal_4701) ) ;
    buf_clk cell_3515 ( .C (clk), .D (signal_4708), .Q (signal_4709) ) ;
    buf_clk cell_3523 ( .C (clk), .D (signal_4716), .Q (signal_4717) ) ;
    buf_clk cell_3531 ( .C (clk), .D (signal_4724), .Q (signal_4725) ) ;
    buf_clk cell_3539 ( .C (clk), .D (signal_4732), .Q (signal_4733) ) ;
    buf_clk cell_3547 ( .C (clk), .D (signal_4740), .Q (signal_4741) ) ;
    buf_clk cell_3555 ( .C (clk), .D (signal_4748), .Q (signal_4749) ) ;
    buf_clk cell_3563 ( .C (clk), .D (signal_4756), .Q (signal_4757) ) ;

    /* cells in depth 5 */
    buf_clk cell_1180 ( .C (clk), .D (signal_2373), .Q (signal_2374) ) ;
    buf_clk cell_1186 ( .C (clk), .D (signal_2379), .Q (signal_2380) ) ;
    buf_clk cell_1192 ( .C (clk), .D (signal_2385), .Q (signal_2386) ) ;
    buf_clk cell_1198 ( .C (clk), .D (signal_2391), .Q (signal_2392) ) ;
    buf_clk cell_1204 ( .C (clk), .D (signal_2397), .Q (signal_2398) ) ;
    buf_clk cell_1210 ( .C (clk), .D (signal_2403), .Q (signal_2404) ) ;
    buf_clk cell_1216 ( .C (clk), .D (signal_2409), .Q (signal_2410) ) ;
    buf_clk cell_1222 ( .C (clk), .D (signal_2415), .Q (signal_2416) ) ;
    buf_clk cell_1228 ( .C (clk), .D (signal_2421), .Q (signal_2422) ) ;
    buf_clk cell_1234 ( .C (clk), .D (signal_2427), .Q (signal_2428) ) ;
    buf_clk cell_1240 ( .C (clk), .D (signal_2433), .Q (signal_2434) ) ;
    buf_clk cell_1246 ( .C (clk), .D (signal_2439), .Q (signal_2440) ) ;
    buf_clk cell_1252 ( .C (clk), .D (signal_2445), .Q (signal_2446) ) ;
    buf_clk cell_1258 ( .C (clk), .D (signal_2451), .Q (signal_2452) ) ;
    buf_clk cell_1264 ( .C (clk), .D (signal_2457), .Q (signal_2458) ) ;
    buf_clk cell_1270 ( .C (clk), .D (signal_2463), .Q (signal_2464) ) ;
    buf_clk cell_1276 ( .C (clk), .D (signal_2469), .Q (signal_2470) ) ;
    buf_clk cell_1282 ( .C (clk), .D (signal_2475), .Q (signal_2476) ) ;
    buf_clk cell_1288 ( .C (clk), .D (signal_2481), .Q (signal_2482) ) ;
    buf_clk cell_1294 ( .C (clk), .D (signal_2487), .Q (signal_2488) ) ;
    buf_clk cell_1300 ( .C (clk), .D (signal_2493), .Q (signal_2494) ) ;
    buf_clk cell_1306 ( .C (clk), .D (signal_2499), .Q (signal_2500) ) ;
    buf_clk cell_1312 ( .C (clk), .D (signal_2505), .Q (signal_2506) ) ;
    buf_clk cell_1318 ( .C (clk), .D (signal_2511), .Q (signal_2512) ) ;
    buf_clk cell_1324 ( .C (clk), .D (signal_2517), .Q (signal_2518) ) ;
    buf_clk cell_1330 ( .C (clk), .D (signal_2523), .Q (signal_2524) ) ;
    buf_clk cell_1336 ( .C (clk), .D (signal_2529), .Q (signal_2530) ) ;
    buf_clk cell_1342 ( .C (clk), .D (signal_2535), .Q (signal_2536) ) ;
    buf_clk cell_1348 ( .C (clk), .D (signal_2541), .Q (signal_2542) ) ;
    buf_clk cell_1354 ( .C (clk), .D (signal_2547), .Q (signal_2548) ) ;
    buf_clk cell_1360 ( .C (clk), .D (signal_2553), .Q (signal_2554) ) ;
    buf_clk cell_1366 ( .C (clk), .D (signal_2559), .Q (signal_2560) ) ;
    buf_clk cell_1372 ( .C (clk), .D (signal_2565), .Q (signal_2566) ) ;
    buf_clk cell_1378 ( .C (clk), .D (signal_2571), .Q (signal_2572) ) ;
    buf_clk cell_1384 ( .C (clk), .D (signal_2577), .Q (signal_2578) ) ;
    buf_clk cell_1390 ( .C (clk), .D (signal_2583), .Q (signal_2584) ) ;
    buf_clk cell_1396 ( .C (clk), .D (signal_2589), .Q (signal_2590) ) ;
    buf_clk cell_1402 ( .C (clk), .D (signal_2595), .Q (signal_2596) ) ;
    buf_clk cell_1408 ( .C (clk), .D (signal_2601), .Q (signal_2602) ) ;
    buf_clk cell_1414 ( .C (clk), .D (signal_2607), .Q (signal_2608) ) ;
    buf_clk cell_1420 ( .C (clk), .D (signal_2613), .Q (signal_2614) ) ;
    buf_clk cell_1426 ( .C (clk), .D (signal_2619), .Q (signal_2620) ) ;
    buf_clk cell_1432 ( .C (clk), .D (signal_2625), .Q (signal_2626) ) ;
    buf_clk cell_1438 ( .C (clk), .D (signal_2631), .Q (signal_2632) ) ;
    buf_clk cell_1444 ( .C (clk), .D (signal_2637), .Q (signal_2638) ) ;
    buf_clk cell_1450 ( .C (clk), .D (signal_2643), .Q (signal_2644) ) ;
    buf_clk cell_1456 ( .C (clk), .D (signal_2649), .Q (signal_2650) ) ;
    buf_clk cell_1462 ( .C (clk), .D (signal_2655), .Q (signal_2656) ) ;
    buf_clk cell_1468 ( .C (clk), .D (signal_2661), .Q (signal_2662) ) ;
    buf_clk cell_1474 ( .C (clk), .D (signal_2667), .Q (signal_2668) ) ;
    buf_clk cell_1480 ( .C (clk), .D (signal_2673), .Q (signal_2674) ) ;
    buf_clk cell_1486 ( .C (clk), .D (signal_2679), .Q (signal_2680) ) ;
    buf_clk cell_1492 ( .C (clk), .D (signal_2685), .Q (signal_2686) ) ;
    buf_clk cell_1498 ( .C (clk), .D (signal_2691), .Q (signal_2692) ) ;
    buf_clk cell_1504 ( .C (clk), .D (signal_2697), .Q (signal_2698) ) ;
    buf_clk cell_1510 ( .C (clk), .D (signal_2703), .Q (signal_2704) ) ;
    buf_clk cell_1516 ( .C (clk), .D (signal_2709), .Q (signal_2710) ) ;
    buf_clk cell_1522 ( .C (clk), .D (signal_2715), .Q (signal_2716) ) ;
    buf_clk cell_1528 ( .C (clk), .D (signal_2721), .Q (signal_2722) ) ;
    buf_clk cell_1534 ( .C (clk), .D (signal_2727), .Q (signal_2728) ) ;
    buf_clk cell_1540 ( .C (clk), .D (signal_2733), .Q (signal_2734) ) ;
    buf_clk cell_1546 ( .C (clk), .D (signal_2739), .Q (signal_2740) ) ;
    buf_clk cell_1552 ( .C (clk), .D (signal_2745), .Q (signal_2746) ) ;
    buf_clk cell_1558 ( .C (clk), .D (signal_2751), .Q (signal_2752) ) ;
    buf_clk cell_1564 ( .C (clk), .D (signal_2757), .Q (signal_2758) ) ;
    buf_clk cell_1570 ( .C (clk), .D (signal_2763), .Q (signal_2764) ) ;
    buf_clk cell_1576 ( .C (clk), .D (signal_2769), .Q (signal_2770) ) ;
    buf_clk cell_1582 ( .C (clk), .D (signal_2775), .Q (signal_2776) ) ;
    buf_clk cell_1588 ( .C (clk), .D (signal_2781), .Q (signal_2782) ) ;
    buf_clk cell_1594 ( .C (clk), .D (signal_2787), .Q (signal_2788) ) ;
    buf_clk cell_1600 ( .C (clk), .D (signal_2793), .Q (signal_2794) ) ;
    buf_clk cell_1606 ( .C (clk), .D (signal_2799), .Q (signal_2800) ) ;
    buf_clk cell_1612 ( .C (clk), .D (signal_2805), .Q (signal_2806) ) ;
    buf_clk cell_1618 ( .C (clk), .D (signal_2811), .Q (signal_2812) ) ;
    buf_clk cell_1624 ( .C (clk), .D (signal_2817), .Q (signal_2818) ) ;
    buf_clk cell_1630 ( .C (clk), .D (signal_2823), .Q (signal_2824) ) ;
    buf_clk cell_1636 ( .C (clk), .D (signal_2829), .Q (signal_2830) ) ;
    buf_clk cell_1642 ( .C (clk), .D (signal_2835), .Q (signal_2836) ) ;
    buf_clk cell_1648 ( .C (clk), .D (signal_2841), .Q (signal_2842) ) ;
    buf_clk cell_1654 ( .C (clk), .D (signal_2847), .Q (signal_2848) ) ;
    buf_clk cell_1660 ( .C (clk), .D (signal_2853), .Q (signal_2854) ) ;
    buf_clk cell_1666 ( .C (clk), .D (signal_2859), .Q (signal_2860) ) ;
    buf_clk cell_1672 ( .C (clk), .D (signal_2865), .Q (signal_2866) ) ;
    buf_clk cell_1678 ( .C (clk), .D (signal_2871), .Q (signal_2872) ) ;
    buf_clk cell_1684 ( .C (clk), .D (signal_2877), .Q (signal_2878) ) ;
    buf_clk cell_1690 ( .C (clk), .D (signal_2883), .Q (signal_2884) ) ;
    buf_clk cell_1696 ( .C (clk), .D (signal_2889), .Q (signal_2890) ) ;
    buf_clk cell_1702 ( .C (clk), .D (signal_2895), .Q (signal_2896) ) ;
    buf_clk cell_1708 ( .C (clk), .D (signal_2901), .Q (signal_2902) ) ;
    buf_clk cell_1714 ( .C (clk), .D (signal_2907), .Q (signal_2908) ) ;
    buf_clk cell_1720 ( .C (clk), .D (signal_2913), .Q (signal_2914) ) ;
    buf_clk cell_1726 ( .C (clk), .D (signal_2919), .Q (signal_2920) ) ;
    buf_clk cell_1732 ( .C (clk), .D (signal_2925), .Q (signal_2926) ) ;
    buf_clk cell_1738 ( .C (clk), .D (signal_2931), .Q (signal_2932) ) ;
    buf_clk cell_1744 ( .C (clk), .D (signal_2937), .Q (signal_2938) ) ;
    buf_clk cell_1750 ( .C (clk), .D (signal_2943), .Q (signal_2944) ) ;
    buf_clk cell_1756 ( .C (clk), .D (signal_2949), .Q (signal_2950) ) ;
    buf_clk cell_1762 ( .C (clk), .D (signal_2955), .Q (signal_2956) ) ;
    buf_clk cell_1768 ( .C (clk), .D (signal_2961), .Q (signal_2962) ) ;
    buf_clk cell_1774 ( .C (clk), .D (signal_2967), .Q (signal_2968) ) ;
    buf_clk cell_1780 ( .C (clk), .D (signal_2973), .Q (signal_2974) ) ;
    buf_clk cell_1786 ( .C (clk), .D (signal_2979), .Q (signal_2980) ) ;
    buf_clk cell_1792 ( .C (clk), .D (signal_2985), .Q (signal_2986) ) ;
    buf_clk cell_1798 ( .C (clk), .D (signal_2991), .Q (signal_2992) ) ;
    buf_clk cell_1804 ( .C (clk), .D (signal_2997), .Q (signal_2998) ) ;
    buf_clk cell_1810 ( .C (clk), .D (signal_3003), .Q (signal_3004) ) ;
    buf_clk cell_1816 ( .C (clk), .D (signal_3009), .Q (signal_3010) ) ;
    buf_clk cell_1822 ( .C (clk), .D (signal_3015), .Q (signal_3016) ) ;
    buf_clk cell_1828 ( .C (clk), .D (signal_3021), .Q (signal_3022) ) ;
    buf_clk cell_1834 ( .C (clk), .D (signal_3027), .Q (signal_3028) ) ;
    buf_clk cell_1840 ( .C (clk), .D (signal_3033), .Q (signal_3034) ) ;
    buf_clk cell_1846 ( .C (clk), .D (signal_3039), .Q (signal_3040) ) ;
    buf_clk cell_1852 ( .C (clk), .D (signal_3045), .Q (signal_3046) ) ;
    buf_clk cell_1858 ( .C (clk), .D (signal_3051), .Q (signal_3052) ) ;
    buf_clk cell_1864 ( .C (clk), .D (signal_3057), .Q (signal_3058) ) ;
    buf_clk cell_1870 ( .C (clk), .D (signal_3063), .Q (signal_3064) ) ;
    buf_clk cell_1876 ( .C (clk), .D (signal_3069), .Q (signal_3070) ) ;
    buf_clk cell_1882 ( .C (clk), .D (signal_3075), .Q (signal_3076) ) ;
    buf_clk cell_1888 ( .C (clk), .D (signal_3081), .Q (signal_3082) ) ;
    buf_clk cell_1894 ( .C (clk), .D (signal_3087), .Q (signal_3088) ) ;
    buf_clk cell_1900 ( .C (clk), .D (signal_3093), .Q (signal_3094) ) ;
    buf_clk cell_1906 ( .C (clk), .D (signal_3099), .Q (signal_3100) ) ;
    buf_clk cell_1912 ( .C (clk), .D (signal_3105), .Q (signal_3106) ) ;
    buf_clk cell_1918 ( .C (clk), .D (signal_3111), .Q (signal_3112) ) ;
    buf_clk cell_1924 ( .C (clk), .D (signal_3117), .Q (signal_3118) ) ;
    buf_clk cell_1930 ( .C (clk), .D (signal_3123), .Q (signal_3124) ) ;
    buf_clk cell_1936 ( .C (clk), .D (signal_3129), .Q (signal_3130) ) ;
    buf_clk cell_1942 ( .C (clk), .D (signal_3135), .Q (signal_3136) ) ;
    buf_clk cell_1948 ( .C (clk), .D (signal_3141), .Q (signal_3142) ) ;
    buf_clk cell_2148 ( .C (clk), .D (signal_3341), .Q (signal_3342) ) ;
    buf_clk cell_2156 ( .C (clk), .D (signal_3349), .Q (signal_3350) ) ;
    buf_clk cell_2164 ( .C (clk), .D (signal_3357), .Q (signal_3358) ) ;
    buf_clk cell_2172 ( .C (clk), .D (signal_3365), .Q (signal_3366) ) ;
    buf_clk cell_2180 ( .C (clk), .D (signal_3373), .Q (signal_3374) ) ;
    buf_clk cell_2188 ( .C (clk), .D (signal_3381), .Q (signal_3382) ) ;
    buf_clk cell_2196 ( .C (clk), .D (signal_3389), .Q (signal_3390) ) ;
    buf_clk cell_2204 ( .C (clk), .D (signal_3397), .Q (signal_3398) ) ;
    buf_clk cell_2212 ( .C (clk), .D (signal_3405), .Q (signal_3406) ) ;
    buf_clk cell_2220 ( .C (clk), .D (signal_3413), .Q (signal_3414) ) ;
    buf_clk cell_2228 ( .C (clk), .D (signal_3421), .Q (signal_3422) ) ;
    buf_clk cell_2236 ( .C (clk), .D (signal_3429), .Q (signal_3430) ) ;
    buf_clk cell_2244 ( .C (clk), .D (signal_3437), .Q (signal_3438) ) ;
    buf_clk cell_2252 ( .C (clk), .D (signal_3445), .Q (signal_3446) ) ;
    buf_clk cell_2260 ( .C (clk), .D (signal_3453), .Q (signal_3454) ) ;
    buf_clk cell_2268 ( .C (clk), .D (signal_3461), .Q (signal_3462) ) ;
    buf_clk cell_2276 ( .C (clk), .D (signal_3469), .Q (signal_3470) ) ;
    buf_clk cell_2284 ( .C (clk), .D (signal_3477), .Q (signal_3478) ) ;
    buf_clk cell_2292 ( .C (clk), .D (signal_3485), .Q (signal_3486) ) ;
    buf_clk cell_2300 ( .C (clk), .D (signal_3493), .Q (signal_3494) ) ;
    buf_clk cell_2308 ( .C (clk), .D (signal_3501), .Q (signal_3502) ) ;
    buf_clk cell_2316 ( .C (clk), .D (signal_3509), .Q (signal_3510) ) ;
    buf_clk cell_2324 ( .C (clk), .D (signal_3517), .Q (signal_3518) ) ;
    buf_clk cell_2332 ( .C (clk), .D (signal_3525), .Q (signal_3526) ) ;
    buf_clk cell_2340 ( .C (clk), .D (signal_3533), .Q (signal_3534) ) ;
    buf_clk cell_2348 ( .C (clk), .D (signal_3541), .Q (signal_3542) ) ;
    buf_clk cell_2356 ( .C (clk), .D (signal_3549), .Q (signal_3550) ) ;
    buf_clk cell_2364 ( .C (clk), .D (signal_3557), .Q (signal_3558) ) ;
    buf_clk cell_2372 ( .C (clk), .D (signal_3565), .Q (signal_3566) ) ;
    buf_clk cell_2380 ( .C (clk), .D (signal_3573), .Q (signal_3574) ) ;
    buf_clk cell_2388 ( .C (clk), .D (signal_3581), .Q (signal_3582) ) ;
    buf_clk cell_2396 ( .C (clk), .D (signal_3589), .Q (signal_3590) ) ;
    buf_clk cell_2404 ( .C (clk), .D (signal_3597), .Q (signal_3598) ) ;
    buf_clk cell_2412 ( .C (clk), .D (signal_3605), .Q (signal_3606) ) ;
    buf_clk cell_2420 ( .C (clk), .D (signal_3613), .Q (signal_3614) ) ;
    buf_clk cell_2428 ( .C (clk), .D (signal_3621), .Q (signal_3622) ) ;
    buf_clk cell_2436 ( .C (clk), .D (signal_3629), .Q (signal_3630) ) ;
    buf_clk cell_2444 ( .C (clk), .D (signal_3637), .Q (signal_3638) ) ;
    buf_clk cell_2452 ( .C (clk), .D (signal_3645), .Q (signal_3646) ) ;
    buf_clk cell_2460 ( .C (clk), .D (signal_3653), .Q (signal_3654) ) ;
    buf_clk cell_2468 ( .C (clk), .D (signal_3661), .Q (signal_3662) ) ;
    buf_clk cell_2476 ( .C (clk), .D (signal_3669), .Q (signal_3670) ) ;
    buf_clk cell_2484 ( .C (clk), .D (signal_3677), .Q (signal_3678) ) ;
    buf_clk cell_2492 ( .C (clk), .D (signal_3685), .Q (signal_3686) ) ;
    buf_clk cell_2500 ( .C (clk), .D (signal_3693), .Q (signal_3694) ) ;
    buf_clk cell_2508 ( .C (clk), .D (signal_3701), .Q (signal_3702) ) ;
    buf_clk cell_2516 ( .C (clk), .D (signal_3709), .Q (signal_3710) ) ;
    buf_clk cell_2524 ( .C (clk), .D (signal_3717), .Q (signal_3718) ) ;
    buf_clk cell_2532 ( .C (clk), .D (signal_3725), .Q (signal_3726) ) ;
    buf_clk cell_2540 ( .C (clk), .D (signal_3733), .Q (signal_3734) ) ;
    buf_clk cell_2548 ( .C (clk), .D (signal_3741), .Q (signal_3742) ) ;
    buf_clk cell_2556 ( .C (clk), .D (signal_3749), .Q (signal_3750) ) ;
    buf_clk cell_2564 ( .C (clk), .D (signal_3757), .Q (signal_3758) ) ;
    buf_clk cell_2572 ( .C (clk), .D (signal_3765), .Q (signal_3766) ) ;
    buf_clk cell_2580 ( .C (clk), .D (signal_3773), .Q (signal_3774) ) ;
    buf_clk cell_2588 ( .C (clk), .D (signal_3781), .Q (signal_3782) ) ;
    buf_clk cell_2596 ( .C (clk), .D (signal_3789), .Q (signal_3790) ) ;
    buf_clk cell_2604 ( .C (clk), .D (signal_3797), .Q (signal_3798) ) ;
    buf_clk cell_2612 ( .C (clk), .D (signal_3805), .Q (signal_3806) ) ;
    buf_clk cell_2620 ( .C (clk), .D (signal_3813), .Q (signal_3814) ) ;
    buf_clk cell_2628 ( .C (clk), .D (signal_3821), .Q (signal_3822) ) ;
    buf_clk cell_2636 ( .C (clk), .D (signal_3829), .Q (signal_3830) ) ;
    buf_clk cell_2644 ( .C (clk), .D (signal_3837), .Q (signal_3838) ) ;
    buf_clk cell_2652 ( .C (clk), .D (signal_3845), .Q (signal_3846) ) ;
    buf_clk cell_2660 ( .C (clk), .D (signal_3853), .Q (signal_3854) ) ;
    buf_clk cell_2668 ( .C (clk), .D (signal_3861), .Q (signal_3862) ) ;
    buf_clk cell_2676 ( .C (clk), .D (signal_3869), .Q (signal_3870) ) ;
    buf_clk cell_2684 ( .C (clk), .D (signal_3877), .Q (signal_3878) ) ;
    buf_clk cell_2692 ( .C (clk), .D (signal_3885), .Q (signal_3886) ) ;
    buf_clk cell_2700 ( .C (clk), .D (signal_3893), .Q (signal_3894) ) ;
    buf_clk cell_2708 ( .C (clk), .D (signal_3901), .Q (signal_3902) ) ;
    buf_clk cell_2716 ( .C (clk), .D (signal_3909), .Q (signal_3910) ) ;
    buf_clk cell_2724 ( .C (clk), .D (signal_3917), .Q (signal_3918) ) ;
    buf_clk cell_2732 ( .C (clk), .D (signal_3925), .Q (signal_3926) ) ;
    buf_clk cell_2740 ( .C (clk), .D (signal_3933), .Q (signal_3934) ) ;
    buf_clk cell_2748 ( .C (clk), .D (signal_3941), .Q (signal_3942) ) ;
    buf_clk cell_2756 ( .C (clk), .D (signal_3949), .Q (signal_3950) ) ;
    buf_clk cell_2764 ( .C (clk), .D (signal_3957), .Q (signal_3958) ) ;
    buf_clk cell_2772 ( .C (clk), .D (signal_3965), .Q (signal_3966) ) ;
    buf_clk cell_2780 ( .C (clk), .D (signal_3973), .Q (signal_3974) ) ;
    buf_clk cell_2788 ( .C (clk), .D (signal_3981), .Q (signal_3982) ) ;
    buf_clk cell_2796 ( .C (clk), .D (signal_3989), .Q (signal_3990) ) ;
    buf_clk cell_2804 ( .C (clk), .D (signal_3997), .Q (signal_3998) ) ;
    buf_clk cell_2812 ( .C (clk), .D (signal_4005), .Q (signal_4006) ) ;
    buf_clk cell_2820 ( .C (clk), .D (signal_4013), .Q (signal_4014) ) ;
    buf_clk cell_2828 ( .C (clk), .D (signal_4021), .Q (signal_4022) ) ;
    buf_clk cell_2836 ( .C (clk), .D (signal_4029), .Q (signal_4030) ) ;
    buf_clk cell_2844 ( .C (clk), .D (signal_4037), .Q (signal_4038) ) ;
    buf_clk cell_2852 ( .C (clk), .D (signal_4045), .Q (signal_4046) ) ;
    buf_clk cell_2860 ( .C (clk), .D (signal_4053), .Q (signal_4054) ) ;
    buf_clk cell_2868 ( .C (clk), .D (signal_4061), .Q (signal_4062) ) ;
    buf_clk cell_2876 ( .C (clk), .D (signal_4069), .Q (signal_4070) ) ;
    buf_clk cell_2884 ( .C (clk), .D (signal_4077), .Q (signal_4078) ) ;
    buf_clk cell_2892 ( .C (clk), .D (signal_4085), .Q (signal_4086) ) ;
    buf_clk cell_2900 ( .C (clk), .D (signal_4093), .Q (signal_4094) ) ;
    buf_clk cell_2908 ( .C (clk), .D (signal_4101), .Q (signal_4102) ) ;
    buf_clk cell_2916 ( .C (clk), .D (signal_4109), .Q (signal_4110) ) ;
    buf_clk cell_2924 ( .C (clk), .D (signal_4117), .Q (signal_4118) ) ;
    buf_clk cell_2932 ( .C (clk), .D (signal_4125), .Q (signal_4126) ) ;
    buf_clk cell_2940 ( .C (clk), .D (signal_4133), .Q (signal_4134) ) ;
    buf_clk cell_2948 ( .C (clk), .D (signal_4141), .Q (signal_4142) ) ;
    buf_clk cell_2956 ( .C (clk), .D (signal_4149), .Q (signal_4150) ) ;
    buf_clk cell_2964 ( .C (clk), .D (signal_4157), .Q (signal_4158) ) ;
    buf_clk cell_2972 ( .C (clk), .D (signal_4165), .Q (signal_4166) ) ;
    buf_clk cell_2980 ( .C (clk), .D (signal_4173), .Q (signal_4174) ) ;
    buf_clk cell_2988 ( .C (clk), .D (signal_4181), .Q (signal_4182) ) ;
    buf_clk cell_2996 ( .C (clk), .D (signal_4189), .Q (signal_4190) ) ;
    buf_clk cell_3004 ( .C (clk), .D (signal_4197), .Q (signal_4198) ) ;
    buf_clk cell_3012 ( .C (clk), .D (signal_4205), .Q (signal_4206) ) ;
    buf_clk cell_3020 ( .C (clk), .D (signal_4213), .Q (signal_4214) ) ;
    buf_clk cell_3028 ( .C (clk), .D (signal_4221), .Q (signal_4222) ) ;
    buf_clk cell_3036 ( .C (clk), .D (signal_4229), .Q (signal_4230) ) ;
    buf_clk cell_3044 ( .C (clk), .D (signal_4237), .Q (signal_4238) ) ;
    buf_clk cell_3052 ( .C (clk), .D (signal_4245), .Q (signal_4246) ) ;
    buf_clk cell_3060 ( .C (clk), .D (signal_4253), .Q (signal_4254) ) ;
    buf_clk cell_3068 ( .C (clk), .D (signal_4261), .Q (signal_4262) ) ;
    buf_clk cell_3076 ( .C (clk), .D (signal_4269), .Q (signal_4270) ) ;
    buf_clk cell_3084 ( .C (clk), .D (signal_4277), .Q (signal_4278) ) ;
    buf_clk cell_3092 ( .C (clk), .D (signal_4285), .Q (signal_4286) ) ;
    buf_clk cell_3100 ( .C (clk), .D (signal_4293), .Q (signal_4294) ) ;
    buf_clk cell_3108 ( .C (clk), .D (signal_4301), .Q (signal_4302) ) ;
    buf_clk cell_3116 ( .C (clk), .D (signal_4309), .Q (signal_4310) ) ;
    buf_clk cell_3124 ( .C (clk), .D (signal_4317), .Q (signal_4318) ) ;
    buf_clk cell_3132 ( .C (clk), .D (signal_4325), .Q (signal_4326) ) ;
    buf_clk cell_3140 ( .C (clk), .D (signal_4333), .Q (signal_4334) ) ;
    buf_clk cell_3148 ( .C (clk), .D (signal_4341), .Q (signal_4342) ) ;
    buf_clk cell_3156 ( .C (clk), .D (signal_4349), .Q (signal_4350) ) ;
    buf_clk cell_3164 ( .C (clk), .D (signal_4357), .Q (signal_4358) ) ;
    buf_clk cell_3168 ( .C (clk), .D (signal_3235), .Q (signal_4362) ) ;
    buf_clk cell_3170 ( .C (clk), .D (signal_3239), .Q (signal_4364) ) ;
    buf_clk cell_3172 ( .C (clk), .D (signal_1114), .Q (signal_4366) ) ;
    buf_clk cell_3174 ( .C (clk), .D (signal_1367), .Q (signal_4368) ) ;
    buf_clk cell_3176 ( .C (clk), .D (signal_3151), .Q (signal_4370) ) ;
    buf_clk cell_3178 ( .C (clk), .D (signal_3155), .Q (signal_4372) ) ;
    buf_clk cell_3180 ( .C (clk), .D (signal_1070), .Q (signal_4374) ) ;
    buf_clk cell_3182 ( .C (clk), .D (signal_1316), .Q (signal_4376) ) ;
    buf_clk cell_3184 ( .C (clk), .D (signal_3183), .Q (signal_4378) ) ;
    buf_clk cell_3186 ( .C (clk), .D (signal_3187), .Q (signal_4380) ) ;
    buf_clk cell_3188 ( .C (clk), .D (signal_1090), .Q (signal_4382) ) ;
    buf_clk cell_3190 ( .C (clk), .D (signal_1338), .Q (signal_4384) ) ;
    buf_clk cell_3192 ( .C (clk), .D (signal_3243), .Q (signal_4386) ) ;
    buf_clk cell_3194 ( .C (clk), .D (signal_3247), .Q (signal_4388) ) ;
    buf_clk cell_3196 ( .C (clk), .D (signal_1093), .Q (signal_4390) ) ;
    buf_clk cell_3198 ( .C (clk), .D (signal_1342), .Q (signal_4392) ) ;
    buf_clk cell_3200 ( .C (clk), .D (signal_1059), .Q (signal_4394) ) ;
    buf_clk cell_3202 ( .C (clk), .D (signal_1296), .Q (signal_4396) ) ;
    buf_clk cell_3204 ( .C (clk), .D (signal_1073), .Q (signal_4398) ) ;
    buf_clk cell_3206 ( .C (clk), .D (signal_1319), .Q (signal_4400) ) ;
    buf_clk cell_3208 ( .C (clk), .D (signal_3227), .Q (signal_4402) ) ;
    buf_clk cell_3210 ( .C (clk), .D (signal_3231), .Q (signal_4404) ) ;
    buf_clk cell_3212 ( .C (clk), .D (signal_1103), .Q (signal_4406) ) ;
    buf_clk cell_3214 ( .C (clk), .D (signal_1353), .Q (signal_4408) ) ;
    buf_clk cell_3216 ( .C (clk), .D (signal_1095), .Q (signal_4410) ) ;
    buf_clk cell_3218 ( .C (clk), .D (signal_1344), .Q (signal_4412) ) ;
    buf_clk cell_3220 ( .C (clk), .D (signal_3251), .Q (signal_4414) ) ;
    buf_clk cell_3222 ( .C (clk), .D (signal_3255), .Q (signal_4416) ) ;
    buf_clk cell_3224 ( .C (clk), .D (signal_1065), .Q (signal_4418) ) ;
    buf_clk cell_3226 ( .C (clk), .D (signal_1308), .Q (signal_4420) ) ;
    buf_clk cell_3228 ( .C (clk), .D (signal_1096), .Q (signal_4422) ) ;
    buf_clk cell_3230 ( .C (clk), .D (signal_1345), .Q (signal_4424) ) ;
    buf_clk cell_3232 ( .C (clk), .D (signal_3259), .Q (signal_4426) ) ;
    buf_clk cell_3234 ( .C (clk), .D (signal_3263), .Q (signal_4428) ) ;
    buf_clk cell_3236 ( .C (clk), .D (signal_1060), .Q (signal_4430) ) ;
    buf_clk cell_3238 ( .C (clk), .D (signal_1298), .Q (signal_4432) ) ;
    buf_clk cell_3240 ( .C (clk), .D (signal_3191), .Q (signal_4434) ) ;
    buf_clk cell_3242 ( .C (clk), .D (signal_3195), .Q (signal_4436) ) ;
    buf_clk cell_3244 ( .C (clk), .D (signal_1058), .Q (signal_4438) ) ;
    buf_clk cell_3246 ( .C (clk), .D (signal_1294), .Q (signal_4440) ) ;
    buf_clk cell_3248 ( .C (clk), .D (signal_3215), .Q (signal_4442) ) ;
    buf_clk cell_3250 ( .C (clk), .D (signal_3219), .Q (signal_4444) ) ;
    buf_clk cell_3252 ( .C (clk), .D (signal_1089), .Q (signal_4446) ) ;
    buf_clk cell_3254 ( .C (clk), .D (signal_1337), .Q (signal_4448) ) ;
    buf_clk cell_3256 ( .C (clk), .D (signal_3207), .Q (signal_4450) ) ;
    buf_clk cell_3258 ( .C (clk), .D (signal_3211), .Q (signal_4452) ) ;
    buf_clk cell_3260 ( .C (clk), .D (signal_1106), .Q (signal_4454) ) ;
    buf_clk cell_3262 ( .C (clk), .D (signal_1357), .Q (signal_4456) ) ;
    buf_clk cell_3264 ( .C (clk), .D (signal_1071), .Q (signal_4458) ) ;
    buf_clk cell_3266 ( .C (clk), .D (signal_1317), .Q (signal_4460) ) ;
    buf_clk cell_3268 ( .C (clk), .D (signal_1063), .Q (signal_4462) ) ;
    buf_clk cell_3270 ( .C (clk), .D (signal_1304), .Q (signal_4464) ) ;
    buf_clk cell_3272 ( .C (clk), .D (signal_1080), .Q (signal_4466) ) ;
    buf_clk cell_3274 ( .C (clk), .D (signal_1327), .Q (signal_4468) ) ;
    buf_clk cell_3276 ( .C (clk), .D (signal_1074), .Q (signal_4470) ) ;
    buf_clk cell_3278 ( .C (clk), .D (signal_1320), .Q (signal_4472) ) ;
    buf_clk cell_3280 ( .C (clk), .D (signal_1067), .Q (signal_4474) ) ;
    buf_clk cell_3282 ( .C (clk), .D (signal_1312), .Q (signal_4476) ) ;
    buf_clk cell_3284 ( .C (clk), .D (signal_1109), .Q (signal_4478) ) ;
    buf_clk cell_3286 ( .C (clk), .D (signal_1361), .Q (signal_4480) ) ;
    buf_clk cell_3288 ( .C (clk), .D (signal_3271), .Q (signal_4482) ) ;
    buf_clk cell_3290 ( .C (clk), .D (signal_3275), .Q (signal_4484) ) ;
    buf_clk cell_3292 ( .C (clk), .D (signal_1116), .Q (signal_4486) ) ;
    buf_clk cell_3294 ( .C (clk), .D (signal_1370), .Q (signal_4488) ) ;
    buf_clk cell_3296 ( .C (clk), .D (signal_1121), .Q (signal_4490) ) ;
    buf_clk cell_3298 ( .C (clk), .D (signal_1376), .Q (signal_4492) ) ;
    buf_clk cell_3300 ( .C (clk), .D (signal_3283), .Q (signal_4494) ) ;
    buf_clk cell_3302 ( .C (clk), .D (signal_3287), .Q (signal_4496) ) ;
    buf_clk cell_3304 ( .C (clk), .D (signal_1122), .Q (signal_4498) ) ;
    buf_clk cell_3306 ( .C (clk), .D (signal_1377), .Q (signal_4500) ) ;
    buf_clk cell_3308 ( .C (clk), .D (signal_1127), .Q (signal_4502) ) ;
    buf_clk cell_3310 ( .C (clk), .D (signal_1383), .Q (signal_4504) ) ;
    buf_clk cell_3312 ( .C (clk), .D (signal_3295), .Q (signal_4506) ) ;
    buf_clk cell_3314 ( .C (clk), .D (signal_3299), .Q (signal_4508) ) ;
    buf_clk cell_3316 ( .C (clk), .D (signal_1128), .Q (signal_4510) ) ;
    buf_clk cell_3318 ( .C (clk), .D (signal_1384), .Q (signal_4512) ) ;
    buf_clk cell_3320 ( .C (clk), .D (signal_1133), .Q (signal_4514) ) ;
    buf_clk cell_3322 ( .C (clk), .D (signal_1390), .Q (signal_4516) ) ;
    buf_clk cell_3324 ( .C (clk), .D (signal_3307), .Q (signal_4518) ) ;
    buf_clk cell_3326 ( .C (clk), .D (signal_3311), .Q (signal_4520) ) ;
    buf_clk cell_3328 ( .C (clk), .D (signal_1134), .Q (signal_4522) ) ;
    buf_clk cell_3330 ( .C (clk), .D (signal_1391), .Q (signal_4524) ) ;
    buf_clk cell_3332 ( .C (clk), .D (signal_1139), .Q (signal_4526) ) ;
    buf_clk cell_3334 ( .C (clk), .D (signal_1397), .Q (signal_4528) ) ;
    buf_clk cell_3336 ( .C (clk), .D (signal_3319), .Q (signal_4530) ) ;
    buf_clk cell_3338 ( .C (clk), .D (signal_3323), .Q (signal_4532) ) ;
    buf_clk cell_3340 ( .C (clk), .D (signal_1140), .Q (signal_4534) ) ;
    buf_clk cell_3342 ( .C (clk), .D (signal_1398), .Q (signal_4536) ) ;
    buf_clk cell_3344 ( .C (clk), .D (signal_1145), .Q (signal_4538) ) ;
    buf_clk cell_3346 ( .C (clk), .D (signal_1404), .Q (signal_4540) ) ;
    buf_clk cell_3348 ( .C (clk), .D (signal_3331), .Q (signal_4542) ) ;
    buf_clk cell_3350 ( .C (clk), .D (signal_3335), .Q (signal_4544) ) ;
    buf_clk cell_3352 ( .C (clk), .D (signal_1146), .Q (signal_4546) ) ;
    buf_clk cell_3354 ( .C (clk), .D (signal_1406), .Q (signal_4548) ) ;
    buf_clk cell_3356 ( .C (clk), .D (signal_1151), .Q (signal_4550) ) ;
    buf_clk cell_3358 ( .C (clk), .D (signal_1412), .Q (signal_4552) ) ;
    buf_clk cell_3492 ( .C (clk), .D (signal_4685), .Q (signal_4686) ) ;
    buf_clk cell_3500 ( .C (clk), .D (signal_4693), .Q (signal_4694) ) ;
    buf_clk cell_3508 ( .C (clk), .D (signal_4701), .Q (signal_4702) ) ;
    buf_clk cell_3516 ( .C (clk), .D (signal_4709), .Q (signal_4710) ) ;
    buf_clk cell_3524 ( .C (clk), .D (signal_4717), .Q (signal_4718) ) ;
    buf_clk cell_3532 ( .C (clk), .D (signal_4725), .Q (signal_4726) ) ;
    buf_clk cell_3540 ( .C (clk), .D (signal_4733), .Q (signal_4734) ) ;
    buf_clk cell_3548 ( .C (clk), .D (signal_4741), .Q (signal_4742) ) ;
    buf_clk cell_3556 ( .C (clk), .D (signal_4749), .Q (signal_4750) ) ;
    buf_clk cell_3564 ( .C (clk), .D (signal_4757), .Q (signal_4758) ) ;

    /* cells in depth 6 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_1 ( .s (signal_2375), .b ({signal_1418, signal_773}), .a ({signal_2387, signal_2381}), .c ({signal_1494, signal_869}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_3 ( .s (signal_2375), .b ({signal_1443, signal_771}), .a ({signal_2399, signal_2393}), .c ({signal_1496, signal_867}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_5 ( .s (signal_2375), .b ({signal_1420, signal_769}), .a ({signal_2411, signal_2405}), .c ({signal_1498, signal_865}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_7 ( .s (signal_2375), .b ({signal_1457, signal_767}), .a ({signal_2423, signal_2417}), .c ({signal_1500, signal_863}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_9 ( .s (signal_2375), .b ({signal_1460, signal_765}), .a ({signal_2435, signal_2429}), .c ({signal_1502, signal_861}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_11 ( .s (signal_2375), .b ({signal_1429, signal_763}), .a ({signal_2447, signal_2441}), .c ({signal_1504, signal_859}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_13 ( .s (signal_2375), .b ({signal_1440, signal_761}), .a ({signal_2459, signal_2453}), .c ({signal_1506, signal_857}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_15 ( .s (signal_2375), .b ({signal_1453, signal_759}), .a ({signal_2471, signal_2465}), .c ({signal_1508, signal_855}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_17 ( .s (signal_2375), .b ({signal_1461, signal_757}), .a ({signal_2483, signal_2477}), .c ({signal_1510, signal_853}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_19 ( .s (signal_2375), .b ({signal_1447, signal_755}), .a ({signal_2495, signal_2489}), .c ({signal_1512, signal_851}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_21 ( .s (signal_2375), .b ({signal_1445, signal_753}), .a ({signal_2507, signal_2501}), .c ({signal_1514, signal_849}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_23 ( .s (signal_2375), .b ({signal_1415, signal_751}), .a ({signal_2519, signal_2513}), .c ({signal_1516, signal_847}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_25 ( .s (signal_2375), .b ({signal_1454, signal_749}), .a ({signal_2531, signal_2525}), .c ({signal_1518, signal_845}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_27 ( .s (signal_2375), .b ({signal_1451, signal_747}), .a ({signal_2543, signal_2537}), .c ({signal_1520, signal_843}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_29 ( .s (signal_2375), .b ({signal_1421, signal_745}), .a ({signal_2555, signal_2549}), .c ({signal_1522, signal_841}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_31 ( .s (signal_2375), .b ({signal_1427, signal_743}), .a ({signal_2567, signal_2561}), .c ({signal_1524, signal_839}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_33 ( .s (signal_2375), .b ({signal_1448, signal_741}), .a ({signal_2579, signal_2573}), .c ({signal_1526, signal_805}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_35 ( .s (signal_2375), .b ({signal_1434, signal_739}), .a ({signal_2591, signal_2585}), .c ({signal_1528, signal_803}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_37 ( .s (signal_2375), .b ({signal_1432, signal_737}), .a ({signal_2603, signal_2597}), .c ({signal_1530, signal_801}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_39 ( .s (signal_2375), .b ({signal_1439, signal_735}), .a ({signal_2615, signal_2609}), .c ({signal_1532, signal_799}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_41 ( .s (signal_2375), .b ({signal_1464, signal_733}), .a ({signal_2627, signal_2621}), .c ({signal_1534, signal_797}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_43 ( .s (signal_2375), .b ({signal_1467, signal_731}), .a ({signal_2639, signal_2633}), .c ({signal_1536, signal_795}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_45 ( .s (signal_2375), .b ({signal_1469, signal_729}), .a ({signal_2651, signal_2645}), .c ({signal_1538, signal_793}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_47 ( .s (signal_2375), .b ({signal_1472, signal_727}), .a ({signal_2663, signal_2657}), .c ({signal_1540, signal_791}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_49 ( .s (signal_2375), .b ({signal_1474, signal_725}), .a ({signal_2675, signal_2669}), .c ({signal_1542, signal_789}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_51 ( .s (signal_2375), .b ({signal_1477, signal_723}), .a ({signal_2687, signal_2681}), .c ({signal_1544, signal_787}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_53 ( .s (signal_2375), .b ({signal_1479, signal_721}), .a ({signal_2699, signal_2693}), .c ({signal_1546, signal_785}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_55 ( .s (signal_2375), .b ({signal_1482, signal_719}), .a ({signal_2711, signal_2705}), .c ({signal_1548, signal_783}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_57 ( .s (signal_2375), .b ({signal_1484, signal_717}), .a ({signal_2723, signal_2717}), .c ({signal_1550, signal_781}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_59 ( .s (signal_2375), .b ({signal_1487, signal_715}), .a ({signal_2735, signal_2729}), .c ({signal_1552, signal_779}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_61 ( .s (signal_2375), .b ({signal_1489, signal_713}), .a ({signal_2747, signal_2741}), .c ({signal_1554, signal_777}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_63 ( .s (signal_2375), .b ({signal_1492, signal_711}), .a ({signal_2759, signal_2753}), .c ({signal_1556, signal_775}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_69 ( .a ({signal_1798, signal_271}), .b ({signal_1797, signal_272}), .c ({signal_1848, signal_821}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_70 ( .a ({signal_1510, signal_853}), .b ({signal_1494, signal_869}), .c ({signal_1797, signal_272}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_71 ( .a ({1'b0, 1'b0}), .b ({signal_1542, signal_789}), .c ({signal_1798, signal_271}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_72 ( .a ({signal_1799, signal_273}), .b ({signal_1494, signal_869}), .c ({signal_1849, signal_837}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_73 ( .a ({1'b0, 1'b0}), .b ({signal_1526, signal_805}), .c ({signal_1799, signal_273}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_79 ( .a ({signal_1801, signal_277}), .b ({signal_1800, signal_278}), .c ({signal_1853, signal_819}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_80 ( .a ({signal_1512, signal_851}), .b ({signal_1496, signal_867}), .c ({signal_1800, signal_278}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_81 ( .a ({1'b0, 1'b0}), .b ({signal_1544, signal_787}), .c ({signal_1801, signal_277}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_82 ( .a ({signal_1802, signal_279}), .b ({signal_1496, signal_867}), .c ({signal_1854, signal_835}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_83 ( .a ({1'b0, 1'b0}), .b ({signal_1528, signal_803}), .c ({signal_1802, signal_279}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_89 ( .a ({signal_1804, signal_283}), .b ({signal_1803, signal_284}), .c ({signal_1858, signal_817}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_90 ( .a ({signal_1514, signal_849}), .b ({signal_1498, signal_865}), .c ({signal_1803, signal_284}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_91 ( .a ({1'b0, 1'b0}), .b ({signal_1546, signal_785}), .c ({signal_1804, signal_283}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_92 ( .a ({signal_1805, signal_285}), .b ({signal_1498, signal_865}), .c ({signal_1859, signal_833}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_93 ( .a ({1'b0, 1'b0}), .b ({signal_1530, signal_801}), .c ({signal_1805, signal_285}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_99 ( .a ({signal_1807, signal_289}), .b ({signal_1806, signal_290}), .c ({signal_1863, signal_815}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_100 ( .a ({signal_1516, signal_847}), .b ({signal_1500, signal_863}), .c ({signal_1806, signal_290}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_101 ( .a ({1'b0, 1'b0}), .b ({signal_1548, signal_783}), .c ({signal_1807, signal_289}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_102 ( .a ({signal_1808, signal_291}), .b ({signal_1500, signal_863}), .c ({signal_1864, signal_831}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_103 ( .a ({1'b0, 1'b0}), .b ({signal_1532, signal_799}), .c ({signal_1808, signal_291}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_109 ( .a ({signal_1810, signal_295}), .b ({signal_1809, signal_296}), .c ({signal_1868, signal_813}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_110 ( .a ({signal_1518, signal_845}), .b ({signal_1502, signal_861}), .c ({signal_1809, signal_296}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_111 ( .a ({1'b0, 1'b0}), .b ({signal_1550, signal_781}), .c ({signal_1810, signal_295}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_112 ( .a ({signal_1811, signal_297}), .b ({signal_1502, signal_861}), .c ({signal_1869, signal_829}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_113 ( .a ({1'b0, 1'b0}), .b ({signal_1534, signal_797}), .c ({signal_1811, signal_297}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_119 ( .a ({signal_1813, signal_301}), .b ({signal_1812, signal_302}), .c ({signal_1873, signal_811}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_120 ( .a ({signal_1520, signal_843}), .b ({signal_1504, signal_859}), .c ({signal_1812, signal_302}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_121 ( .a ({1'b0, 1'b0}), .b ({signal_1552, signal_779}), .c ({signal_1813, signal_301}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_122 ( .a ({signal_1814, signal_303}), .b ({signal_1504, signal_859}), .c ({signal_1874, signal_827}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_123 ( .a ({1'b0, 1'b0}), .b ({signal_1536, signal_795}), .c ({signal_1814, signal_303}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_129 ( .a ({signal_1816, signal_307}), .b ({signal_1815, signal_308}), .c ({signal_1878, signal_809}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_130 ( .a ({signal_1522, signal_841}), .b ({signal_1506, signal_857}), .c ({signal_1815, signal_308}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_131 ( .a ({1'b0, 1'b0}), .b ({signal_1554, signal_777}), .c ({signal_1816, signal_307}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_132 ( .a ({signal_1817, signal_309}), .b ({signal_1506, signal_857}), .c ({signal_1879, signal_825}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_133 ( .a ({1'b0, 1'b0}), .b ({signal_1538, signal_793}), .c ({signal_1817, signal_309}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_139 ( .a ({signal_1819, signal_313}), .b ({signal_1818, signal_314}), .c ({signal_1883, signal_807}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_140 ( .a ({signal_1524, signal_839}), .b ({signal_1508, signal_855}), .c ({signal_1818, signal_314}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_141 ( .a ({1'b0, 1'b0}), .b ({signal_1556, signal_775}), .c ({signal_1819, signal_313}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_142 ( .a ({signal_1820, signal_315}), .b ({signal_1508, signal_855}), .c ({signal_1884, signal_823}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_143 ( .a ({1'b0, 1'b0}), .b ({signal_1540, signal_791}), .c ({signal_1820, signal_315}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_146 ( .a ({signal_1933, signal_317}), .b ({signal_2771, signal_2765}), .c ({signal_1966, signal_949}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_147 ( .a ({1'b0, 1'b0}), .b ({signal_1848, signal_821}), .c ({signal_1933, signal_317}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_150 ( .a ({signal_1934, signal_319}), .b ({signal_2783, signal_2777}), .c ({signal_1968, signal_947}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_151 ( .a ({1'b0, 1'b0}), .b ({signal_1853, signal_819}), .c ({signal_1934, signal_319}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_154 ( .a ({signal_1935, signal_321}), .b ({signal_2795, signal_2789}), .c ({signal_1970, signal_945}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_155 ( .a ({1'b0, 1'b0}), .b ({signal_1858, signal_817}), .c ({signal_1935, signal_321}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_158 ( .a ({signal_1936, signal_323}), .b ({signal_2807, signal_2801}), .c ({signal_1972, signal_943}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_159 ( .a ({1'b0, 1'b0}), .b ({signal_1863, signal_815}), .c ({signal_1936, signal_323}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_162 ( .a ({signal_1937, signal_325}), .b ({signal_2819, signal_2813}), .c ({signal_1974, signal_941}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_163 ( .a ({1'b0, 1'b0}), .b ({signal_1868, signal_813}), .c ({signal_1937, signal_325}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_166 ( .a ({signal_1938, signal_327}), .b ({signal_2831, signal_2825}), .c ({signal_1976, signal_939}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_167 ( .a ({1'b0, 1'b0}), .b ({signal_1873, signal_811}), .c ({signal_1938, signal_327}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_170 ( .a ({signal_1939, signal_329}), .b ({signal_2843, signal_2837}), .c ({signal_1978, signal_937}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_171 ( .a ({1'b0, 1'b0}), .b ({signal_1878, signal_809}), .c ({signal_1939, signal_329}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_174 ( .a ({signal_1940, signal_331}), .b ({signal_2855, signal_2849}), .c ({signal_1980, signal_935}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_175 ( .a ({1'b0, 1'b0}), .b ({signal_1883, signal_807}), .c ({signal_1940, signal_331}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_179 ( .a ({signal_1941, signal_334}), .b ({signal_2867, signal_2861}), .c ({signal_1982, signal_957}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_181 ( .a ({1'b0, 1'b0}), .b ({signal_1869, signal_829}), .c ({signal_1941, signal_334}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_185 ( .a ({signal_1942, signal_338}), .b ({signal_2879, signal_2873}), .c ({signal_1984, signal_955}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_187 ( .a ({1'b0, 1'b0}), .b ({signal_1874, signal_827}), .c ({signal_1942, signal_338}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_191 ( .a ({signal_1943, signal_342}), .b ({signal_2891, signal_2885}), .c ({signal_1986, signal_953}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_193 ( .a ({1'b0, 1'b0}), .b ({signal_1879, signal_825}), .c ({signal_1943, signal_342}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_197 ( .a ({signal_1944, signal_346}), .b ({signal_2903, signal_2897}), .c ({signal_1988, signal_951}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_199 ( .a ({1'b0, 1'b0}), .b ({signal_1884, signal_823}), .c ({signal_1944, signal_346}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_202 ( .a ({signal_1829, signal_349}), .b ({signal_2915, signal_2909}), .c ({signal_1886, signal_997}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_203 ( .a ({1'b0, 1'b0}), .b ({signal_1494, signal_869}), .c ({signal_1829, signal_349}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_206 ( .a ({signal_1830, signal_351}), .b ({signal_2927, signal_2921}), .c ({signal_1888, signal_995}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_207 ( .a ({1'b0, 1'b0}), .b ({signal_1496, signal_867}), .c ({signal_1830, signal_351}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_210 ( .a ({signal_1831, signal_353}), .b ({signal_2939, signal_2933}), .c ({signal_1890, signal_993}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_211 ( .a ({1'b0, 1'b0}), .b ({signal_1498, signal_865}), .c ({signal_1831, signal_353}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_214 ( .a ({signal_1832, signal_355}), .b ({signal_2951, signal_2945}), .c ({signal_1892, signal_991}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_215 ( .a ({1'b0, 1'b0}), .b ({signal_1500, signal_863}), .c ({signal_1832, signal_355}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_218 ( .a ({signal_1833, signal_357}), .b ({signal_2963, signal_2957}), .c ({signal_1894, signal_989}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_219 ( .a ({1'b0, 1'b0}), .b ({signal_1502, signal_861}), .c ({signal_1833, signal_357}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_222 ( .a ({signal_1834, signal_359}), .b ({signal_2975, signal_2969}), .c ({signal_1896, signal_987}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_223 ( .a ({1'b0, 1'b0}), .b ({signal_1504, signal_859}), .c ({signal_1834, signal_359}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_226 ( .a ({signal_1835, signal_361}), .b ({signal_2987, signal_2981}), .c ({signal_1898, signal_985}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_227 ( .a ({1'b0, 1'b0}), .b ({signal_1506, signal_857}), .c ({signal_1835, signal_361}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_230 ( .a ({signal_1836, signal_363}), .b ({signal_2999, signal_2993}), .c ({signal_1900, signal_983}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_231 ( .a ({1'b0, 1'b0}), .b ({signal_1508, signal_855}), .c ({signal_1836, signal_363}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_234 ( .a ({signal_1837, signal_365}), .b ({signal_3011, signal_3005}), .c ({signal_1902, signal_981}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_235 ( .a ({1'b0, 1'b0}), .b ({signal_1510, signal_853}), .c ({signal_1837, signal_365}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_238 ( .a ({signal_1838, signal_367}), .b ({signal_3023, signal_3017}), .c ({signal_1904, signal_979}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_239 ( .a ({1'b0, 1'b0}), .b ({signal_1512, signal_851}), .c ({signal_1838, signal_367}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_242 ( .a ({signal_1839, signal_369}), .b ({signal_3035, signal_3029}), .c ({signal_1906, signal_977}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_243 ( .a ({1'b0, 1'b0}), .b ({signal_1514, signal_849}), .c ({signal_1839, signal_369}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_246 ( .a ({signal_1840, signal_371}), .b ({signal_3047, signal_3041}), .c ({signal_1908, signal_975}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_247 ( .a ({1'b0, 1'b0}), .b ({signal_1516, signal_847}), .c ({signal_1840, signal_371}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_250 ( .a ({signal_1841, signal_373}), .b ({signal_3059, signal_3053}), .c ({signal_1910, signal_973}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_251 ( .a ({1'b0, 1'b0}), .b ({signal_1518, signal_845}), .c ({signal_1841, signal_373}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_254 ( .a ({signal_1842, signal_375}), .b ({signal_3071, signal_3065}), .c ({signal_1912, signal_971}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_255 ( .a ({1'b0, 1'b0}), .b ({signal_1520, signal_843}), .c ({signal_1842, signal_375}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_258 ( .a ({signal_1843, signal_377}), .b ({signal_3083, signal_3077}), .c ({signal_1914, signal_969}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_259 ( .a ({1'b0, 1'b0}), .b ({signal_1522, signal_841}), .c ({signal_1843, signal_377}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_262 ( .a ({signal_1844, signal_379}), .b ({signal_3095, signal_3089}), .c ({signal_1916, signal_967}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_263 ( .a ({1'b0, 1'b0}), .b ({signal_1524, signal_839}), .c ({signal_1844, signal_379}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_266 ( .a ({signal_1961, signal_381}), .b ({signal_3107, signal_3101}), .c ({signal_1990, signal_965}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_267 ( .a ({1'b0, 1'b0}), .b ({signal_1849, signal_837}), .c ({signal_1961, signal_381}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_270 ( .a ({signal_1962, signal_383}), .b ({signal_3119, signal_3113}), .c ({signal_1992, signal_963}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_271 ( .a ({1'b0, 1'b0}), .b ({signal_1854, signal_835}), .c ({signal_1962, signal_383}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_274 ( .a ({signal_1963, signal_385}), .b ({signal_3131, signal_3125}), .c ({signal_1994, signal_961}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_275 ( .a ({1'b0, 1'b0}), .b ({signal_1859, signal_833}), .c ({signal_1963, signal_385}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_278 ( .a ({signal_1964, signal_387}), .b ({signal_3143, signal_3137}), .c ({signal_1996, signal_959}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_279 ( .a ({1'b0, 1'b0}), .b ({signal_1864, signal_831}), .c ({signal_1964, signal_387}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_952 ( .s ({signal_3147, signal_3145}), .b ({signal_1350, signal_1101}), .a ({signal_1302, signal_1062}), .clk (clk), .r (Fresh[133]), .c ({signal_1413, signal_1152}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_953 ( .s ({signal_3155, signal_3151}), .b ({signal_1316, signal_1070}), .a ({signal_1304, signal_1063}), .clk (clk), .r (Fresh[134]), .c ({signal_1415, signal_751}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_954 ( .s ({signal_3147, signal_3145}), .b ({1'b0, 1'b0}), .a ({signal_1347, signal_1098}), .clk (clk), .r (Fresh[135]), .c ({signal_1416, signal_1153}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_955 ( .s ({signal_3159, signal_3157}), .b ({1'b0, 1'b0}), .a ({signal_1368, signal_1115}), .clk (clk), .r (Fresh[136]), .c ({signal_1417, signal_1154}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_956 ( .s ({signal_3159, signal_3157}), .b ({signal_1322, signal_1076}), .a ({signal_1346, signal_1097}), .clk (clk), .r (Fresh[137]), .c ({signal_1418, signal_773}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_957 ( .s ({signal_3163, signal_3161}), .b ({1'b0, 1'b0}), .a ({signal_1349, signal_1100}), .clk (clk), .r (Fresh[138]), .c ({signal_1419, signal_1155}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_958 ( .s ({signal_3163, signal_3161}), .b ({signal_1330, signal_1083}), .a ({signal_1335, signal_1087}), .clk (clk), .r (Fresh[139]), .c ({signal_1420, signal_769}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_959 ( .s ({signal_3167, signal_3165}), .b ({signal_1351, signal_1102}), .a ({signal_1355, signal_1105}), .clk (clk), .r (Fresh[140]), .c ({signal_1421, signal_745}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_960 ( .s ({signal_3171, signal_3169}), .b ({1'b0, 1'b0}), .a ({signal_1362, signal_1110}), .clk (clk), .r (Fresh[141]), .c ({signal_1422, signal_1156}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_961 ( .s ({signal_3175, signal_3173}), .b ({signal_1348, signal_1099}), .a ({signal_1324, signal_1078}), .clk (clk), .r (Fresh[142]), .c ({signal_1423, signal_1157}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_962 ( .s ({signal_3167, signal_3165}), .b ({signal_1355, signal_1105}), .a ({signal_1334, signal_1086}), .clk (clk), .r (Fresh[143]), .c ({signal_1424, signal_1158}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_963 ( .s ({signal_3179, signal_3177}), .b ({1'b0, 1'b0}), .a ({signal_1340, signal_1092}), .clk (clk), .r (Fresh[144]), .c ({signal_1425, signal_1159}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_964 ( .s ({signal_3187, signal_3183}), .b ({signal_1338, signal_1090}), .a ({signal_1296, signal_1059}), .clk (clk), .r (Fresh[145]), .c ({signal_1427, signal_743}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_965 ( .s ({signal_3195, signal_3191}), .b ({signal_1312, signal_1067}), .a ({signal_1294, signal_1058}), .clk (clk), .r (Fresh[146]), .c ({signal_1429, signal_763}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_966 ( .s ({signal_3199, signal_3197}), .b ({1'b0, 1'b0}), .a ({signal_1339, signal_1091}), .clk (clk), .r (Fresh[147]), .c ({signal_1430, signal_1160}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_967 ( .s ({signal_3203, signal_3201}), .b ({1'b0, 1'b0}), .a ({signal_1323, signal_1077}), .clk (clk), .r (Fresh[148]), .c ({signal_1431, signal_1161}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_968 ( .s ({signal_3147, signal_3145}), .b ({signal_1313, signal_1068}), .a ({signal_1350, signal_1101}), .clk (clk), .r (Fresh[149]), .c ({signal_1432, signal_737}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_969 ( .s ({signal_3211, signal_3207}), .b ({signal_1317, signal_1071}), .a ({signal_1357, signal_1106}), .clk (clk), .r (Fresh[150]), .c ({signal_1434, signal_739}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_970 ( .s ({signal_3199, signal_3197}), .b ({signal_1300, signal_1061}), .a ({signal_1365, signal_1113}), .clk (clk), .r (Fresh[151]), .c ({signal_1435, signal_1162}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_971 ( .s ({signal_3179, signal_3177}), .b ({signal_1321, signal_1075}), .a ({signal_1328, signal_1081}), .clk (clk), .r (Fresh[152]), .c ({signal_1436, signal_1163}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_972 ( .s ({signal_3159, signal_3157}), .b ({signal_1346, signal_1097}), .a ({signal_1315, signal_1069}), .clk (clk), .r (Fresh[153]), .c ({signal_1437, signal_1164}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_973 ( .s ({signal_3219, signal_3215}), .b ({signal_1337, signal_1089}), .a ({signal_1361, signal_1109}), .clk (clk), .r (Fresh[154]), .c ({signal_1439, signal_735}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_974 ( .s ({signal_3223, signal_3221}), .b ({signal_1343, signal_1094}), .a ({signal_1329, signal_1082}), .clk (clk), .r (Fresh[155]), .c ({signal_1440, signal_761}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_975 ( .s ({signal_3163, signal_3161}), .b ({signal_1335, signal_1087}), .a ({signal_1363, signal_1111}), .clk (clk), .r (Fresh[156]), .c ({signal_1441, signal_1165}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_976 ( .s ({signal_3231, signal_3227}), .b ({signal_1344, signal_1095}), .a ({signal_1353, signal_1103}), .clk (clk), .r (Fresh[157]), .c ({signal_1443, signal_771}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_977 ( .s ({signal_3223, signal_3221}), .b ({1'b0, 1'b0}), .a ({signal_1333, signal_1085}), .clk (clk), .r (Fresh[158]), .c ({signal_1444, signal_1166}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_978 ( .s ({signal_3175, signal_3173}), .b ({signal_1310, signal_1066}), .a ({signal_1348, signal_1099}), .clk (clk), .r (Fresh[159]), .c ({signal_1445, signal_753}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_979 ( .s ({signal_3239, signal_3235}), .b ({signal_1319, signal_1073}), .a ({signal_1367, signal_1114}), .clk (clk), .r (Fresh[160]), .c ({signal_1447, signal_755}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_980 ( .s ({signal_3203, signal_3201}), .b ({signal_1292, signal_1057}), .a ({signal_1325, signal_1079}), .clk (clk), .r (Fresh[161]), .c ({signal_1448, signal_741}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_981 ( .s ({signal_3167, signal_3165}), .b ({1'b0, 1'b0}), .a ({signal_1332, signal_1084}), .clk (clk), .r (Fresh[162]), .c ({signal_1449, signal_1167}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_982 ( .s ({signal_3247, signal_3243}), .b ({signal_1345, signal_1096}), .a ({signal_1342, signal_1093}), .clk (clk), .r (Fresh[163]), .c ({signal_1451, signal_747}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_983 ( .s ({signal_3255, signal_3251}), .b ({signal_1320, signal_1074}), .a ({signal_1308, signal_1065}), .clk (clk), .r (Fresh[164]), .c ({signal_1453, signal_759}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_984 ( .s ({signal_3171, signal_3169}), .b ({signal_1336, signal_1088}), .a ({signal_1291, signal_1056}), .clk (clk), .r (Fresh[165]), .c ({signal_1454, signal_749}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_985 ( .s ({signal_3203, signal_3201}), .b ({signal_1325, signal_1079}), .a ({signal_1358, signal_1107}), .clk (clk), .r (Fresh[166]), .c ({signal_1455, signal_1168}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_986 ( .s ({signal_3263, signal_3259}), .b ({signal_1327, signal_1080}), .a ({signal_1298, signal_1060}), .clk (clk), .r (Fresh[167]), .c ({signal_1457, signal_767}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_987 ( .s ({signal_3175, signal_3173}), .b ({1'b0, 1'b0}), .a ({signal_1318, signal_1072}), .clk (clk), .r (Fresh[168]), .c ({signal_1458, signal_1169}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_988 ( .s ({signal_3223, signal_3221}), .b ({signal_1329, signal_1082}), .a ({signal_1306, signal_1064}), .clk (clk), .r (Fresh[169]), .c ({signal_1459, signal_1170}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_989 ( .s ({signal_3179, signal_3177}), .b ({signal_1364, signal_1112}), .a ({signal_1321, signal_1075}), .clk (clk), .r (Fresh[170]), .c ({signal_1460, signal_765}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_990 ( .s ({signal_3199, signal_3197}), .b ({signal_1359, signal_1108}), .a ({signal_1300, signal_1061}), .clk (clk), .r (Fresh[171]), .c ({signal_1461, signal_757}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_991 ( .s ({signal_3171, signal_3169}), .b ({signal_1291, signal_1056}), .a ({signal_1354, signal_1104}), .clk (clk), .r (Fresh[172]), .c ({signal_1462, signal_1171}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_992 ( .s ({signal_3267, signal_3265}), .b ({1'b0, 1'b0}), .a ({signal_1371, signal_1117}), .clk (clk), .r (Fresh[173]), .c ({signal_1463, signal_1172}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_993 ( .s ({signal_3267, signal_3265}), .b ({signal_1373, signal_1119}), .a ({signal_1372, signal_1118}), .clk (clk), .r (Fresh[174]), .c ({signal_1464, signal_733}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_994 ( .s ({signal_3267, signal_3265}), .b ({signal_1372, signal_1118}), .a ({signal_1374, signal_1120}), .clk (clk), .r (Fresh[175]), .c ({signal_1465, signal_1173}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_995 ( .s ({signal_3275, signal_3271}), .b ({signal_1370, signal_1116}), .a ({signal_1376, signal_1121}), .clk (clk), .r (Fresh[176]), .c ({signal_1467, signal_731}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_996 ( .s ({signal_3279, signal_3277}), .b ({1'b0, 1'b0}), .a ({signal_1378, signal_1123}), .clk (clk), .r (Fresh[177]), .c ({signal_1468, signal_1174}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_997 ( .s ({signal_3279, signal_3277}), .b ({signal_1380, signal_1125}), .a ({signal_1379, signal_1124}), .clk (clk), .r (Fresh[178]), .c ({signal_1469, signal_729}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_998 ( .s ({signal_3279, signal_3277}), .b ({signal_1379, signal_1124}), .a ({signal_1381, signal_1126}), .clk (clk), .r (Fresh[179]), .c ({signal_1470, signal_1175}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_999 ( .s ({signal_3287, signal_3283}), .b ({signal_1377, signal_1122}), .a ({signal_1383, signal_1127}), .clk (clk), .r (Fresh[180]), .c ({signal_1472, signal_727}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1000 ( .s ({signal_3291, signal_3289}), .b ({1'b0, 1'b0}), .a ({signal_1385, signal_1129}), .clk (clk), .r (Fresh[181]), .c ({signal_1473, signal_1176}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1001 ( .s ({signal_3291, signal_3289}), .b ({signal_1387, signal_1131}), .a ({signal_1386, signal_1130}), .clk (clk), .r (Fresh[182]), .c ({signal_1474, signal_725}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1002 ( .s ({signal_3291, signal_3289}), .b ({signal_1386, signal_1130}), .a ({signal_1388, signal_1132}), .clk (clk), .r (Fresh[183]), .c ({signal_1475, signal_1177}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1003 ( .s ({signal_3299, signal_3295}), .b ({signal_1384, signal_1128}), .a ({signal_1390, signal_1133}), .clk (clk), .r (Fresh[184]), .c ({signal_1477, signal_723}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1004 ( .s ({signal_3303, signal_3301}), .b ({1'b0, 1'b0}), .a ({signal_1392, signal_1135}), .clk (clk), .r (Fresh[185]), .c ({signal_1478, signal_1178}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1005 ( .s ({signal_3303, signal_3301}), .b ({signal_1394, signal_1137}), .a ({signal_1393, signal_1136}), .clk (clk), .r (Fresh[186]), .c ({signal_1479, signal_721}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1006 ( .s ({signal_3303, signal_3301}), .b ({signal_1393, signal_1136}), .a ({signal_1395, signal_1138}), .clk (clk), .r (Fresh[187]), .c ({signal_1480, signal_1179}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1007 ( .s ({signal_3311, signal_3307}), .b ({signal_1391, signal_1134}), .a ({signal_1397, signal_1139}), .clk (clk), .r (Fresh[188]), .c ({signal_1482, signal_719}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1008 ( .s ({signal_3315, signal_3313}), .b ({1'b0, 1'b0}), .a ({signal_1399, signal_1141}), .clk (clk), .r (Fresh[189]), .c ({signal_1483, signal_1180}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1009 ( .s ({signal_3315, signal_3313}), .b ({signal_1401, signal_1143}), .a ({signal_1400, signal_1142}), .clk (clk), .r (Fresh[190]), .c ({signal_1484, signal_717}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1010 ( .s ({signal_3315, signal_3313}), .b ({signal_1400, signal_1142}), .a ({signal_1402, signal_1144}), .clk (clk), .r (Fresh[191]), .c ({signal_1485, signal_1181}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1011 ( .s ({signal_3323, signal_3319}), .b ({signal_1398, signal_1140}), .a ({signal_1404, signal_1145}), .clk (clk), .r (Fresh[192]), .c ({signal_1487, signal_715}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1012 ( .s ({signal_3327, signal_3325}), .b ({1'b0, 1'b0}), .a ({signal_1407, signal_1147}), .clk (clk), .r (Fresh[193]), .c ({signal_1488, signal_1182}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1013 ( .s ({signal_3327, signal_3325}), .b ({signal_1409, signal_1149}), .a ({signal_1408, signal_1148}), .clk (clk), .r (Fresh[194]), .c ({signal_1489, signal_713}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1014 ( .s ({signal_3327, signal_3325}), .b ({signal_1408, signal_1148}), .a ({signal_1410, signal_1150}), .clk (clk), .r (Fresh[195]), .c ({signal_1490, signal_1183}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1015 ( .s ({signal_3335, signal_3331}), .b ({signal_1406, signal_1146}), .a ({signal_1412, signal_1151}), .clk (clk), .r (Fresh[196]), .c ({signal_1492, signal_711}) ) ;
    buf_clk cell_1181 ( .C (clk), .D (signal_2374), .Q (signal_2375) ) ;
    buf_clk cell_1187 ( .C (clk), .D (signal_2380), .Q (signal_2381) ) ;
    buf_clk cell_1193 ( .C (clk), .D (signal_2386), .Q (signal_2387) ) ;
    buf_clk cell_1199 ( .C (clk), .D (signal_2392), .Q (signal_2393) ) ;
    buf_clk cell_1205 ( .C (clk), .D (signal_2398), .Q (signal_2399) ) ;
    buf_clk cell_1211 ( .C (clk), .D (signal_2404), .Q (signal_2405) ) ;
    buf_clk cell_1217 ( .C (clk), .D (signal_2410), .Q (signal_2411) ) ;
    buf_clk cell_1223 ( .C (clk), .D (signal_2416), .Q (signal_2417) ) ;
    buf_clk cell_1229 ( .C (clk), .D (signal_2422), .Q (signal_2423) ) ;
    buf_clk cell_1235 ( .C (clk), .D (signal_2428), .Q (signal_2429) ) ;
    buf_clk cell_1241 ( .C (clk), .D (signal_2434), .Q (signal_2435) ) ;
    buf_clk cell_1247 ( .C (clk), .D (signal_2440), .Q (signal_2441) ) ;
    buf_clk cell_1253 ( .C (clk), .D (signal_2446), .Q (signal_2447) ) ;
    buf_clk cell_1259 ( .C (clk), .D (signal_2452), .Q (signal_2453) ) ;
    buf_clk cell_1265 ( .C (clk), .D (signal_2458), .Q (signal_2459) ) ;
    buf_clk cell_1271 ( .C (clk), .D (signal_2464), .Q (signal_2465) ) ;
    buf_clk cell_1277 ( .C (clk), .D (signal_2470), .Q (signal_2471) ) ;
    buf_clk cell_1283 ( .C (clk), .D (signal_2476), .Q (signal_2477) ) ;
    buf_clk cell_1289 ( .C (clk), .D (signal_2482), .Q (signal_2483) ) ;
    buf_clk cell_1295 ( .C (clk), .D (signal_2488), .Q (signal_2489) ) ;
    buf_clk cell_1301 ( .C (clk), .D (signal_2494), .Q (signal_2495) ) ;
    buf_clk cell_1307 ( .C (clk), .D (signal_2500), .Q (signal_2501) ) ;
    buf_clk cell_1313 ( .C (clk), .D (signal_2506), .Q (signal_2507) ) ;
    buf_clk cell_1319 ( .C (clk), .D (signal_2512), .Q (signal_2513) ) ;
    buf_clk cell_1325 ( .C (clk), .D (signal_2518), .Q (signal_2519) ) ;
    buf_clk cell_1331 ( .C (clk), .D (signal_2524), .Q (signal_2525) ) ;
    buf_clk cell_1337 ( .C (clk), .D (signal_2530), .Q (signal_2531) ) ;
    buf_clk cell_1343 ( .C (clk), .D (signal_2536), .Q (signal_2537) ) ;
    buf_clk cell_1349 ( .C (clk), .D (signal_2542), .Q (signal_2543) ) ;
    buf_clk cell_1355 ( .C (clk), .D (signal_2548), .Q (signal_2549) ) ;
    buf_clk cell_1361 ( .C (clk), .D (signal_2554), .Q (signal_2555) ) ;
    buf_clk cell_1367 ( .C (clk), .D (signal_2560), .Q (signal_2561) ) ;
    buf_clk cell_1373 ( .C (clk), .D (signal_2566), .Q (signal_2567) ) ;
    buf_clk cell_1379 ( .C (clk), .D (signal_2572), .Q (signal_2573) ) ;
    buf_clk cell_1385 ( .C (clk), .D (signal_2578), .Q (signal_2579) ) ;
    buf_clk cell_1391 ( .C (clk), .D (signal_2584), .Q (signal_2585) ) ;
    buf_clk cell_1397 ( .C (clk), .D (signal_2590), .Q (signal_2591) ) ;
    buf_clk cell_1403 ( .C (clk), .D (signal_2596), .Q (signal_2597) ) ;
    buf_clk cell_1409 ( .C (clk), .D (signal_2602), .Q (signal_2603) ) ;
    buf_clk cell_1415 ( .C (clk), .D (signal_2608), .Q (signal_2609) ) ;
    buf_clk cell_1421 ( .C (clk), .D (signal_2614), .Q (signal_2615) ) ;
    buf_clk cell_1427 ( .C (clk), .D (signal_2620), .Q (signal_2621) ) ;
    buf_clk cell_1433 ( .C (clk), .D (signal_2626), .Q (signal_2627) ) ;
    buf_clk cell_1439 ( .C (clk), .D (signal_2632), .Q (signal_2633) ) ;
    buf_clk cell_1445 ( .C (clk), .D (signal_2638), .Q (signal_2639) ) ;
    buf_clk cell_1451 ( .C (clk), .D (signal_2644), .Q (signal_2645) ) ;
    buf_clk cell_1457 ( .C (clk), .D (signal_2650), .Q (signal_2651) ) ;
    buf_clk cell_1463 ( .C (clk), .D (signal_2656), .Q (signal_2657) ) ;
    buf_clk cell_1469 ( .C (clk), .D (signal_2662), .Q (signal_2663) ) ;
    buf_clk cell_1475 ( .C (clk), .D (signal_2668), .Q (signal_2669) ) ;
    buf_clk cell_1481 ( .C (clk), .D (signal_2674), .Q (signal_2675) ) ;
    buf_clk cell_1487 ( .C (clk), .D (signal_2680), .Q (signal_2681) ) ;
    buf_clk cell_1493 ( .C (clk), .D (signal_2686), .Q (signal_2687) ) ;
    buf_clk cell_1499 ( .C (clk), .D (signal_2692), .Q (signal_2693) ) ;
    buf_clk cell_1505 ( .C (clk), .D (signal_2698), .Q (signal_2699) ) ;
    buf_clk cell_1511 ( .C (clk), .D (signal_2704), .Q (signal_2705) ) ;
    buf_clk cell_1517 ( .C (clk), .D (signal_2710), .Q (signal_2711) ) ;
    buf_clk cell_1523 ( .C (clk), .D (signal_2716), .Q (signal_2717) ) ;
    buf_clk cell_1529 ( .C (clk), .D (signal_2722), .Q (signal_2723) ) ;
    buf_clk cell_1535 ( .C (clk), .D (signal_2728), .Q (signal_2729) ) ;
    buf_clk cell_1541 ( .C (clk), .D (signal_2734), .Q (signal_2735) ) ;
    buf_clk cell_1547 ( .C (clk), .D (signal_2740), .Q (signal_2741) ) ;
    buf_clk cell_1553 ( .C (clk), .D (signal_2746), .Q (signal_2747) ) ;
    buf_clk cell_1559 ( .C (clk), .D (signal_2752), .Q (signal_2753) ) ;
    buf_clk cell_1565 ( .C (clk), .D (signal_2758), .Q (signal_2759) ) ;
    buf_clk cell_1571 ( .C (clk), .D (signal_2764), .Q (signal_2765) ) ;
    buf_clk cell_1577 ( .C (clk), .D (signal_2770), .Q (signal_2771) ) ;
    buf_clk cell_1583 ( .C (clk), .D (signal_2776), .Q (signal_2777) ) ;
    buf_clk cell_1589 ( .C (clk), .D (signal_2782), .Q (signal_2783) ) ;
    buf_clk cell_1595 ( .C (clk), .D (signal_2788), .Q (signal_2789) ) ;
    buf_clk cell_1601 ( .C (clk), .D (signal_2794), .Q (signal_2795) ) ;
    buf_clk cell_1607 ( .C (clk), .D (signal_2800), .Q (signal_2801) ) ;
    buf_clk cell_1613 ( .C (clk), .D (signal_2806), .Q (signal_2807) ) ;
    buf_clk cell_1619 ( .C (clk), .D (signal_2812), .Q (signal_2813) ) ;
    buf_clk cell_1625 ( .C (clk), .D (signal_2818), .Q (signal_2819) ) ;
    buf_clk cell_1631 ( .C (clk), .D (signal_2824), .Q (signal_2825) ) ;
    buf_clk cell_1637 ( .C (clk), .D (signal_2830), .Q (signal_2831) ) ;
    buf_clk cell_1643 ( .C (clk), .D (signal_2836), .Q (signal_2837) ) ;
    buf_clk cell_1649 ( .C (clk), .D (signal_2842), .Q (signal_2843) ) ;
    buf_clk cell_1655 ( .C (clk), .D (signal_2848), .Q (signal_2849) ) ;
    buf_clk cell_1661 ( .C (clk), .D (signal_2854), .Q (signal_2855) ) ;
    buf_clk cell_1667 ( .C (clk), .D (signal_2860), .Q (signal_2861) ) ;
    buf_clk cell_1673 ( .C (clk), .D (signal_2866), .Q (signal_2867) ) ;
    buf_clk cell_1679 ( .C (clk), .D (signal_2872), .Q (signal_2873) ) ;
    buf_clk cell_1685 ( .C (clk), .D (signal_2878), .Q (signal_2879) ) ;
    buf_clk cell_1691 ( .C (clk), .D (signal_2884), .Q (signal_2885) ) ;
    buf_clk cell_1697 ( .C (clk), .D (signal_2890), .Q (signal_2891) ) ;
    buf_clk cell_1703 ( .C (clk), .D (signal_2896), .Q (signal_2897) ) ;
    buf_clk cell_1709 ( .C (clk), .D (signal_2902), .Q (signal_2903) ) ;
    buf_clk cell_1715 ( .C (clk), .D (signal_2908), .Q (signal_2909) ) ;
    buf_clk cell_1721 ( .C (clk), .D (signal_2914), .Q (signal_2915) ) ;
    buf_clk cell_1727 ( .C (clk), .D (signal_2920), .Q (signal_2921) ) ;
    buf_clk cell_1733 ( .C (clk), .D (signal_2926), .Q (signal_2927) ) ;
    buf_clk cell_1739 ( .C (clk), .D (signal_2932), .Q (signal_2933) ) ;
    buf_clk cell_1745 ( .C (clk), .D (signal_2938), .Q (signal_2939) ) ;
    buf_clk cell_1751 ( .C (clk), .D (signal_2944), .Q (signal_2945) ) ;
    buf_clk cell_1757 ( .C (clk), .D (signal_2950), .Q (signal_2951) ) ;
    buf_clk cell_1763 ( .C (clk), .D (signal_2956), .Q (signal_2957) ) ;
    buf_clk cell_1769 ( .C (clk), .D (signal_2962), .Q (signal_2963) ) ;
    buf_clk cell_1775 ( .C (clk), .D (signal_2968), .Q (signal_2969) ) ;
    buf_clk cell_1781 ( .C (clk), .D (signal_2974), .Q (signal_2975) ) ;
    buf_clk cell_1787 ( .C (clk), .D (signal_2980), .Q (signal_2981) ) ;
    buf_clk cell_1793 ( .C (clk), .D (signal_2986), .Q (signal_2987) ) ;
    buf_clk cell_1799 ( .C (clk), .D (signal_2992), .Q (signal_2993) ) ;
    buf_clk cell_1805 ( .C (clk), .D (signal_2998), .Q (signal_2999) ) ;
    buf_clk cell_1811 ( .C (clk), .D (signal_3004), .Q (signal_3005) ) ;
    buf_clk cell_1817 ( .C (clk), .D (signal_3010), .Q (signal_3011) ) ;
    buf_clk cell_1823 ( .C (clk), .D (signal_3016), .Q (signal_3017) ) ;
    buf_clk cell_1829 ( .C (clk), .D (signal_3022), .Q (signal_3023) ) ;
    buf_clk cell_1835 ( .C (clk), .D (signal_3028), .Q (signal_3029) ) ;
    buf_clk cell_1841 ( .C (clk), .D (signal_3034), .Q (signal_3035) ) ;
    buf_clk cell_1847 ( .C (clk), .D (signal_3040), .Q (signal_3041) ) ;
    buf_clk cell_1853 ( .C (clk), .D (signal_3046), .Q (signal_3047) ) ;
    buf_clk cell_1859 ( .C (clk), .D (signal_3052), .Q (signal_3053) ) ;
    buf_clk cell_1865 ( .C (clk), .D (signal_3058), .Q (signal_3059) ) ;
    buf_clk cell_1871 ( .C (clk), .D (signal_3064), .Q (signal_3065) ) ;
    buf_clk cell_1877 ( .C (clk), .D (signal_3070), .Q (signal_3071) ) ;
    buf_clk cell_1883 ( .C (clk), .D (signal_3076), .Q (signal_3077) ) ;
    buf_clk cell_1889 ( .C (clk), .D (signal_3082), .Q (signal_3083) ) ;
    buf_clk cell_1895 ( .C (clk), .D (signal_3088), .Q (signal_3089) ) ;
    buf_clk cell_1901 ( .C (clk), .D (signal_3094), .Q (signal_3095) ) ;
    buf_clk cell_1907 ( .C (clk), .D (signal_3100), .Q (signal_3101) ) ;
    buf_clk cell_1913 ( .C (clk), .D (signal_3106), .Q (signal_3107) ) ;
    buf_clk cell_1919 ( .C (clk), .D (signal_3112), .Q (signal_3113) ) ;
    buf_clk cell_1925 ( .C (clk), .D (signal_3118), .Q (signal_3119) ) ;
    buf_clk cell_1931 ( .C (clk), .D (signal_3124), .Q (signal_3125) ) ;
    buf_clk cell_1937 ( .C (clk), .D (signal_3130), .Q (signal_3131) ) ;
    buf_clk cell_1943 ( .C (clk), .D (signal_3136), .Q (signal_3137) ) ;
    buf_clk cell_1949 ( .C (clk), .D (signal_3142), .Q (signal_3143) ) ;
    buf_clk cell_2149 ( .C (clk), .D (signal_3342), .Q (signal_3343) ) ;
    buf_clk cell_2157 ( .C (clk), .D (signal_3350), .Q (signal_3351) ) ;
    buf_clk cell_2165 ( .C (clk), .D (signal_3358), .Q (signal_3359) ) ;
    buf_clk cell_2173 ( .C (clk), .D (signal_3366), .Q (signal_3367) ) ;
    buf_clk cell_2181 ( .C (clk), .D (signal_3374), .Q (signal_3375) ) ;
    buf_clk cell_2189 ( .C (clk), .D (signal_3382), .Q (signal_3383) ) ;
    buf_clk cell_2197 ( .C (clk), .D (signal_3390), .Q (signal_3391) ) ;
    buf_clk cell_2205 ( .C (clk), .D (signal_3398), .Q (signal_3399) ) ;
    buf_clk cell_2213 ( .C (clk), .D (signal_3406), .Q (signal_3407) ) ;
    buf_clk cell_2221 ( .C (clk), .D (signal_3414), .Q (signal_3415) ) ;
    buf_clk cell_2229 ( .C (clk), .D (signal_3422), .Q (signal_3423) ) ;
    buf_clk cell_2237 ( .C (clk), .D (signal_3430), .Q (signal_3431) ) ;
    buf_clk cell_2245 ( .C (clk), .D (signal_3438), .Q (signal_3439) ) ;
    buf_clk cell_2253 ( .C (clk), .D (signal_3446), .Q (signal_3447) ) ;
    buf_clk cell_2261 ( .C (clk), .D (signal_3454), .Q (signal_3455) ) ;
    buf_clk cell_2269 ( .C (clk), .D (signal_3462), .Q (signal_3463) ) ;
    buf_clk cell_2277 ( .C (clk), .D (signal_3470), .Q (signal_3471) ) ;
    buf_clk cell_2285 ( .C (clk), .D (signal_3478), .Q (signal_3479) ) ;
    buf_clk cell_2293 ( .C (clk), .D (signal_3486), .Q (signal_3487) ) ;
    buf_clk cell_2301 ( .C (clk), .D (signal_3494), .Q (signal_3495) ) ;
    buf_clk cell_2309 ( .C (clk), .D (signal_3502), .Q (signal_3503) ) ;
    buf_clk cell_2317 ( .C (clk), .D (signal_3510), .Q (signal_3511) ) ;
    buf_clk cell_2325 ( .C (clk), .D (signal_3518), .Q (signal_3519) ) ;
    buf_clk cell_2333 ( .C (clk), .D (signal_3526), .Q (signal_3527) ) ;
    buf_clk cell_2341 ( .C (clk), .D (signal_3534), .Q (signal_3535) ) ;
    buf_clk cell_2349 ( .C (clk), .D (signal_3542), .Q (signal_3543) ) ;
    buf_clk cell_2357 ( .C (clk), .D (signal_3550), .Q (signal_3551) ) ;
    buf_clk cell_2365 ( .C (clk), .D (signal_3558), .Q (signal_3559) ) ;
    buf_clk cell_2373 ( .C (clk), .D (signal_3566), .Q (signal_3567) ) ;
    buf_clk cell_2381 ( .C (clk), .D (signal_3574), .Q (signal_3575) ) ;
    buf_clk cell_2389 ( .C (clk), .D (signal_3582), .Q (signal_3583) ) ;
    buf_clk cell_2397 ( .C (clk), .D (signal_3590), .Q (signal_3591) ) ;
    buf_clk cell_2405 ( .C (clk), .D (signal_3598), .Q (signal_3599) ) ;
    buf_clk cell_2413 ( .C (clk), .D (signal_3606), .Q (signal_3607) ) ;
    buf_clk cell_2421 ( .C (clk), .D (signal_3614), .Q (signal_3615) ) ;
    buf_clk cell_2429 ( .C (clk), .D (signal_3622), .Q (signal_3623) ) ;
    buf_clk cell_2437 ( .C (clk), .D (signal_3630), .Q (signal_3631) ) ;
    buf_clk cell_2445 ( .C (clk), .D (signal_3638), .Q (signal_3639) ) ;
    buf_clk cell_2453 ( .C (clk), .D (signal_3646), .Q (signal_3647) ) ;
    buf_clk cell_2461 ( .C (clk), .D (signal_3654), .Q (signal_3655) ) ;
    buf_clk cell_2469 ( .C (clk), .D (signal_3662), .Q (signal_3663) ) ;
    buf_clk cell_2477 ( .C (clk), .D (signal_3670), .Q (signal_3671) ) ;
    buf_clk cell_2485 ( .C (clk), .D (signal_3678), .Q (signal_3679) ) ;
    buf_clk cell_2493 ( .C (clk), .D (signal_3686), .Q (signal_3687) ) ;
    buf_clk cell_2501 ( .C (clk), .D (signal_3694), .Q (signal_3695) ) ;
    buf_clk cell_2509 ( .C (clk), .D (signal_3702), .Q (signal_3703) ) ;
    buf_clk cell_2517 ( .C (clk), .D (signal_3710), .Q (signal_3711) ) ;
    buf_clk cell_2525 ( .C (clk), .D (signal_3718), .Q (signal_3719) ) ;
    buf_clk cell_2533 ( .C (clk), .D (signal_3726), .Q (signal_3727) ) ;
    buf_clk cell_2541 ( .C (clk), .D (signal_3734), .Q (signal_3735) ) ;
    buf_clk cell_2549 ( .C (clk), .D (signal_3742), .Q (signal_3743) ) ;
    buf_clk cell_2557 ( .C (clk), .D (signal_3750), .Q (signal_3751) ) ;
    buf_clk cell_2565 ( .C (clk), .D (signal_3758), .Q (signal_3759) ) ;
    buf_clk cell_2573 ( .C (clk), .D (signal_3766), .Q (signal_3767) ) ;
    buf_clk cell_2581 ( .C (clk), .D (signal_3774), .Q (signal_3775) ) ;
    buf_clk cell_2589 ( .C (clk), .D (signal_3782), .Q (signal_3783) ) ;
    buf_clk cell_2597 ( .C (clk), .D (signal_3790), .Q (signal_3791) ) ;
    buf_clk cell_2605 ( .C (clk), .D (signal_3798), .Q (signal_3799) ) ;
    buf_clk cell_2613 ( .C (clk), .D (signal_3806), .Q (signal_3807) ) ;
    buf_clk cell_2621 ( .C (clk), .D (signal_3814), .Q (signal_3815) ) ;
    buf_clk cell_2629 ( .C (clk), .D (signal_3822), .Q (signal_3823) ) ;
    buf_clk cell_2637 ( .C (clk), .D (signal_3830), .Q (signal_3831) ) ;
    buf_clk cell_2645 ( .C (clk), .D (signal_3838), .Q (signal_3839) ) ;
    buf_clk cell_2653 ( .C (clk), .D (signal_3846), .Q (signal_3847) ) ;
    buf_clk cell_2661 ( .C (clk), .D (signal_3854), .Q (signal_3855) ) ;
    buf_clk cell_2669 ( .C (clk), .D (signal_3862), .Q (signal_3863) ) ;
    buf_clk cell_2677 ( .C (clk), .D (signal_3870), .Q (signal_3871) ) ;
    buf_clk cell_2685 ( .C (clk), .D (signal_3878), .Q (signal_3879) ) ;
    buf_clk cell_2693 ( .C (clk), .D (signal_3886), .Q (signal_3887) ) ;
    buf_clk cell_2701 ( .C (clk), .D (signal_3894), .Q (signal_3895) ) ;
    buf_clk cell_2709 ( .C (clk), .D (signal_3902), .Q (signal_3903) ) ;
    buf_clk cell_2717 ( .C (clk), .D (signal_3910), .Q (signal_3911) ) ;
    buf_clk cell_2725 ( .C (clk), .D (signal_3918), .Q (signal_3919) ) ;
    buf_clk cell_2733 ( .C (clk), .D (signal_3926), .Q (signal_3927) ) ;
    buf_clk cell_2741 ( .C (clk), .D (signal_3934), .Q (signal_3935) ) ;
    buf_clk cell_2749 ( .C (clk), .D (signal_3942), .Q (signal_3943) ) ;
    buf_clk cell_2757 ( .C (clk), .D (signal_3950), .Q (signal_3951) ) ;
    buf_clk cell_2765 ( .C (clk), .D (signal_3958), .Q (signal_3959) ) ;
    buf_clk cell_2773 ( .C (clk), .D (signal_3966), .Q (signal_3967) ) ;
    buf_clk cell_2781 ( .C (clk), .D (signal_3974), .Q (signal_3975) ) ;
    buf_clk cell_2789 ( .C (clk), .D (signal_3982), .Q (signal_3983) ) ;
    buf_clk cell_2797 ( .C (clk), .D (signal_3990), .Q (signal_3991) ) ;
    buf_clk cell_2805 ( .C (clk), .D (signal_3998), .Q (signal_3999) ) ;
    buf_clk cell_2813 ( .C (clk), .D (signal_4006), .Q (signal_4007) ) ;
    buf_clk cell_2821 ( .C (clk), .D (signal_4014), .Q (signal_4015) ) ;
    buf_clk cell_2829 ( .C (clk), .D (signal_4022), .Q (signal_4023) ) ;
    buf_clk cell_2837 ( .C (clk), .D (signal_4030), .Q (signal_4031) ) ;
    buf_clk cell_2845 ( .C (clk), .D (signal_4038), .Q (signal_4039) ) ;
    buf_clk cell_2853 ( .C (clk), .D (signal_4046), .Q (signal_4047) ) ;
    buf_clk cell_2861 ( .C (clk), .D (signal_4054), .Q (signal_4055) ) ;
    buf_clk cell_2869 ( .C (clk), .D (signal_4062), .Q (signal_4063) ) ;
    buf_clk cell_2877 ( .C (clk), .D (signal_4070), .Q (signal_4071) ) ;
    buf_clk cell_2885 ( .C (clk), .D (signal_4078), .Q (signal_4079) ) ;
    buf_clk cell_2893 ( .C (clk), .D (signal_4086), .Q (signal_4087) ) ;
    buf_clk cell_2901 ( .C (clk), .D (signal_4094), .Q (signal_4095) ) ;
    buf_clk cell_2909 ( .C (clk), .D (signal_4102), .Q (signal_4103) ) ;
    buf_clk cell_2917 ( .C (clk), .D (signal_4110), .Q (signal_4111) ) ;
    buf_clk cell_2925 ( .C (clk), .D (signal_4118), .Q (signal_4119) ) ;
    buf_clk cell_2933 ( .C (clk), .D (signal_4126), .Q (signal_4127) ) ;
    buf_clk cell_2941 ( .C (clk), .D (signal_4134), .Q (signal_4135) ) ;
    buf_clk cell_2949 ( .C (clk), .D (signal_4142), .Q (signal_4143) ) ;
    buf_clk cell_2957 ( .C (clk), .D (signal_4150), .Q (signal_4151) ) ;
    buf_clk cell_2965 ( .C (clk), .D (signal_4158), .Q (signal_4159) ) ;
    buf_clk cell_2973 ( .C (clk), .D (signal_4166), .Q (signal_4167) ) ;
    buf_clk cell_2981 ( .C (clk), .D (signal_4174), .Q (signal_4175) ) ;
    buf_clk cell_2989 ( .C (clk), .D (signal_4182), .Q (signal_4183) ) ;
    buf_clk cell_2997 ( .C (clk), .D (signal_4190), .Q (signal_4191) ) ;
    buf_clk cell_3005 ( .C (clk), .D (signal_4198), .Q (signal_4199) ) ;
    buf_clk cell_3013 ( .C (clk), .D (signal_4206), .Q (signal_4207) ) ;
    buf_clk cell_3021 ( .C (clk), .D (signal_4214), .Q (signal_4215) ) ;
    buf_clk cell_3029 ( .C (clk), .D (signal_4222), .Q (signal_4223) ) ;
    buf_clk cell_3037 ( .C (clk), .D (signal_4230), .Q (signal_4231) ) ;
    buf_clk cell_3045 ( .C (clk), .D (signal_4238), .Q (signal_4239) ) ;
    buf_clk cell_3053 ( .C (clk), .D (signal_4246), .Q (signal_4247) ) ;
    buf_clk cell_3061 ( .C (clk), .D (signal_4254), .Q (signal_4255) ) ;
    buf_clk cell_3069 ( .C (clk), .D (signal_4262), .Q (signal_4263) ) ;
    buf_clk cell_3077 ( .C (clk), .D (signal_4270), .Q (signal_4271) ) ;
    buf_clk cell_3085 ( .C (clk), .D (signal_4278), .Q (signal_4279) ) ;
    buf_clk cell_3093 ( .C (clk), .D (signal_4286), .Q (signal_4287) ) ;
    buf_clk cell_3101 ( .C (clk), .D (signal_4294), .Q (signal_4295) ) ;
    buf_clk cell_3109 ( .C (clk), .D (signal_4302), .Q (signal_4303) ) ;
    buf_clk cell_3117 ( .C (clk), .D (signal_4310), .Q (signal_4311) ) ;
    buf_clk cell_3125 ( .C (clk), .D (signal_4318), .Q (signal_4319) ) ;
    buf_clk cell_3133 ( .C (clk), .D (signal_4326), .Q (signal_4327) ) ;
    buf_clk cell_3141 ( .C (clk), .D (signal_4334), .Q (signal_4335) ) ;
    buf_clk cell_3149 ( .C (clk), .D (signal_4342), .Q (signal_4343) ) ;
    buf_clk cell_3157 ( .C (clk), .D (signal_4350), .Q (signal_4351) ) ;
    buf_clk cell_3165 ( .C (clk), .D (signal_4358), .Q (signal_4359) ) ;
    buf_clk cell_3169 ( .C (clk), .D (signal_4362), .Q (signal_4363) ) ;
    buf_clk cell_3171 ( .C (clk), .D (signal_4364), .Q (signal_4365) ) ;
    buf_clk cell_3173 ( .C (clk), .D (signal_4366), .Q (signal_4367) ) ;
    buf_clk cell_3175 ( .C (clk), .D (signal_4368), .Q (signal_4369) ) ;
    buf_clk cell_3177 ( .C (clk), .D (signal_4370), .Q (signal_4371) ) ;
    buf_clk cell_3179 ( .C (clk), .D (signal_4372), .Q (signal_4373) ) ;
    buf_clk cell_3181 ( .C (clk), .D (signal_4374), .Q (signal_4375) ) ;
    buf_clk cell_3183 ( .C (clk), .D (signal_4376), .Q (signal_4377) ) ;
    buf_clk cell_3185 ( .C (clk), .D (signal_4378), .Q (signal_4379) ) ;
    buf_clk cell_3187 ( .C (clk), .D (signal_4380), .Q (signal_4381) ) ;
    buf_clk cell_3189 ( .C (clk), .D (signal_4382), .Q (signal_4383) ) ;
    buf_clk cell_3191 ( .C (clk), .D (signal_4384), .Q (signal_4385) ) ;
    buf_clk cell_3193 ( .C (clk), .D (signal_4386), .Q (signal_4387) ) ;
    buf_clk cell_3195 ( .C (clk), .D (signal_4388), .Q (signal_4389) ) ;
    buf_clk cell_3197 ( .C (clk), .D (signal_4390), .Q (signal_4391) ) ;
    buf_clk cell_3199 ( .C (clk), .D (signal_4392), .Q (signal_4393) ) ;
    buf_clk cell_3201 ( .C (clk), .D (signal_4394), .Q (signal_4395) ) ;
    buf_clk cell_3203 ( .C (clk), .D (signal_4396), .Q (signal_4397) ) ;
    buf_clk cell_3205 ( .C (clk), .D (signal_4398), .Q (signal_4399) ) ;
    buf_clk cell_3207 ( .C (clk), .D (signal_4400), .Q (signal_4401) ) ;
    buf_clk cell_3209 ( .C (clk), .D (signal_4402), .Q (signal_4403) ) ;
    buf_clk cell_3211 ( .C (clk), .D (signal_4404), .Q (signal_4405) ) ;
    buf_clk cell_3213 ( .C (clk), .D (signal_4406), .Q (signal_4407) ) ;
    buf_clk cell_3215 ( .C (clk), .D (signal_4408), .Q (signal_4409) ) ;
    buf_clk cell_3217 ( .C (clk), .D (signal_4410), .Q (signal_4411) ) ;
    buf_clk cell_3219 ( .C (clk), .D (signal_4412), .Q (signal_4413) ) ;
    buf_clk cell_3221 ( .C (clk), .D (signal_4414), .Q (signal_4415) ) ;
    buf_clk cell_3223 ( .C (clk), .D (signal_4416), .Q (signal_4417) ) ;
    buf_clk cell_3225 ( .C (clk), .D (signal_4418), .Q (signal_4419) ) ;
    buf_clk cell_3227 ( .C (clk), .D (signal_4420), .Q (signal_4421) ) ;
    buf_clk cell_3229 ( .C (clk), .D (signal_4422), .Q (signal_4423) ) ;
    buf_clk cell_3231 ( .C (clk), .D (signal_4424), .Q (signal_4425) ) ;
    buf_clk cell_3233 ( .C (clk), .D (signal_4426), .Q (signal_4427) ) ;
    buf_clk cell_3235 ( .C (clk), .D (signal_4428), .Q (signal_4429) ) ;
    buf_clk cell_3237 ( .C (clk), .D (signal_4430), .Q (signal_4431) ) ;
    buf_clk cell_3239 ( .C (clk), .D (signal_4432), .Q (signal_4433) ) ;
    buf_clk cell_3241 ( .C (clk), .D (signal_4434), .Q (signal_4435) ) ;
    buf_clk cell_3243 ( .C (clk), .D (signal_4436), .Q (signal_4437) ) ;
    buf_clk cell_3245 ( .C (clk), .D (signal_4438), .Q (signal_4439) ) ;
    buf_clk cell_3247 ( .C (clk), .D (signal_4440), .Q (signal_4441) ) ;
    buf_clk cell_3249 ( .C (clk), .D (signal_4442), .Q (signal_4443) ) ;
    buf_clk cell_3251 ( .C (clk), .D (signal_4444), .Q (signal_4445) ) ;
    buf_clk cell_3253 ( .C (clk), .D (signal_4446), .Q (signal_4447) ) ;
    buf_clk cell_3255 ( .C (clk), .D (signal_4448), .Q (signal_4449) ) ;
    buf_clk cell_3257 ( .C (clk), .D (signal_4450), .Q (signal_4451) ) ;
    buf_clk cell_3259 ( .C (clk), .D (signal_4452), .Q (signal_4453) ) ;
    buf_clk cell_3261 ( .C (clk), .D (signal_4454), .Q (signal_4455) ) ;
    buf_clk cell_3263 ( .C (clk), .D (signal_4456), .Q (signal_4457) ) ;
    buf_clk cell_3265 ( .C (clk), .D (signal_4458), .Q (signal_4459) ) ;
    buf_clk cell_3267 ( .C (clk), .D (signal_4460), .Q (signal_4461) ) ;
    buf_clk cell_3269 ( .C (clk), .D (signal_4462), .Q (signal_4463) ) ;
    buf_clk cell_3271 ( .C (clk), .D (signal_4464), .Q (signal_4465) ) ;
    buf_clk cell_3273 ( .C (clk), .D (signal_4466), .Q (signal_4467) ) ;
    buf_clk cell_3275 ( .C (clk), .D (signal_4468), .Q (signal_4469) ) ;
    buf_clk cell_3277 ( .C (clk), .D (signal_4470), .Q (signal_4471) ) ;
    buf_clk cell_3279 ( .C (clk), .D (signal_4472), .Q (signal_4473) ) ;
    buf_clk cell_3281 ( .C (clk), .D (signal_4474), .Q (signal_4475) ) ;
    buf_clk cell_3283 ( .C (clk), .D (signal_4476), .Q (signal_4477) ) ;
    buf_clk cell_3285 ( .C (clk), .D (signal_4478), .Q (signal_4479) ) ;
    buf_clk cell_3287 ( .C (clk), .D (signal_4480), .Q (signal_4481) ) ;
    buf_clk cell_3289 ( .C (clk), .D (signal_4482), .Q (signal_4483) ) ;
    buf_clk cell_3291 ( .C (clk), .D (signal_4484), .Q (signal_4485) ) ;
    buf_clk cell_3293 ( .C (clk), .D (signal_4486), .Q (signal_4487) ) ;
    buf_clk cell_3295 ( .C (clk), .D (signal_4488), .Q (signal_4489) ) ;
    buf_clk cell_3297 ( .C (clk), .D (signal_4490), .Q (signal_4491) ) ;
    buf_clk cell_3299 ( .C (clk), .D (signal_4492), .Q (signal_4493) ) ;
    buf_clk cell_3301 ( .C (clk), .D (signal_4494), .Q (signal_4495) ) ;
    buf_clk cell_3303 ( .C (clk), .D (signal_4496), .Q (signal_4497) ) ;
    buf_clk cell_3305 ( .C (clk), .D (signal_4498), .Q (signal_4499) ) ;
    buf_clk cell_3307 ( .C (clk), .D (signal_4500), .Q (signal_4501) ) ;
    buf_clk cell_3309 ( .C (clk), .D (signal_4502), .Q (signal_4503) ) ;
    buf_clk cell_3311 ( .C (clk), .D (signal_4504), .Q (signal_4505) ) ;
    buf_clk cell_3313 ( .C (clk), .D (signal_4506), .Q (signal_4507) ) ;
    buf_clk cell_3315 ( .C (clk), .D (signal_4508), .Q (signal_4509) ) ;
    buf_clk cell_3317 ( .C (clk), .D (signal_4510), .Q (signal_4511) ) ;
    buf_clk cell_3319 ( .C (clk), .D (signal_4512), .Q (signal_4513) ) ;
    buf_clk cell_3321 ( .C (clk), .D (signal_4514), .Q (signal_4515) ) ;
    buf_clk cell_3323 ( .C (clk), .D (signal_4516), .Q (signal_4517) ) ;
    buf_clk cell_3325 ( .C (clk), .D (signal_4518), .Q (signal_4519) ) ;
    buf_clk cell_3327 ( .C (clk), .D (signal_4520), .Q (signal_4521) ) ;
    buf_clk cell_3329 ( .C (clk), .D (signal_4522), .Q (signal_4523) ) ;
    buf_clk cell_3331 ( .C (clk), .D (signal_4524), .Q (signal_4525) ) ;
    buf_clk cell_3333 ( .C (clk), .D (signal_4526), .Q (signal_4527) ) ;
    buf_clk cell_3335 ( .C (clk), .D (signal_4528), .Q (signal_4529) ) ;
    buf_clk cell_3337 ( .C (clk), .D (signal_4530), .Q (signal_4531) ) ;
    buf_clk cell_3339 ( .C (clk), .D (signal_4532), .Q (signal_4533) ) ;
    buf_clk cell_3341 ( .C (clk), .D (signal_4534), .Q (signal_4535) ) ;
    buf_clk cell_3343 ( .C (clk), .D (signal_4536), .Q (signal_4537) ) ;
    buf_clk cell_3345 ( .C (clk), .D (signal_4538), .Q (signal_4539) ) ;
    buf_clk cell_3347 ( .C (clk), .D (signal_4540), .Q (signal_4541) ) ;
    buf_clk cell_3349 ( .C (clk), .D (signal_4542), .Q (signal_4543) ) ;
    buf_clk cell_3351 ( .C (clk), .D (signal_4544), .Q (signal_4545) ) ;
    buf_clk cell_3353 ( .C (clk), .D (signal_4546), .Q (signal_4547) ) ;
    buf_clk cell_3355 ( .C (clk), .D (signal_4548), .Q (signal_4549) ) ;
    buf_clk cell_3357 ( .C (clk), .D (signal_4550), .Q (signal_4551) ) ;
    buf_clk cell_3359 ( .C (clk), .D (signal_4552), .Q (signal_4553) ) ;
    buf_clk cell_3493 ( .C (clk), .D (signal_4686), .Q (signal_4687) ) ;
    buf_clk cell_3501 ( .C (clk), .D (signal_4694), .Q (signal_4695) ) ;
    buf_clk cell_3509 ( .C (clk), .D (signal_4702), .Q (signal_4703) ) ;
    buf_clk cell_3517 ( .C (clk), .D (signal_4710), .Q (signal_4711) ) ;
    buf_clk cell_3525 ( .C (clk), .D (signal_4718), .Q (signal_4719) ) ;
    buf_clk cell_3533 ( .C (clk), .D (signal_4726), .Q (signal_4727) ) ;
    buf_clk cell_3541 ( .C (clk), .D (signal_4734), .Q (signal_4735) ) ;
    buf_clk cell_3549 ( .C (clk), .D (signal_4742), .Q (signal_4743) ) ;
    buf_clk cell_3557 ( .C (clk), .D (signal_4750), .Q (signal_4751) ) ;
    buf_clk cell_3565 ( .C (clk), .D (signal_4758), .Q (signal_4759) ) ;

    /* cells in depth 7 */
    buf_clk cell_2142 ( .C (clk), .D (signal_2375), .Q (signal_3336) ) ;
    buf_clk cell_2150 ( .C (clk), .D (signal_3343), .Q (signal_3344) ) ;
    buf_clk cell_2158 ( .C (clk), .D (signal_3351), .Q (signal_3352) ) ;
    buf_clk cell_2166 ( .C (clk), .D (signal_3359), .Q (signal_3360) ) ;
    buf_clk cell_2174 ( .C (clk), .D (signal_3367), .Q (signal_3368) ) ;
    buf_clk cell_2182 ( .C (clk), .D (signal_3375), .Q (signal_3376) ) ;
    buf_clk cell_2190 ( .C (clk), .D (signal_3383), .Q (signal_3384) ) ;
    buf_clk cell_2198 ( .C (clk), .D (signal_3391), .Q (signal_3392) ) ;
    buf_clk cell_2206 ( .C (clk), .D (signal_3399), .Q (signal_3400) ) ;
    buf_clk cell_2214 ( .C (clk), .D (signal_3407), .Q (signal_3408) ) ;
    buf_clk cell_2222 ( .C (clk), .D (signal_3415), .Q (signal_3416) ) ;
    buf_clk cell_2230 ( .C (clk), .D (signal_3423), .Q (signal_3424) ) ;
    buf_clk cell_2238 ( .C (clk), .D (signal_3431), .Q (signal_3432) ) ;
    buf_clk cell_2246 ( .C (clk), .D (signal_3439), .Q (signal_3440) ) ;
    buf_clk cell_2254 ( .C (clk), .D (signal_3447), .Q (signal_3448) ) ;
    buf_clk cell_2262 ( .C (clk), .D (signal_3455), .Q (signal_3456) ) ;
    buf_clk cell_2270 ( .C (clk), .D (signal_3463), .Q (signal_3464) ) ;
    buf_clk cell_2278 ( .C (clk), .D (signal_3471), .Q (signal_3472) ) ;
    buf_clk cell_2286 ( .C (clk), .D (signal_3479), .Q (signal_3480) ) ;
    buf_clk cell_2294 ( .C (clk), .D (signal_3487), .Q (signal_3488) ) ;
    buf_clk cell_2302 ( .C (clk), .D (signal_3495), .Q (signal_3496) ) ;
    buf_clk cell_2310 ( .C (clk), .D (signal_3503), .Q (signal_3504) ) ;
    buf_clk cell_2318 ( .C (clk), .D (signal_3511), .Q (signal_3512) ) ;
    buf_clk cell_2326 ( .C (clk), .D (signal_3519), .Q (signal_3520) ) ;
    buf_clk cell_2334 ( .C (clk), .D (signal_3527), .Q (signal_3528) ) ;
    buf_clk cell_2342 ( .C (clk), .D (signal_3535), .Q (signal_3536) ) ;
    buf_clk cell_2350 ( .C (clk), .D (signal_3543), .Q (signal_3544) ) ;
    buf_clk cell_2358 ( .C (clk), .D (signal_3551), .Q (signal_3552) ) ;
    buf_clk cell_2366 ( .C (clk), .D (signal_3559), .Q (signal_3560) ) ;
    buf_clk cell_2374 ( .C (clk), .D (signal_3567), .Q (signal_3568) ) ;
    buf_clk cell_2382 ( .C (clk), .D (signal_3575), .Q (signal_3576) ) ;
    buf_clk cell_2390 ( .C (clk), .D (signal_3583), .Q (signal_3584) ) ;
    buf_clk cell_2398 ( .C (clk), .D (signal_3591), .Q (signal_3592) ) ;
    buf_clk cell_2406 ( .C (clk), .D (signal_3599), .Q (signal_3600) ) ;
    buf_clk cell_2414 ( .C (clk), .D (signal_3607), .Q (signal_3608) ) ;
    buf_clk cell_2422 ( .C (clk), .D (signal_3615), .Q (signal_3616) ) ;
    buf_clk cell_2430 ( .C (clk), .D (signal_3623), .Q (signal_3624) ) ;
    buf_clk cell_2438 ( .C (clk), .D (signal_3631), .Q (signal_3632) ) ;
    buf_clk cell_2446 ( .C (clk), .D (signal_3639), .Q (signal_3640) ) ;
    buf_clk cell_2454 ( .C (clk), .D (signal_3647), .Q (signal_3648) ) ;
    buf_clk cell_2462 ( .C (clk), .D (signal_3655), .Q (signal_3656) ) ;
    buf_clk cell_2470 ( .C (clk), .D (signal_3663), .Q (signal_3664) ) ;
    buf_clk cell_2478 ( .C (clk), .D (signal_3671), .Q (signal_3672) ) ;
    buf_clk cell_2486 ( .C (clk), .D (signal_3679), .Q (signal_3680) ) ;
    buf_clk cell_2494 ( .C (clk), .D (signal_3687), .Q (signal_3688) ) ;
    buf_clk cell_2502 ( .C (clk), .D (signal_3695), .Q (signal_3696) ) ;
    buf_clk cell_2510 ( .C (clk), .D (signal_3703), .Q (signal_3704) ) ;
    buf_clk cell_2518 ( .C (clk), .D (signal_3711), .Q (signal_3712) ) ;
    buf_clk cell_2526 ( .C (clk), .D (signal_3719), .Q (signal_3720) ) ;
    buf_clk cell_2534 ( .C (clk), .D (signal_3727), .Q (signal_3728) ) ;
    buf_clk cell_2542 ( .C (clk), .D (signal_3735), .Q (signal_3736) ) ;
    buf_clk cell_2550 ( .C (clk), .D (signal_3743), .Q (signal_3744) ) ;
    buf_clk cell_2558 ( .C (clk), .D (signal_3751), .Q (signal_3752) ) ;
    buf_clk cell_2566 ( .C (clk), .D (signal_3759), .Q (signal_3760) ) ;
    buf_clk cell_2574 ( .C (clk), .D (signal_3767), .Q (signal_3768) ) ;
    buf_clk cell_2582 ( .C (clk), .D (signal_3775), .Q (signal_3776) ) ;
    buf_clk cell_2590 ( .C (clk), .D (signal_3783), .Q (signal_3784) ) ;
    buf_clk cell_2598 ( .C (clk), .D (signal_3791), .Q (signal_3792) ) ;
    buf_clk cell_2606 ( .C (clk), .D (signal_3799), .Q (signal_3800) ) ;
    buf_clk cell_2614 ( .C (clk), .D (signal_3807), .Q (signal_3808) ) ;
    buf_clk cell_2622 ( .C (clk), .D (signal_3815), .Q (signal_3816) ) ;
    buf_clk cell_2630 ( .C (clk), .D (signal_3823), .Q (signal_3824) ) ;
    buf_clk cell_2638 ( .C (clk), .D (signal_3831), .Q (signal_3832) ) ;
    buf_clk cell_2646 ( .C (clk), .D (signal_3839), .Q (signal_3840) ) ;
    buf_clk cell_2654 ( .C (clk), .D (signal_3847), .Q (signal_3848) ) ;
    buf_clk cell_2662 ( .C (clk), .D (signal_3855), .Q (signal_3856) ) ;
    buf_clk cell_2670 ( .C (clk), .D (signal_3863), .Q (signal_3864) ) ;
    buf_clk cell_2678 ( .C (clk), .D (signal_3871), .Q (signal_3872) ) ;
    buf_clk cell_2686 ( .C (clk), .D (signal_3879), .Q (signal_3880) ) ;
    buf_clk cell_2694 ( .C (clk), .D (signal_3887), .Q (signal_3888) ) ;
    buf_clk cell_2702 ( .C (clk), .D (signal_3895), .Q (signal_3896) ) ;
    buf_clk cell_2710 ( .C (clk), .D (signal_3903), .Q (signal_3904) ) ;
    buf_clk cell_2718 ( .C (clk), .D (signal_3911), .Q (signal_3912) ) ;
    buf_clk cell_2726 ( .C (clk), .D (signal_3919), .Q (signal_3920) ) ;
    buf_clk cell_2734 ( .C (clk), .D (signal_3927), .Q (signal_3928) ) ;
    buf_clk cell_2742 ( .C (clk), .D (signal_3935), .Q (signal_3936) ) ;
    buf_clk cell_2750 ( .C (clk), .D (signal_3943), .Q (signal_3944) ) ;
    buf_clk cell_2758 ( .C (clk), .D (signal_3951), .Q (signal_3952) ) ;
    buf_clk cell_2766 ( .C (clk), .D (signal_3959), .Q (signal_3960) ) ;
    buf_clk cell_2774 ( .C (clk), .D (signal_3967), .Q (signal_3968) ) ;
    buf_clk cell_2782 ( .C (clk), .D (signal_3975), .Q (signal_3976) ) ;
    buf_clk cell_2790 ( .C (clk), .D (signal_3983), .Q (signal_3984) ) ;
    buf_clk cell_2798 ( .C (clk), .D (signal_3991), .Q (signal_3992) ) ;
    buf_clk cell_2806 ( .C (clk), .D (signal_3999), .Q (signal_4000) ) ;
    buf_clk cell_2814 ( .C (clk), .D (signal_4007), .Q (signal_4008) ) ;
    buf_clk cell_2822 ( .C (clk), .D (signal_4015), .Q (signal_4016) ) ;
    buf_clk cell_2830 ( .C (clk), .D (signal_4023), .Q (signal_4024) ) ;
    buf_clk cell_2838 ( .C (clk), .D (signal_4031), .Q (signal_4032) ) ;
    buf_clk cell_2846 ( .C (clk), .D (signal_4039), .Q (signal_4040) ) ;
    buf_clk cell_2854 ( .C (clk), .D (signal_4047), .Q (signal_4048) ) ;
    buf_clk cell_2862 ( .C (clk), .D (signal_4055), .Q (signal_4056) ) ;
    buf_clk cell_2870 ( .C (clk), .D (signal_4063), .Q (signal_4064) ) ;
    buf_clk cell_2878 ( .C (clk), .D (signal_4071), .Q (signal_4072) ) ;
    buf_clk cell_2886 ( .C (clk), .D (signal_4079), .Q (signal_4080) ) ;
    buf_clk cell_2894 ( .C (clk), .D (signal_4087), .Q (signal_4088) ) ;
    buf_clk cell_2902 ( .C (clk), .D (signal_4095), .Q (signal_4096) ) ;
    buf_clk cell_2910 ( .C (clk), .D (signal_4103), .Q (signal_4104) ) ;
    buf_clk cell_2918 ( .C (clk), .D (signal_4111), .Q (signal_4112) ) ;
    buf_clk cell_2926 ( .C (clk), .D (signal_4119), .Q (signal_4120) ) ;
    buf_clk cell_2934 ( .C (clk), .D (signal_4127), .Q (signal_4128) ) ;
    buf_clk cell_2942 ( .C (clk), .D (signal_4135), .Q (signal_4136) ) ;
    buf_clk cell_2950 ( .C (clk), .D (signal_4143), .Q (signal_4144) ) ;
    buf_clk cell_2958 ( .C (clk), .D (signal_4151), .Q (signal_4152) ) ;
    buf_clk cell_2966 ( .C (clk), .D (signal_4159), .Q (signal_4160) ) ;
    buf_clk cell_2974 ( .C (clk), .D (signal_4167), .Q (signal_4168) ) ;
    buf_clk cell_2982 ( .C (clk), .D (signal_4175), .Q (signal_4176) ) ;
    buf_clk cell_2990 ( .C (clk), .D (signal_4183), .Q (signal_4184) ) ;
    buf_clk cell_2998 ( .C (clk), .D (signal_4191), .Q (signal_4192) ) ;
    buf_clk cell_3006 ( .C (clk), .D (signal_4199), .Q (signal_4200) ) ;
    buf_clk cell_3014 ( .C (clk), .D (signal_4207), .Q (signal_4208) ) ;
    buf_clk cell_3022 ( .C (clk), .D (signal_4215), .Q (signal_4216) ) ;
    buf_clk cell_3030 ( .C (clk), .D (signal_4223), .Q (signal_4224) ) ;
    buf_clk cell_3038 ( .C (clk), .D (signal_4231), .Q (signal_4232) ) ;
    buf_clk cell_3046 ( .C (clk), .D (signal_4239), .Q (signal_4240) ) ;
    buf_clk cell_3054 ( .C (clk), .D (signal_4247), .Q (signal_4248) ) ;
    buf_clk cell_3062 ( .C (clk), .D (signal_4255), .Q (signal_4256) ) ;
    buf_clk cell_3070 ( .C (clk), .D (signal_4263), .Q (signal_4264) ) ;
    buf_clk cell_3078 ( .C (clk), .D (signal_4271), .Q (signal_4272) ) ;
    buf_clk cell_3086 ( .C (clk), .D (signal_4279), .Q (signal_4280) ) ;
    buf_clk cell_3094 ( .C (clk), .D (signal_4287), .Q (signal_4288) ) ;
    buf_clk cell_3102 ( .C (clk), .D (signal_4295), .Q (signal_4296) ) ;
    buf_clk cell_3110 ( .C (clk), .D (signal_4303), .Q (signal_4304) ) ;
    buf_clk cell_3118 ( .C (clk), .D (signal_4311), .Q (signal_4312) ) ;
    buf_clk cell_3126 ( .C (clk), .D (signal_4319), .Q (signal_4320) ) ;
    buf_clk cell_3134 ( .C (clk), .D (signal_4327), .Q (signal_4328) ) ;
    buf_clk cell_3142 ( .C (clk), .D (signal_4335), .Q (signal_4336) ) ;
    buf_clk cell_3150 ( .C (clk), .D (signal_4343), .Q (signal_4344) ) ;
    buf_clk cell_3158 ( .C (clk), .D (signal_4351), .Q (signal_4352) ) ;
    buf_clk cell_3166 ( .C (clk), .D (signal_4359), .Q (signal_4360) ) ;
    buf_clk cell_3360 ( .C (clk), .D (signal_935), .Q (signal_4554) ) ;
    buf_clk cell_3362 ( .C (clk), .D (signal_1980), .Q (signal_4556) ) ;
    buf_clk cell_3364 ( .C (clk), .D (signal_937), .Q (signal_4558) ) ;
    buf_clk cell_3366 ( .C (clk), .D (signal_1978), .Q (signal_4560) ) ;
    buf_clk cell_3368 ( .C (clk), .D (signal_939), .Q (signal_4562) ) ;
    buf_clk cell_3370 ( .C (clk), .D (signal_1976), .Q (signal_4564) ) ;
    buf_clk cell_3372 ( .C (clk), .D (signal_941), .Q (signal_4566) ) ;
    buf_clk cell_3374 ( .C (clk), .D (signal_1974), .Q (signal_4568) ) ;
    buf_clk cell_3376 ( .C (clk), .D (signal_943), .Q (signal_4570) ) ;
    buf_clk cell_3378 ( .C (clk), .D (signal_1972), .Q (signal_4572) ) ;
    buf_clk cell_3380 ( .C (clk), .D (signal_945), .Q (signal_4574) ) ;
    buf_clk cell_3382 ( .C (clk), .D (signal_1970), .Q (signal_4576) ) ;
    buf_clk cell_3384 ( .C (clk), .D (signal_947), .Q (signal_4578) ) ;
    buf_clk cell_3386 ( .C (clk), .D (signal_1968), .Q (signal_4580) ) ;
    buf_clk cell_3388 ( .C (clk), .D (signal_949), .Q (signal_4582) ) ;
    buf_clk cell_3390 ( .C (clk), .D (signal_1966), .Q (signal_4584) ) ;
    buf_clk cell_3392 ( .C (clk), .D (signal_951), .Q (signal_4586) ) ;
    buf_clk cell_3394 ( .C (clk), .D (signal_1988), .Q (signal_4588) ) ;
    buf_clk cell_3396 ( .C (clk), .D (signal_953), .Q (signal_4590) ) ;
    buf_clk cell_3398 ( .C (clk), .D (signal_1986), .Q (signal_4592) ) ;
    buf_clk cell_3400 ( .C (clk), .D (signal_955), .Q (signal_4594) ) ;
    buf_clk cell_3402 ( .C (clk), .D (signal_1984), .Q (signal_4596) ) ;
    buf_clk cell_3404 ( .C (clk), .D (signal_957), .Q (signal_4598) ) ;
    buf_clk cell_3406 ( .C (clk), .D (signal_1982), .Q (signal_4600) ) ;
    buf_clk cell_3408 ( .C (clk), .D (signal_959), .Q (signal_4602) ) ;
    buf_clk cell_3410 ( .C (clk), .D (signal_1996), .Q (signal_4604) ) ;
    buf_clk cell_3412 ( .C (clk), .D (signal_961), .Q (signal_4606) ) ;
    buf_clk cell_3414 ( .C (clk), .D (signal_1994), .Q (signal_4608) ) ;
    buf_clk cell_3416 ( .C (clk), .D (signal_963), .Q (signal_4610) ) ;
    buf_clk cell_3418 ( .C (clk), .D (signal_1992), .Q (signal_4612) ) ;
    buf_clk cell_3420 ( .C (clk), .D (signal_965), .Q (signal_4614) ) ;
    buf_clk cell_3422 ( .C (clk), .D (signal_1990), .Q (signal_4616) ) ;
    buf_clk cell_3424 ( .C (clk), .D (signal_967), .Q (signal_4618) ) ;
    buf_clk cell_3426 ( .C (clk), .D (signal_1916), .Q (signal_4620) ) ;
    buf_clk cell_3428 ( .C (clk), .D (signal_969), .Q (signal_4622) ) ;
    buf_clk cell_3430 ( .C (clk), .D (signal_1914), .Q (signal_4624) ) ;
    buf_clk cell_3432 ( .C (clk), .D (signal_971), .Q (signal_4626) ) ;
    buf_clk cell_3434 ( .C (clk), .D (signal_1912), .Q (signal_4628) ) ;
    buf_clk cell_3436 ( .C (clk), .D (signal_973), .Q (signal_4630) ) ;
    buf_clk cell_3438 ( .C (clk), .D (signal_1910), .Q (signal_4632) ) ;
    buf_clk cell_3440 ( .C (clk), .D (signal_975), .Q (signal_4634) ) ;
    buf_clk cell_3442 ( .C (clk), .D (signal_1908), .Q (signal_4636) ) ;
    buf_clk cell_3444 ( .C (clk), .D (signal_977), .Q (signal_4638) ) ;
    buf_clk cell_3446 ( .C (clk), .D (signal_1906), .Q (signal_4640) ) ;
    buf_clk cell_3448 ( .C (clk), .D (signal_979), .Q (signal_4642) ) ;
    buf_clk cell_3450 ( .C (clk), .D (signal_1904), .Q (signal_4644) ) ;
    buf_clk cell_3452 ( .C (clk), .D (signal_981), .Q (signal_4646) ) ;
    buf_clk cell_3454 ( .C (clk), .D (signal_1902), .Q (signal_4648) ) ;
    buf_clk cell_3456 ( .C (clk), .D (signal_983), .Q (signal_4650) ) ;
    buf_clk cell_3458 ( .C (clk), .D (signal_1900), .Q (signal_4652) ) ;
    buf_clk cell_3460 ( .C (clk), .D (signal_985), .Q (signal_4654) ) ;
    buf_clk cell_3462 ( .C (clk), .D (signal_1898), .Q (signal_4656) ) ;
    buf_clk cell_3464 ( .C (clk), .D (signal_987), .Q (signal_4658) ) ;
    buf_clk cell_3466 ( .C (clk), .D (signal_1896), .Q (signal_4660) ) ;
    buf_clk cell_3468 ( .C (clk), .D (signal_989), .Q (signal_4662) ) ;
    buf_clk cell_3470 ( .C (clk), .D (signal_1894), .Q (signal_4664) ) ;
    buf_clk cell_3472 ( .C (clk), .D (signal_991), .Q (signal_4666) ) ;
    buf_clk cell_3474 ( .C (clk), .D (signal_1892), .Q (signal_4668) ) ;
    buf_clk cell_3476 ( .C (clk), .D (signal_993), .Q (signal_4670) ) ;
    buf_clk cell_3478 ( .C (clk), .D (signal_1890), .Q (signal_4672) ) ;
    buf_clk cell_3480 ( .C (clk), .D (signal_995), .Q (signal_4674) ) ;
    buf_clk cell_3482 ( .C (clk), .D (signal_1888), .Q (signal_4676) ) ;
    buf_clk cell_3484 ( .C (clk), .D (signal_997), .Q (signal_4678) ) ;
    buf_clk cell_3486 ( .C (clk), .D (signal_1886), .Q (signal_4680) ) ;
    buf_clk cell_3494 ( .C (clk), .D (signal_4687), .Q (signal_4688) ) ;
    buf_clk cell_3502 ( .C (clk), .D (signal_4695), .Q (signal_4696) ) ;
    buf_clk cell_3510 ( .C (clk), .D (signal_4703), .Q (signal_4704) ) ;
    buf_clk cell_3518 ( .C (clk), .D (signal_4711), .Q (signal_4712) ) ;
    buf_clk cell_3526 ( .C (clk), .D (signal_4719), .Q (signal_4720) ) ;
    buf_clk cell_3534 ( .C (clk), .D (signal_4727), .Q (signal_4728) ) ;
    buf_clk cell_3542 ( .C (clk), .D (signal_4735), .Q (signal_4736) ) ;
    buf_clk cell_3550 ( .C (clk), .D (signal_4743), .Q (signal_4744) ) ;
    buf_clk cell_3558 ( .C (clk), .D (signal_4751), .Q (signal_4752) ) ;
    buf_clk cell_3566 ( .C (clk), .D (signal_4759), .Q (signal_4760) ) ;

    /* cells in depth 8 */
    mux2_masked #(.security_order(1), .pipeline(1)) cell_0 ( .s (signal_3337), .b ({signal_1708, signal_774}), .a ({signal_3353, signal_3345}), .c ({signal_1734, signal_870}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_2 ( .s (signal_3337), .b ({signal_1707, signal_772}), .a ({signal_3369, signal_3361}), .c ({signal_1736, signal_868}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_4 ( .s (signal_3337), .b ({signal_1717, signal_770}), .a ({signal_3385, signal_3377}), .c ({signal_1738, signal_866}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_6 ( .s (signal_3337), .b ({signal_1711, signal_768}), .a ({signal_3401, signal_3393}), .c ({signal_1740, signal_864}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_8 ( .s (signal_3337), .b ({signal_1719, signal_766}), .a ({signal_3417, signal_3409}), .c ({signal_1742, signal_862}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_10 ( .s (signal_3337), .b ({signal_1712, signal_764}), .a ({signal_3433, signal_3425}), .c ({signal_1744, signal_860}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_12 ( .s (signal_3337), .b ({signal_1718, signal_762}), .a ({signal_3449, signal_3441}), .c ({signal_1746, signal_858}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_14 ( .s (signal_3337), .b ({signal_1709, signal_760}), .a ({signal_3465, signal_3457}), .c ({signal_1748, signal_856}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_16 ( .s (signal_3337), .b ({signal_1706, signal_758}), .a ({signal_3481, signal_3473}), .c ({signal_1750, signal_854}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_18 ( .s (signal_3337), .b ({signal_1701, signal_756}), .a ({signal_3497, signal_3489}), .c ({signal_1752, signal_852}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_20 ( .s (signal_3337), .b ({signal_1702, signal_754}), .a ({signal_3513, signal_3505}), .c ({signal_1754, signal_850}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_22 ( .s (signal_3337), .b ({signal_1716, signal_752}), .a ({signal_3529, signal_3521}), .c ({signal_1756, signal_848}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_24 ( .s (signal_3337), .b ({signal_1710, signal_750}), .a ({signal_3545, signal_3537}), .c ({signal_1758, signal_846}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_26 ( .s (signal_3337), .b ({signal_1704, signal_748}), .a ({signal_3561, signal_3553}), .c ({signal_1760, signal_844}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_28 ( .s (signal_3337), .b ({signal_1703, signal_746}), .a ({signal_3577, signal_3569}), .c ({signal_1762, signal_842}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_30 ( .s (signal_3337), .b ({signal_1705, signal_744}), .a ({signal_3593, signal_3585}), .c ({signal_1764, signal_840}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_32 ( .s (signal_3337), .b ({signal_1715, signal_742}), .a ({signal_3609, signal_3601}), .c ({signal_1766, signal_806}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_34 ( .s (signal_3337), .b ({signal_1714, signal_740}), .a ({signal_3625, signal_3617}), .c ({signal_1768, signal_804}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_36 ( .s (signal_3337), .b ({signal_1713, signal_738}), .a ({signal_3641, signal_3633}), .c ({signal_1770, signal_802}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_38 ( .s (signal_3337), .b ({signal_1720, signal_736}), .a ({signal_3657, signal_3649}), .c ({signal_1772, signal_800}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_40 ( .s (signal_3337), .b ({signal_1721, signal_734}), .a ({signal_3673, signal_3665}), .c ({signal_1774, signal_798}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_42 ( .s (signal_3337), .b ({signal_1722, signal_732}), .a ({signal_3689, signal_3681}), .c ({signal_1776, signal_796}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_44 ( .s (signal_3337), .b ({signal_1723, signal_730}), .a ({signal_3705, signal_3697}), .c ({signal_1778, signal_794}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_46 ( .s (signal_3337), .b ({signal_1724, signal_728}), .a ({signal_3721, signal_3713}), .c ({signal_1780, signal_792}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_48 ( .s (signal_3337), .b ({signal_1725, signal_726}), .a ({signal_3737, signal_3729}), .c ({signal_1782, signal_790}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_50 ( .s (signal_3337), .b ({signal_1726, signal_724}), .a ({signal_3753, signal_3745}), .c ({signal_1784, signal_788}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_52 ( .s (signal_3337), .b ({signal_1727, signal_722}), .a ({signal_3769, signal_3761}), .c ({signal_1786, signal_786}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_54 ( .s (signal_3337), .b ({signal_1728, signal_720}), .a ({signal_3785, signal_3777}), .c ({signal_1788, signal_784}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_56 ( .s (signal_3337), .b ({signal_1729, signal_718}), .a ({signal_3801, signal_3793}), .c ({signal_1790, signal_782}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_58 ( .s (signal_3337), .b ({signal_1730, signal_716}), .a ({signal_3817, signal_3809}), .c ({signal_1792, signal_780}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_60 ( .s (signal_3337), .b ({signal_1731, signal_714}), .a ({signal_3833, signal_3825}), .c ({signal_1794, signal_778}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) cell_62 ( .s (signal_3337), .b ({signal_1732, signal_712}), .a ({signal_3849, signal_3841}), .c ({signal_1796, signal_776}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_64 ( .a ({signal_1846, signal_268}), .b ({signal_1845, signal_269}), .c ({signal_1917, signal_822}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_65 ( .a ({signal_1750, signal_854}), .b ({signal_1734, signal_870}), .c ({signal_1845, signal_269}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_66 ( .a ({1'b0, 1'b0}), .b ({signal_1782, signal_790}), .c ({signal_1846, signal_268}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_67 ( .a ({signal_1847, signal_270}), .b ({signal_1734, signal_870}), .c ({signal_1918, signal_838}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_68 ( .a ({1'b0, 1'b0}), .b ({signal_1766, signal_806}), .c ({signal_1847, signal_270}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_74 ( .a ({signal_1851, signal_274}), .b ({signal_1850, signal_275}), .c ({signal_1919, signal_820}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_75 ( .a ({signal_1752, signal_852}), .b ({signal_1736, signal_868}), .c ({signal_1850, signal_275}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_76 ( .a ({1'b0, 1'b0}), .b ({signal_1784, signal_788}), .c ({signal_1851, signal_274}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_77 ( .a ({signal_1852, signal_276}), .b ({signal_1736, signal_868}), .c ({signal_1920, signal_836}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_78 ( .a ({1'b0, 1'b0}), .b ({signal_1768, signal_804}), .c ({signal_1852, signal_276}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_84 ( .a ({signal_1856, signal_280}), .b ({signal_1855, signal_281}), .c ({signal_1921, signal_818}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_85 ( .a ({signal_1754, signal_850}), .b ({signal_1738, signal_866}), .c ({signal_1855, signal_281}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_86 ( .a ({1'b0, 1'b0}), .b ({signal_1786, signal_786}), .c ({signal_1856, signal_280}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_87 ( .a ({signal_1857, signal_282}), .b ({signal_1738, signal_866}), .c ({signal_1922, signal_834}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_88 ( .a ({1'b0, 1'b0}), .b ({signal_1770, signal_802}), .c ({signal_1857, signal_282}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_94 ( .a ({signal_1861, signal_286}), .b ({signal_1860, signal_287}), .c ({signal_1923, signal_816}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_95 ( .a ({signal_1756, signal_848}), .b ({signal_1740, signal_864}), .c ({signal_1860, signal_287}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_96 ( .a ({1'b0, 1'b0}), .b ({signal_1788, signal_784}), .c ({signal_1861, signal_286}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_97 ( .a ({signal_1862, signal_288}), .b ({signal_1740, signal_864}), .c ({signal_1924, signal_832}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_98 ( .a ({1'b0, 1'b0}), .b ({signal_1772, signal_800}), .c ({signal_1862, signal_288}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_104 ( .a ({signal_1866, signal_292}), .b ({signal_1865, signal_293}), .c ({signal_1925, signal_814}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_105 ( .a ({signal_1758, signal_846}), .b ({signal_1742, signal_862}), .c ({signal_1865, signal_293}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_106 ( .a ({1'b0, 1'b0}), .b ({signal_1790, signal_782}), .c ({signal_1866, signal_292}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_107 ( .a ({signal_1867, signal_294}), .b ({signal_1742, signal_862}), .c ({signal_1926, signal_830}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_108 ( .a ({1'b0, 1'b0}), .b ({signal_1774, signal_798}), .c ({signal_1867, signal_294}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_114 ( .a ({signal_1871, signal_298}), .b ({signal_1870, signal_299}), .c ({signal_1927, signal_812}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_115 ( .a ({signal_1760, signal_844}), .b ({signal_1744, signal_860}), .c ({signal_1870, signal_299}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_116 ( .a ({1'b0, 1'b0}), .b ({signal_1792, signal_780}), .c ({signal_1871, signal_298}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_117 ( .a ({signal_1872, signal_300}), .b ({signal_1744, signal_860}), .c ({signal_1928, signal_828}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_118 ( .a ({1'b0, 1'b0}), .b ({signal_1776, signal_796}), .c ({signal_1872, signal_300}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_124 ( .a ({signal_1876, signal_304}), .b ({signal_1875, signal_305}), .c ({signal_1929, signal_810}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_125 ( .a ({signal_1762, signal_842}), .b ({signal_1746, signal_858}), .c ({signal_1875, signal_305}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_126 ( .a ({1'b0, 1'b0}), .b ({signal_1794, signal_778}), .c ({signal_1876, signal_304}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_127 ( .a ({signal_1877, signal_306}), .b ({signal_1746, signal_858}), .c ({signal_1930, signal_826}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_128 ( .a ({1'b0, 1'b0}), .b ({signal_1778, signal_794}), .c ({signal_1877, signal_306}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_134 ( .a ({signal_1881, signal_310}), .b ({signal_1880, signal_311}), .c ({signal_1931, signal_808}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_135 ( .a ({signal_1764, signal_840}), .b ({signal_1748, signal_856}), .c ({signal_1880, signal_311}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_136 ( .a ({1'b0, 1'b0}), .b ({signal_1796, signal_776}), .c ({signal_1881, signal_310}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_137 ( .a ({signal_1882, signal_312}), .b ({signal_1748, signal_856}), .c ({signal_1932, signal_824}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_138 ( .a ({1'b0, 1'b0}), .b ({signal_1780, signal_792}), .c ({signal_1882, signal_312}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_144 ( .a ({signal_1965, signal_316}), .b ({signal_3865, signal_3857}), .c ({signal_1997, signal_950}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_145 ( .a ({1'b0, 1'b0}), .b ({signal_1917, signal_822}), .c ({signal_1965, signal_316}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_148 ( .a ({signal_1967, signal_318}), .b ({signal_3881, signal_3873}), .c ({signal_1998, signal_948}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_149 ( .a ({1'b0, 1'b0}), .b ({signal_1919, signal_820}), .c ({signal_1967, signal_318}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_152 ( .a ({signal_1969, signal_320}), .b ({signal_3897, signal_3889}), .c ({signal_1999, signal_946}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_153 ( .a ({1'b0, 1'b0}), .b ({signal_1921, signal_818}), .c ({signal_1969, signal_320}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_156 ( .a ({signal_1971, signal_322}), .b ({signal_3913, signal_3905}), .c ({signal_2000, signal_944}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_157 ( .a ({1'b0, 1'b0}), .b ({signal_1923, signal_816}), .c ({signal_1971, signal_322}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_160 ( .a ({signal_1973, signal_324}), .b ({signal_3929, signal_3921}), .c ({signal_2001, signal_942}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_161 ( .a ({1'b0, 1'b0}), .b ({signal_1925, signal_814}), .c ({signal_1973, signal_324}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_164 ( .a ({signal_1975, signal_326}), .b ({signal_3945, signal_3937}), .c ({signal_2002, signal_940}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_165 ( .a ({1'b0, 1'b0}), .b ({signal_1927, signal_812}), .c ({signal_1975, signal_326}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_168 ( .a ({signal_1977, signal_328}), .b ({signal_3961, signal_3953}), .c ({signal_2003, signal_938}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_169 ( .a ({1'b0, 1'b0}), .b ({signal_1929, signal_810}), .c ({signal_1977, signal_328}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_172 ( .a ({signal_1979, signal_330}), .b ({signal_3977, signal_3969}), .c ({signal_2004, signal_936}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_173 ( .a ({1'b0, 1'b0}), .b ({signal_1931, signal_808}), .c ({signal_1979, signal_330}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_176 ( .a ({signal_1981, signal_332}), .b ({signal_3993, signal_3985}), .c ({signal_2005, signal_958}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_178 ( .a ({1'b0, 1'b0}), .b ({signal_1926, signal_830}), .c ({signal_1981, signal_332}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_182 ( .a ({signal_1983, signal_336}), .b ({signal_4009, signal_4001}), .c ({signal_2006, signal_956}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_184 ( .a ({1'b0, 1'b0}), .b ({signal_1928, signal_828}), .c ({signal_1983, signal_336}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_188 ( .a ({signal_1985, signal_340}), .b ({signal_4025, signal_4017}), .c ({signal_2007, signal_954}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_190 ( .a ({1'b0, 1'b0}), .b ({signal_1930, signal_826}), .c ({signal_1985, signal_340}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_194 ( .a ({signal_1987, signal_344}), .b ({signal_4041, signal_4033}), .c ({signal_2008, signal_952}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_196 ( .a ({1'b0, 1'b0}), .b ({signal_1932, signal_824}), .c ({signal_1987, signal_344}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_200 ( .a ({signal_1885, signal_348}), .b ({signal_4057, signal_4049}), .c ({signal_1945, signal_998}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_201 ( .a ({1'b0, 1'b0}), .b ({signal_1734, signal_870}), .c ({signal_1885, signal_348}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_204 ( .a ({signal_1887, signal_350}), .b ({signal_4073, signal_4065}), .c ({signal_1946, signal_996}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_205 ( .a ({1'b0, 1'b0}), .b ({signal_1736, signal_868}), .c ({signal_1887, signal_350}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_208 ( .a ({signal_1889, signal_352}), .b ({signal_4089, signal_4081}), .c ({signal_1947, signal_994}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_209 ( .a ({1'b0, 1'b0}), .b ({signal_1738, signal_866}), .c ({signal_1889, signal_352}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_212 ( .a ({signal_1891, signal_354}), .b ({signal_4105, signal_4097}), .c ({signal_1948, signal_992}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_213 ( .a ({1'b0, 1'b0}), .b ({signal_1740, signal_864}), .c ({signal_1891, signal_354}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_216 ( .a ({signal_1893, signal_356}), .b ({signal_4121, signal_4113}), .c ({signal_1949, signal_990}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_217 ( .a ({1'b0, 1'b0}), .b ({signal_1742, signal_862}), .c ({signal_1893, signal_356}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_220 ( .a ({signal_1895, signal_358}), .b ({signal_4137, signal_4129}), .c ({signal_1950, signal_988}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_221 ( .a ({1'b0, 1'b0}), .b ({signal_1744, signal_860}), .c ({signal_1895, signal_358}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_224 ( .a ({signal_1897, signal_360}), .b ({signal_4153, signal_4145}), .c ({signal_1951, signal_986}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_225 ( .a ({1'b0, 1'b0}), .b ({signal_1746, signal_858}), .c ({signal_1897, signal_360}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_228 ( .a ({signal_1899, signal_362}), .b ({signal_4169, signal_4161}), .c ({signal_1952, signal_984}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_229 ( .a ({1'b0, 1'b0}), .b ({signal_1748, signal_856}), .c ({signal_1899, signal_362}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_232 ( .a ({signal_1901, signal_364}), .b ({signal_4185, signal_4177}), .c ({signal_1953, signal_982}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_233 ( .a ({1'b0, 1'b0}), .b ({signal_1750, signal_854}), .c ({signal_1901, signal_364}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_236 ( .a ({signal_1903, signal_366}), .b ({signal_4201, signal_4193}), .c ({signal_1954, signal_980}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_237 ( .a ({1'b0, 1'b0}), .b ({signal_1752, signal_852}), .c ({signal_1903, signal_366}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_240 ( .a ({signal_1905, signal_368}), .b ({signal_4217, signal_4209}), .c ({signal_1955, signal_978}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_241 ( .a ({1'b0, 1'b0}), .b ({signal_1754, signal_850}), .c ({signal_1905, signal_368}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_244 ( .a ({signal_1907, signal_370}), .b ({signal_4233, signal_4225}), .c ({signal_1956, signal_976}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_245 ( .a ({1'b0, 1'b0}), .b ({signal_1756, signal_848}), .c ({signal_1907, signal_370}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_248 ( .a ({signal_1909, signal_372}), .b ({signal_4249, signal_4241}), .c ({signal_1957, signal_974}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_249 ( .a ({1'b0, 1'b0}), .b ({signal_1758, signal_846}), .c ({signal_1909, signal_372}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_252 ( .a ({signal_1911, signal_374}), .b ({signal_4265, signal_4257}), .c ({signal_1958, signal_972}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_253 ( .a ({1'b0, 1'b0}), .b ({signal_1760, signal_844}), .c ({signal_1911, signal_374}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_256 ( .a ({signal_1913, signal_376}), .b ({signal_4281, signal_4273}), .c ({signal_1959, signal_970}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_257 ( .a ({1'b0, 1'b0}), .b ({signal_1762, signal_842}), .c ({signal_1913, signal_376}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_260 ( .a ({signal_1915, signal_378}), .b ({signal_4297, signal_4289}), .c ({signal_1960, signal_968}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_261 ( .a ({1'b0, 1'b0}), .b ({signal_1764, signal_840}), .c ({signal_1915, signal_378}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_264 ( .a ({signal_1989, signal_380}), .b ({signal_4313, signal_4305}), .c ({signal_2009, signal_966}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_265 ( .a ({1'b0, 1'b0}), .b ({signal_1918, signal_838}), .c ({signal_1989, signal_380}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_268 ( .a ({signal_1991, signal_382}), .b ({signal_4329, signal_4321}), .c ({signal_2010, signal_964}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_269 ( .a ({1'b0, 1'b0}), .b ({signal_1920, signal_836}), .c ({signal_1991, signal_382}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_272 ( .a ({signal_1993, signal_384}), .b ({signal_4345, signal_4337}), .c ({signal_2011, signal_962}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_273 ( .a ({1'b0, 1'b0}), .b ({signal_1922, signal_834}), .c ({signal_1993, signal_384}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_276 ( .a ({signal_1995, signal_386}), .b ({signal_4361, signal_4353}), .c ({signal_2012, signal_960}) ) ;
    xnor_HPC2 #(.security_order(1), .pipeline(1)) cell_277 ( .a ({1'b0, 1'b0}), .b ({signal_1924, signal_832}), .c ({signal_1995, signal_386}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1016 ( .s ({signal_4365, signal_4363}), .b ({signal_4369, signal_4367}), .a ({signal_1435, signal_1162}), .clk (clk), .r (Fresh[197]), .c ({signal_1701, signal_756}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1017 ( .s ({signal_4373, signal_4371}), .b ({signal_1458, signal_1169}), .a ({signal_4377, signal_4375}), .clk (clk), .r (Fresh[198]), .c ({signal_1702, signal_754}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1018 ( .s ({signal_4381, signal_4379}), .b ({signal_1449, signal_1167}), .a ({signal_4385, signal_4383}), .clk (clk), .r (Fresh[199]), .c ({signal_1703, signal_746}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1019 ( .s ({signal_4389, signal_4387}), .b ({signal_4393, signal_4391}), .a ({signal_1462, signal_1171}), .clk (clk), .r (Fresh[200]), .c ({signal_1704, signal_748}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1020 ( .s ({signal_4381, signal_4379}), .b ({signal_4397, signal_4395}), .a ({signal_1424, signal_1158}), .clk (clk), .r (Fresh[201]), .c ({signal_1705, signal_744}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1021 ( .s ({signal_4365, signal_4363}), .b ({signal_1430, signal_1160}), .a ({signal_4401, signal_4399}), .clk (clk), .r (Fresh[202]), .c ({signal_1706, signal_758}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1022 ( .s ({signal_4405, signal_4403}), .b ({signal_4409, signal_4407}), .a ({signal_1437, signal_1164}), .clk (clk), .r (Fresh[203]), .c ({signal_1707, signal_772}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1023 ( .s ({signal_4405, signal_4403}), .b ({signal_1417, signal_1154}), .a ({signal_4413, signal_4411}), .clk (clk), .r (Fresh[204]), .c ({signal_1708, signal_774}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1024 ( .s ({signal_4417, signal_4415}), .b ({signal_4421, signal_4419}), .a ({signal_1459, signal_1170}), .clk (clk), .r (Fresh[205]), .c ({signal_1709, signal_760}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1025 ( .s ({signal_4389, signal_4387}), .b ({signal_1422, signal_1156}), .a ({signal_4425, signal_4423}), .clk (clk), .r (Fresh[206]), .c ({signal_1710, signal_750}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1026 ( .s ({signal_4429, signal_4427}), .b ({signal_4433, signal_4431}), .a ({signal_1441, signal_1165}), .clk (clk), .r (Fresh[207]), .c ({signal_1711, signal_768}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1027 ( .s ({signal_4437, signal_4435}), .b ({signal_4441, signal_4439}), .a ({signal_1436, signal_1163}), .clk (clk), .r (Fresh[208]), .c ({signal_1712, signal_764}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1028 ( .s ({signal_4445, signal_4443}), .b ({signal_1416, signal_1153}), .a ({signal_4449, signal_4447}), .clk (clk), .r (Fresh[209]), .c ({signal_1713, signal_738}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1029 ( .s ({signal_4453, signal_4451}), .b ({signal_4457, signal_4455}), .a ({signal_1455, signal_1168}), .clk (clk), .r (Fresh[210]), .c ({signal_1714, signal_740}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1030 ( .s ({signal_4453, signal_4451}), .b ({signal_1431, signal_1161}), .a ({signal_4461, signal_4459}), .clk (clk), .r (Fresh[211]), .c ({signal_1715, signal_742}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1031 ( .s ({signal_4373, signal_4371}), .b ({signal_4465, signal_4463}), .a ({signal_1423, signal_1157}), .clk (clk), .r (Fresh[212]), .c ({signal_1716, signal_752}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1032 ( .s ({signal_4429, signal_4427}), .b ({signal_1419, signal_1155}), .a ({signal_4469, signal_4467}), .clk (clk), .r (Fresh[213]), .c ({signal_1717, signal_770}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1033 ( .s ({signal_4417, signal_4415}), .b ({signal_1444, signal_1166}), .a ({signal_4473, signal_4471}), .clk (clk), .r (Fresh[214]), .c ({signal_1718, signal_762}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1034 ( .s ({signal_4437, signal_4435}), .b ({signal_1425, signal_1159}), .a ({signal_4477, signal_4475}), .clk (clk), .r (Fresh[215]), .c ({signal_1719, signal_766}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1035 ( .s ({signal_4445, signal_4443}), .b ({signal_4481, signal_4479}), .a ({signal_1413, signal_1152}), .clk (clk), .r (Fresh[216]), .c ({signal_1720, signal_736}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1036 ( .s ({signal_4485, signal_4483}), .b ({signal_1463, signal_1172}), .a ({signal_4489, signal_4487}), .clk (clk), .r (Fresh[217]), .c ({signal_1721, signal_734}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1037 ( .s ({signal_4485, signal_4483}), .b ({signal_4493, signal_4491}), .a ({signal_1465, signal_1173}), .clk (clk), .r (Fresh[218]), .c ({signal_1722, signal_732}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1038 ( .s ({signal_4497, signal_4495}), .b ({signal_1468, signal_1174}), .a ({signal_4501, signal_4499}), .clk (clk), .r (Fresh[219]), .c ({signal_1723, signal_730}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1039 ( .s ({signal_4497, signal_4495}), .b ({signal_4505, signal_4503}), .a ({signal_1470, signal_1175}), .clk (clk), .r (Fresh[220]), .c ({signal_1724, signal_728}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1040 ( .s ({signal_4509, signal_4507}), .b ({signal_1473, signal_1176}), .a ({signal_4513, signal_4511}), .clk (clk), .r (Fresh[221]), .c ({signal_1725, signal_726}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1041 ( .s ({signal_4509, signal_4507}), .b ({signal_4517, signal_4515}), .a ({signal_1475, signal_1177}), .clk (clk), .r (Fresh[222]), .c ({signal_1726, signal_724}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1042 ( .s ({signal_4521, signal_4519}), .b ({signal_1478, signal_1178}), .a ({signal_4525, signal_4523}), .clk (clk), .r (Fresh[223]), .c ({signal_1727, signal_722}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1043 ( .s ({signal_4521, signal_4519}), .b ({signal_4529, signal_4527}), .a ({signal_1480, signal_1179}), .clk (clk), .r (Fresh[224]), .c ({signal_1728, signal_720}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1044 ( .s ({signal_4533, signal_4531}), .b ({signal_1483, signal_1180}), .a ({signal_4537, signal_4535}), .clk (clk), .r (Fresh[225]), .c ({signal_1729, signal_718}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1045 ( .s ({signal_4533, signal_4531}), .b ({signal_4541, signal_4539}), .a ({signal_1485, signal_1181}), .clk (clk), .r (Fresh[226]), .c ({signal_1730, signal_716}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1046 ( .s ({signal_4545, signal_4543}), .b ({signal_1488, signal_1182}), .a ({signal_4549, signal_4547}), .clk (clk), .r (Fresh[227]), .c ({signal_1731, signal_714}) ) ;
    mux2_HPC2 #(.security_order(1), .pipeline(1)) cell_1047 ( .s ({signal_4545, signal_4543}), .b ({signal_4553, signal_4551}), .a ({signal_1490, signal_1183}), .clk (clk), .r (Fresh[228]), .c ({signal_1732, signal_712}) ) ;
    buf_clk cell_2143 ( .C (clk), .D (signal_3336), .Q (signal_3337) ) ;
    buf_clk cell_2151 ( .C (clk), .D (signal_3344), .Q (signal_3345) ) ;
    buf_clk cell_2159 ( .C (clk), .D (signal_3352), .Q (signal_3353) ) ;
    buf_clk cell_2167 ( .C (clk), .D (signal_3360), .Q (signal_3361) ) ;
    buf_clk cell_2175 ( .C (clk), .D (signal_3368), .Q (signal_3369) ) ;
    buf_clk cell_2183 ( .C (clk), .D (signal_3376), .Q (signal_3377) ) ;
    buf_clk cell_2191 ( .C (clk), .D (signal_3384), .Q (signal_3385) ) ;
    buf_clk cell_2199 ( .C (clk), .D (signal_3392), .Q (signal_3393) ) ;
    buf_clk cell_2207 ( .C (clk), .D (signal_3400), .Q (signal_3401) ) ;
    buf_clk cell_2215 ( .C (clk), .D (signal_3408), .Q (signal_3409) ) ;
    buf_clk cell_2223 ( .C (clk), .D (signal_3416), .Q (signal_3417) ) ;
    buf_clk cell_2231 ( .C (clk), .D (signal_3424), .Q (signal_3425) ) ;
    buf_clk cell_2239 ( .C (clk), .D (signal_3432), .Q (signal_3433) ) ;
    buf_clk cell_2247 ( .C (clk), .D (signal_3440), .Q (signal_3441) ) ;
    buf_clk cell_2255 ( .C (clk), .D (signal_3448), .Q (signal_3449) ) ;
    buf_clk cell_2263 ( .C (clk), .D (signal_3456), .Q (signal_3457) ) ;
    buf_clk cell_2271 ( .C (clk), .D (signal_3464), .Q (signal_3465) ) ;
    buf_clk cell_2279 ( .C (clk), .D (signal_3472), .Q (signal_3473) ) ;
    buf_clk cell_2287 ( .C (clk), .D (signal_3480), .Q (signal_3481) ) ;
    buf_clk cell_2295 ( .C (clk), .D (signal_3488), .Q (signal_3489) ) ;
    buf_clk cell_2303 ( .C (clk), .D (signal_3496), .Q (signal_3497) ) ;
    buf_clk cell_2311 ( .C (clk), .D (signal_3504), .Q (signal_3505) ) ;
    buf_clk cell_2319 ( .C (clk), .D (signal_3512), .Q (signal_3513) ) ;
    buf_clk cell_2327 ( .C (clk), .D (signal_3520), .Q (signal_3521) ) ;
    buf_clk cell_2335 ( .C (clk), .D (signal_3528), .Q (signal_3529) ) ;
    buf_clk cell_2343 ( .C (clk), .D (signal_3536), .Q (signal_3537) ) ;
    buf_clk cell_2351 ( .C (clk), .D (signal_3544), .Q (signal_3545) ) ;
    buf_clk cell_2359 ( .C (clk), .D (signal_3552), .Q (signal_3553) ) ;
    buf_clk cell_2367 ( .C (clk), .D (signal_3560), .Q (signal_3561) ) ;
    buf_clk cell_2375 ( .C (clk), .D (signal_3568), .Q (signal_3569) ) ;
    buf_clk cell_2383 ( .C (clk), .D (signal_3576), .Q (signal_3577) ) ;
    buf_clk cell_2391 ( .C (clk), .D (signal_3584), .Q (signal_3585) ) ;
    buf_clk cell_2399 ( .C (clk), .D (signal_3592), .Q (signal_3593) ) ;
    buf_clk cell_2407 ( .C (clk), .D (signal_3600), .Q (signal_3601) ) ;
    buf_clk cell_2415 ( .C (clk), .D (signal_3608), .Q (signal_3609) ) ;
    buf_clk cell_2423 ( .C (clk), .D (signal_3616), .Q (signal_3617) ) ;
    buf_clk cell_2431 ( .C (clk), .D (signal_3624), .Q (signal_3625) ) ;
    buf_clk cell_2439 ( .C (clk), .D (signal_3632), .Q (signal_3633) ) ;
    buf_clk cell_2447 ( .C (clk), .D (signal_3640), .Q (signal_3641) ) ;
    buf_clk cell_2455 ( .C (clk), .D (signal_3648), .Q (signal_3649) ) ;
    buf_clk cell_2463 ( .C (clk), .D (signal_3656), .Q (signal_3657) ) ;
    buf_clk cell_2471 ( .C (clk), .D (signal_3664), .Q (signal_3665) ) ;
    buf_clk cell_2479 ( .C (clk), .D (signal_3672), .Q (signal_3673) ) ;
    buf_clk cell_2487 ( .C (clk), .D (signal_3680), .Q (signal_3681) ) ;
    buf_clk cell_2495 ( .C (clk), .D (signal_3688), .Q (signal_3689) ) ;
    buf_clk cell_2503 ( .C (clk), .D (signal_3696), .Q (signal_3697) ) ;
    buf_clk cell_2511 ( .C (clk), .D (signal_3704), .Q (signal_3705) ) ;
    buf_clk cell_2519 ( .C (clk), .D (signal_3712), .Q (signal_3713) ) ;
    buf_clk cell_2527 ( .C (clk), .D (signal_3720), .Q (signal_3721) ) ;
    buf_clk cell_2535 ( .C (clk), .D (signal_3728), .Q (signal_3729) ) ;
    buf_clk cell_2543 ( .C (clk), .D (signal_3736), .Q (signal_3737) ) ;
    buf_clk cell_2551 ( .C (clk), .D (signal_3744), .Q (signal_3745) ) ;
    buf_clk cell_2559 ( .C (clk), .D (signal_3752), .Q (signal_3753) ) ;
    buf_clk cell_2567 ( .C (clk), .D (signal_3760), .Q (signal_3761) ) ;
    buf_clk cell_2575 ( .C (clk), .D (signal_3768), .Q (signal_3769) ) ;
    buf_clk cell_2583 ( .C (clk), .D (signal_3776), .Q (signal_3777) ) ;
    buf_clk cell_2591 ( .C (clk), .D (signal_3784), .Q (signal_3785) ) ;
    buf_clk cell_2599 ( .C (clk), .D (signal_3792), .Q (signal_3793) ) ;
    buf_clk cell_2607 ( .C (clk), .D (signal_3800), .Q (signal_3801) ) ;
    buf_clk cell_2615 ( .C (clk), .D (signal_3808), .Q (signal_3809) ) ;
    buf_clk cell_2623 ( .C (clk), .D (signal_3816), .Q (signal_3817) ) ;
    buf_clk cell_2631 ( .C (clk), .D (signal_3824), .Q (signal_3825) ) ;
    buf_clk cell_2639 ( .C (clk), .D (signal_3832), .Q (signal_3833) ) ;
    buf_clk cell_2647 ( .C (clk), .D (signal_3840), .Q (signal_3841) ) ;
    buf_clk cell_2655 ( .C (clk), .D (signal_3848), .Q (signal_3849) ) ;
    buf_clk cell_2663 ( .C (clk), .D (signal_3856), .Q (signal_3857) ) ;
    buf_clk cell_2671 ( .C (clk), .D (signal_3864), .Q (signal_3865) ) ;
    buf_clk cell_2679 ( .C (clk), .D (signal_3872), .Q (signal_3873) ) ;
    buf_clk cell_2687 ( .C (clk), .D (signal_3880), .Q (signal_3881) ) ;
    buf_clk cell_2695 ( .C (clk), .D (signal_3888), .Q (signal_3889) ) ;
    buf_clk cell_2703 ( .C (clk), .D (signal_3896), .Q (signal_3897) ) ;
    buf_clk cell_2711 ( .C (clk), .D (signal_3904), .Q (signal_3905) ) ;
    buf_clk cell_2719 ( .C (clk), .D (signal_3912), .Q (signal_3913) ) ;
    buf_clk cell_2727 ( .C (clk), .D (signal_3920), .Q (signal_3921) ) ;
    buf_clk cell_2735 ( .C (clk), .D (signal_3928), .Q (signal_3929) ) ;
    buf_clk cell_2743 ( .C (clk), .D (signal_3936), .Q (signal_3937) ) ;
    buf_clk cell_2751 ( .C (clk), .D (signal_3944), .Q (signal_3945) ) ;
    buf_clk cell_2759 ( .C (clk), .D (signal_3952), .Q (signal_3953) ) ;
    buf_clk cell_2767 ( .C (clk), .D (signal_3960), .Q (signal_3961) ) ;
    buf_clk cell_2775 ( .C (clk), .D (signal_3968), .Q (signal_3969) ) ;
    buf_clk cell_2783 ( .C (clk), .D (signal_3976), .Q (signal_3977) ) ;
    buf_clk cell_2791 ( .C (clk), .D (signal_3984), .Q (signal_3985) ) ;
    buf_clk cell_2799 ( .C (clk), .D (signal_3992), .Q (signal_3993) ) ;
    buf_clk cell_2807 ( .C (clk), .D (signal_4000), .Q (signal_4001) ) ;
    buf_clk cell_2815 ( .C (clk), .D (signal_4008), .Q (signal_4009) ) ;
    buf_clk cell_2823 ( .C (clk), .D (signal_4016), .Q (signal_4017) ) ;
    buf_clk cell_2831 ( .C (clk), .D (signal_4024), .Q (signal_4025) ) ;
    buf_clk cell_2839 ( .C (clk), .D (signal_4032), .Q (signal_4033) ) ;
    buf_clk cell_2847 ( .C (clk), .D (signal_4040), .Q (signal_4041) ) ;
    buf_clk cell_2855 ( .C (clk), .D (signal_4048), .Q (signal_4049) ) ;
    buf_clk cell_2863 ( .C (clk), .D (signal_4056), .Q (signal_4057) ) ;
    buf_clk cell_2871 ( .C (clk), .D (signal_4064), .Q (signal_4065) ) ;
    buf_clk cell_2879 ( .C (clk), .D (signal_4072), .Q (signal_4073) ) ;
    buf_clk cell_2887 ( .C (clk), .D (signal_4080), .Q (signal_4081) ) ;
    buf_clk cell_2895 ( .C (clk), .D (signal_4088), .Q (signal_4089) ) ;
    buf_clk cell_2903 ( .C (clk), .D (signal_4096), .Q (signal_4097) ) ;
    buf_clk cell_2911 ( .C (clk), .D (signal_4104), .Q (signal_4105) ) ;
    buf_clk cell_2919 ( .C (clk), .D (signal_4112), .Q (signal_4113) ) ;
    buf_clk cell_2927 ( .C (clk), .D (signal_4120), .Q (signal_4121) ) ;
    buf_clk cell_2935 ( .C (clk), .D (signal_4128), .Q (signal_4129) ) ;
    buf_clk cell_2943 ( .C (clk), .D (signal_4136), .Q (signal_4137) ) ;
    buf_clk cell_2951 ( .C (clk), .D (signal_4144), .Q (signal_4145) ) ;
    buf_clk cell_2959 ( .C (clk), .D (signal_4152), .Q (signal_4153) ) ;
    buf_clk cell_2967 ( .C (clk), .D (signal_4160), .Q (signal_4161) ) ;
    buf_clk cell_2975 ( .C (clk), .D (signal_4168), .Q (signal_4169) ) ;
    buf_clk cell_2983 ( .C (clk), .D (signal_4176), .Q (signal_4177) ) ;
    buf_clk cell_2991 ( .C (clk), .D (signal_4184), .Q (signal_4185) ) ;
    buf_clk cell_2999 ( .C (clk), .D (signal_4192), .Q (signal_4193) ) ;
    buf_clk cell_3007 ( .C (clk), .D (signal_4200), .Q (signal_4201) ) ;
    buf_clk cell_3015 ( .C (clk), .D (signal_4208), .Q (signal_4209) ) ;
    buf_clk cell_3023 ( .C (clk), .D (signal_4216), .Q (signal_4217) ) ;
    buf_clk cell_3031 ( .C (clk), .D (signal_4224), .Q (signal_4225) ) ;
    buf_clk cell_3039 ( .C (clk), .D (signal_4232), .Q (signal_4233) ) ;
    buf_clk cell_3047 ( .C (clk), .D (signal_4240), .Q (signal_4241) ) ;
    buf_clk cell_3055 ( .C (clk), .D (signal_4248), .Q (signal_4249) ) ;
    buf_clk cell_3063 ( .C (clk), .D (signal_4256), .Q (signal_4257) ) ;
    buf_clk cell_3071 ( .C (clk), .D (signal_4264), .Q (signal_4265) ) ;
    buf_clk cell_3079 ( .C (clk), .D (signal_4272), .Q (signal_4273) ) ;
    buf_clk cell_3087 ( .C (clk), .D (signal_4280), .Q (signal_4281) ) ;
    buf_clk cell_3095 ( .C (clk), .D (signal_4288), .Q (signal_4289) ) ;
    buf_clk cell_3103 ( .C (clk), .D (signal_4296), .Q (signal_4297) ) ;
    buf_clk cell_3111 ( .C (clk), .D (signal_4304), .Q (signal_4305) ) ;
    buf_clk cell_3119 ( .C (clk), .D (signal_4312), .Q (signal_4313) ) ;
    buf_clk cell_3127 ( .C (clk), .D (signal_4320), .Q (signal_4321) ) ;
    buf_clk cell_3135 ( .C (clk), .D (signal_4328), .Q (signal_4329) ) ;
    buf_clk cell_3143 ( .C (clk), .D (signal_4336), .Q (signal_4337) ) ;
    buf_clk cell_3151 ( .C (clk), .D (signal_4344), .Q (signal_4345) ) ;
    buf_clk cell_3159 ( .C (clk), .D (signal_4352), .Q (signal_4353) ) ;
    buf_clk cell_3167 ( .C (clk), .D (signal_4360), .Q (signal_4361) ) ;
    buf_clk cell_3361 ( .C (clk), .D (signal_4554), .Q (signal_4555) ) ;
    buf_clk cell_3363 ( .C (clk), .D (signal_4556), .Q (signal_4557) ) ;
    buf_clk cell_3365 ( .C (clk), .D (signal_4558), .Q (signal_4559) ) ;
    buf_clk cell_3367 ( .C (clk), .D (signal_4560), .Q (signal_4561) ) ;
    buf_clk cell_3369 ( .C (clk), .D (signal_4562), .Q (signal_4563) ) ;
    buf_clk cell_3371 ( .C (clk), .D (signal_4564), .Q (signal_4565) ) ;
    buf_clk cell_3373 ( .C (clk), .D (signal_4566), .Q (signal_4567) ) ;
    buf_clk cell_3375 ( .C (clk), .D (signal_4568), .Q (signal_4569) ) ;
    buf_clk cell_3377 ( .C (clk), .D (signal_4570), .Q (signal_4571) ) ;
    buf_clk cell_3379 ( .C (clk), .D (signal_4572), .Q (signal_4573) ) ;
    buf_clk cell_3381 ( .C (clk), .D (signal_4574), .Q (signal_4575) ) ;
    buf_clk cell_3383 ( .C (clk), .D (signal_4576), .Q (signal_4577) ) ;
    buf_clk cell_3385 ( .C (clk), .D (signal_4578), .Q (signal_4579) ) ;
    buf_clk cell_3387 ( .C (clk), .D (signal_4580), .Q (signal_4581) ) ;
    buf_clk cell_3389 ( .C (clk), .D (signal_4582), .Q (signal_4583) ) ;
    buf_clk cell_3391 ( .C (clk), .D (signal_4584), .Q (signal_4585) ) ;
    buf_clk cell_3393 ( .C (clk), .D (signal_4586), .Q (signal_4587) ) ;
    buf_clk cell_3395 ( .C (clk), .D (signal_4588), .Q (signal_4589) ) ;
    buf_clk cell_3397 ( .C (clk), .D (signal_4590), .Q (signal_4591) ) ;
    buf_clk cell_3399 ( .C (clk), .D (signal_4592), .Q (signal_4593) ) ;
    buf_clk cell_3401 ( .C (clk), .D (signal_4594), .Q (signal_4595) ) ;
    buf_clk cell_3403 ( .C (clk), .D (signal_4596), .Q (signal_4597) ) ;
    buf_clk cell_3405 ( .C (clk), .D (signal_4598), .Q (signal_4599) ) ;
    buf_clk cell_3407 ( .C (clk), .D (signal_4600), .Q (signal_4601) ) ;
    buf_clk cell_3409 ( .C (clk), .D (signal_4602), .Q (signal_4603) ) ;
    buf_clk cell_3411 ( .C (clk), .D (signal_4604), .Q (signal_4605) ) ;
    buf_clk cell_3413 ( .C (clk), .D (signal_4606), .Q (signal_4607) ) ;
    buf_clk cell_3415 ( .C (clk), .D (signal_4608), .Q (signal_4609) ) ;
    buf_clk cell_3417 ( .C (clk), .D (signal_4610), .Q (signal_4611) ) ;
    buf_clk cell_3419 ( .C (clk), .D (signal_4612), .Q (signal_4613) ) ;
    buf_clk cell_3421 ( .C (clk), .D (signal_4614), .Q (signal_4615) ) ;
    buf_clk cell_3423 ( .C (clk), .D (signal_4616), .Q (signal_4617) ) ;
    buf_clk cell_3425 ( .C (clk), .D (signal_4618), .Q (signal_4619) ) ;
    buf_clk cell_3427 ( .C (clk), .D (signal_4620), .Q (signal_4621) ) ;
    buf_clk cell_3429 ( .C (clk), .D (signal_4622), .Q (signal_4623) ) ;
    buf_clk cell_3431 ( .C (clk), .D (signal_4624), .Q (signal_4625) ) ;
    buf_clk cell_3433 ( .C (clk), .D (signal_4626), .Q (signal_4627) ) ;
    buf_clk cell_3435 ( .C (clk), .D (signal_4628), .Q (signal_4629) ) ;
    buf_clk cell_3437 ( .C (clk), .D (signal_4630), .Q (signal_4631) ) ;
    buf_clk cell_3439 ( .C (clk), .D (signal_4632), .Q (signal_4633) ) ;
    buf_clk cell_3441 ( .C (clk), .D (signal_4634), .Q (signal_4635) ) ;
    buf_clk cell_3443 ( .C (clk), .D (signal_4636), .Q (signal_4637) ) ;
    buf_clk cell_3445 ( .C (clk), .D (signal_4638), .Q (signal_4639) ) ;
    buf_clk cell_3447 ( .C (clk), .D (signal_4640), .Q (signal_4641) ) ;
    buf_clk cell_3449 ( .C (clk), .D (signal_4642), .Q (signal_4643) ) ;
    buf_clk cell_3451 ( .C (clk), .D (signal_4644), .Q (signal_4645) ) ;
    buf_clk cell_3453 ( .C (clk), .D (signal_4646), .Q (signal_4647) ) ;
    buf_clk cell_3455 ( .C (clk), .D (signal_4648), .Q (signal_4649) ) ;
    buf_clk cell_3457 ( .C (clk), .D (signal_4650), .Q (signal_4651) ) ;
    buf_clk cell_3459 ( .C (clk), .D (signal_4652), .Q (signal_4653) ) ;
    buf_clk cell_3461 ( .C (clk), .D (signal_4654), .Q (signal_4655) ) ;
    buf_clk cell_3463 ( .C (clk), .D (signal_4656), .Q (signal_4657) ) ;
    buf_clk cell_3465 ( .C (clk), .D (signal_4658), .Q (signal_4659) ) ;
    buf_clk cell_3467 ( .C (clk), .D (signal_4660), .Q (signal_4661) ) ;
    buf_clk cell_3469 ( .C (clk), .D (signal_4662), .Q (signal_4663) ) ;
    buf_clk cell_3471 ( .C (clk), .D (signal_4664), .Q (signal_4665) ) ;
    buf_clk cell_3473 ( .C (clk), .D (signal_4666), .Q (signal_4667) ) ;
    buf_clk cell_3475 ( .C (clk), .D (signal_4668), .Q (signal_4669) ) ;
    buf_clk cell_3477 ( .C (clk), .D (signal_4670), .Q (signal_4671) ) ;
    buf_clk cell_3479 ( .C (clk), .D (signal_4672), .Q (signal_4673) ) ;
    buf_clk cell_3481 ( .C (clk), .D (signal_4674), .Q (signal_4675) ) ;
    buf_clk cell_3483 ( .C (clk), .D (signal_4676), .Q (signal_4677) ) ;
    buf_clk cell_3485 ( .C (clk), .D (signal_4678), .Q (signal_4679) ) ;
    buf_clk cell_3487 ( .C (clk), .D (signal_4680), .Q (signal_4681) ) ;
    buf_clk cell_3495 ( .C (clk), .D (signal_4688), .Q (signal_4689) ) ;
    buf_clk cell_3503 ( .C (clk), .D (signal_4696), .Q (signal_4697) ) ;
    buf_clk cell_3511 ( .C (clk), .D (signal_4704), .Q (signal_4705) ) ;
    buf_clk cell_3519 ( .C (clk), .D (signal_4712), .Q (signal_4713) ) ;
    buf_clk cell_3527 ( .C (clk), .D (signal_4720), .Q (signal_4721) ) ;
    buf_clk cell_3535 ( .C (clk), .D (signal_4728), .Q (signal_4729) ) ;
    buf_clk cell_3543 ( .C (clk), .D (signal_4736), .Q (signal_4737) ) ;
    buf_clk cell_3551 ( .C (clk), .D (signal_4744), .Q (signal_4745) ) ;
    buf_clk cell_3559 ( .C (clk), .D (signal_4752), .Q (signal_4753) ) ;
    buf_clk cell_3567 ( .C (clk), .D (signal_4760), .Q (signal_4761) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_281 ( .clk (clk), .D ({signal_4557, signal_4555}), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_283 ( .clk (clk), .D ({signal_2004, signal_936}), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_285 ( .clk (clk), .D ({signal_4561, signal_4559}), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_287 ( .clk (clk), .D ({signal_2003, signal_938}), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_289 ( .clk (clk), .D ({signal_4565, signal_4563}), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_291 ( .clk (clk), .D ({signal_2002, signal_940}), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_293 ( .clk (clk), .D ({signal_4569, signal_4567}), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_295 ( .clk (clk), .D ({signal_2001, signal_942}), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_297 ( .clk (clk), .D ({signal_4573, signal_4571}), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_299 ( .clk (clk), .D ({signal_2000, signal_944}), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_301 ( .clk (clk), .D ({signal_4577, signal_4575}), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_303 ( .clk (clk), .D ({signal_1999, signal_946}), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_305 ( .clk (clk), .D ({signal_4581, signal_4579}), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_307 ( .clk (clk), .D ({signal_1998, signal_948}), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_309 ( .clk (clk), .D ({signal_4585, signal_4583}), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_311 ( .clk (clk), .D ({signal_1997, signal_950}), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_313 ( .clk (clk), .D ({signal_4589, signal_4587}), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_315 ( .clk (clk), .D ({signal_2008, signal_952}), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_317 ( .clk (clk), .D ({signal_4593, signal_4591}), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_319 ( .clk (clk), .D ({signal_2007, signal_954}), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_321 ( .clk (clk), .D ({signal_4597, signal_4595}), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_323 ( .clk (clk), .D ({signal_2006, signal_956}), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_325 ( .clk (clk), .D ({signal_4601, signal_4599}), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_327 ( .clk (clk), .D ({signal_2005, signal_958}), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_329 ( .clk (clk), .D ({signal_4605, signal_4603}), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_331 ( .clk (clk), .D ({signal_2012, signal_960}), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_333 ( .clk (clk), .D ({signal_4609, signal_4607}), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_335 ( .clk (clk), .D ({signal_2011, signal_962}), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_337 ( .clk (clk), .D ({signal_4613, signal_4611}), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_339 ( .clk (clk), .D ({signal_2010, signal_964}), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_341 ( .clk (clk), .D ({signal_4617, signal_4615}), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_343 ( .clk (clk), .D ({signal_2009, signal_966}), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_345 ( .clk (clk), .D ({signal_4621, signal_4619}), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_347 ( .clk (clk), .D ({signal_1960, signal_968}), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_349 ( .clk (clk), .D ({signal_4625, signal_4623}), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_351 ( .clk (clk), .D ({signal_1959, signal_970}), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_353 ( .clk (clk), .D ({signal_4629, signal_4627}), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_355 ( .clk (clk), .D ({signal_1958, signal_972}), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_357 ( .clk (clk), .D ({signal_4633, signal_4631}), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_359 ( .clk (clk), .D ({signal_1957, signal_974}), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_361 ( .clk (clk), .D ({signal_4637, signal_4635}), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_363 ( .clk (clk), .D ({signal_1956, signal_976}), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_365 ( .clk (clk), .D ({signal_4641, signal_4639}), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_367 ( .clk (clk), .D ({signal_1955, signal_978}), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_369 ( .clk (clk), .D ({signal_4645, signal_4643}), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_371 ( .clk (clk), .D ({signal_1954, signal_980}), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_373 ( .clk (clk), .D ({signal_4649, signal_4647}), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_375 ( .clk (clk), .D ({signal_1953, signal_982}), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_377 ( .clk (clk), .D ({signal_4653, signal_4651}), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_379 ( .clk (clk), .D ({signal_1952, signal_984}), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_381 ( .clk (clk), .D ({signal_4657, signal_4655}), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_383 ( .clk (clk), .D ({signal_1951, signal_986}), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_385 ( .clk (clk), .D ({signal_4661, signal_4659}), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_387 ( .clk (clk), .D ({signal_1950, signal_988}), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_389 ( .clk (clk), .D ({signal_4665, signal_4663}), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_391 ( .clk (clk), .D ({signal_1949, signal_990}), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_393 ( .clk (clk), .D ({signal_4669, signal_4667}), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_395 ( .clk (clk), .D ({signal_1948, signal_992}), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_397 ( .clk (clk), .D ({signal_4673, signal_4671}), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_399 ( .clk (clk), .D ({signal_1947, signal_994}), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_401 ( .clk (clk), .D ({signal_4677, signal_4675}), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_403 ( .clk (clk), .D ({signal_1946, signal_996}), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_405 ( .clk (clk), .D ({signal_4681, signal_4679}), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_407 ( .clk (clk), .D ({signal_1945, signal_998}), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    DFF_X1 cell_789 ( .CK (clk), .D (signal_4689), .Q (signal_1001), .QN () ) ;
    DFF_X1 cell_791 ( .CK (clk), .D (signal_4697), .Q (signal_1002), .QN () ) ;
    DFF_X1 cell_793 ( .CK (clk), .D (signal_4705), .Q (signal_1003), .QN () ) ;
    DFF_X1 cell_795 ( .CK (clk), .D (signal_4713), .Q (signal_1004), .QN () ) ;
    DFF_X1 cell_797 ( .CK (clk), .D (signal_4721), .Q (signal_1005), .QN () ) ;
    DFF_X1 cell_799 ( .CK (clk), .D (signal_4729), .Q (signal_1006), .QN () ) ;
    DFF_X1 cell_801 ( .CK (clk), .D (signal_4737), .Q (signal_1007), .QN () ) ;
    DFF_X1 cell_814 ( .CK (clk), .D (signal_4745), .Q (signal_1015), .QN () ) ;
    DFF_X1 cell_816 ( .CK (clk), .D (signal_4753), .Q (signal_1016), .QN () ) ;
    DFF_X1 cell_818 ( .CK (clk), .D (signal_4761), .Q (done), .QN () ) ;
endmodule
